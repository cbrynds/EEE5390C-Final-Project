/*module AND2X1 (Y, A, B);
	output Y;
	input A, B;

	// Function
	and (Y, A, B);

	// Timing
	specify
		(A => Y) = 0;
		(B => Y) = 0;
	endspecify
endmodule*/

module AND2X1 (Y, A, B);
	output Y;
	input A, B;

	// Function
	reg Y=0;
	always@(*) begin
		Y = A&B;
	end
endmodule
/*module AND2XL (Y, A, B);
	output Y;
	input A, B;

	// Function
	and (Y, A, B);

	// Timing
	specify
		(A => Y) = 0;
		(B => Y) = 0;
	endspecify
endmodule*/

module AND2XL (Y, A, B);
	output Y;
	input A, B;

	// Function
	assign Y = A & B;
endmodule
/*module AOI21X1 (Y, A0, A1, B0);
	output Y;
	input A0, A1, B0;

	// Function
	wire int_fwire_0, int_fwire_1;

	and (int_fwire_0, A0, A1);
	or (int_fwire_1, int_fwire_0, B0);
	not (Y, int_fwire_1);

	// Timing
	specify
		(A0 => Y) = 0;
		(A1 => Y) = 0;
		(B0 => Y) = 0;
	endspecify
endmodule*/


module AOI21X1 (Y, A0, A1, B0);
	output Y;
	input A0, A1, B0;

	// Function
	reg Y=0;
	always@(*) begin
		Y = ~((A0&A1)|B0);
	end
endmodule
/*module AOI22X1 (Y, A0, A1, B0, B1);
	output Y;
	input A0, A1, B0, B1;

	// Function
	wire int_fwire_0, int_fwire_1, int_fwire_2;

	and (int_fwire_0, A0, A1);
	and (int_fwire_1, B0, B1);
	or (int_fwire_2, int_fwire_1, int_fwire_0);
	not (Y, int_fwire_2);

	// Timing
	specify
		(A0 => Y) = 0;
		(A1 => Y) = 0;
		(B0 => Y) = 0;
		(B1 => Y) = 0;
	endspecify
endmodule*/


module AOI22X1 (Y, A0, A1, B0, B1);
	output Y;
	input A0, A1, B0, B1;

	// Function
	reg Y=0;
	always@(*) begin
		Y = ~((A0&A1)|(B0&B1));
	end
endmodule
module BUFX1 (Y, A);
        output Y;
        input A;

 

        assign Y = A;
endmodule
/*module BUFX3 (Y, A);
	output Y;
	input A;

	// Function
	buf (Y, A);

	// Timing
	specify
		(A => Y) = 0;
	endspecify
endmodule*/


module BUFX3 (Y, A);
	output Y;
	input A;

	assign Y = A;
endmodule
/*module CLKBUFX2 (Y, A);
	output Y;
	input A;

	// Function
	buf (Y, A);

	// Timing
	specify
		(A => Y) = 0;
	endspecify
endmodule*/


module CLKBUFX2 (Y, A);
	output Y;
	input A;

	// Function
	reg Y=0;
	always@(*) begin
		Y <= A;
	end

endmodule
/*module DFFHQX1 (Q, D, CK);
	output Q;
	input D, CK;
	reg notifier;
	wire delayed_D, delayed_CK;

	// Function
	wire int_fwire_N30, xcr_0;

	altos_dff_err (xcr_0, delayed_CK, delayed_D);
	altos_dff (int_fwire_N30, notifier, delayed_CK, delayed_D, xcr_0);
	buf (Q, int_fwire_N30);

	// Timing
	specify
		(posedge CK => (Q+:D)) = 0;
		$setuphold (posedge CK, posedge D, 0, 0, notifier,,, delayed_CK, delayed_D);
		$setuphold (posedge CK, negedge D, 0, 0, notifier,,, delayed_CK, delayed_D);
		$width (posedge CK, 0, 0, notifier);
		$width (negedge CK, 0, 0, notifier);
	endspecify
endmodule*/


module DFFHQX1 (Q, D, CK);
	output Q;
	input D, CK;

	// Function
	reg Q=0;
	always@(posedge CK) begin
		Q <= D;
	end
endmodule
/*module DFFRHQX1 (Q, D, RN, CK);
	output Q;
	input D, RN, CK;
	reg notifier;
	wire delayed_D, delayed_CK;

	// Function
	wire int_fwire_N30, int_fwire_r, xcr_0;

	not (int_fwire_r, RN);
	altos_dff_r_err (xcr_0, delayed_CK, delayed_D, int_fwire_r);
	altos_dff_r (int_fwire_N30, notifier, delayed_CK, delayed_D, int_fwire_r, xcr_0);
	buf (Q, int_fwire_N30);

	// Timing
	specify
		(negedge RN => (Q+:1'b0)) = 0;
		(posedge CK => (Q+:D)) = 0;
		$setuphold (posedge CK, posedge D, 0, 0, notifier,,, delayed_CK, delayed_D);
		$setuphold (posedge CK, negedge D, 0, 0, notifier,,, delayed_CK, delayed_D);
		$recovery (posedge RN, posedge CK, 0, notifier);
		$hold (posedge CK, posedge RN, 0, notifier);
		$width (negedge RN, 0, 0, notifier);
		$width (posedge CK, 0, 0, notifier);
		$width (negedge CK, 0, 0, notifier);
	endspecify
endmodule*/



module DFFRHQX1 (Q, D, RN, CK);
	output Q;
	input D, RN, CK;
	
	// Function
	reg Q=0;
	always@(posedge CK or negedge RN) begin
		if(!RN) begin
			Q <= 0;
		end
		else begin
			Q <= D;
		end
	end
endmodule
/*module DFFRX1 (Q, QN, D, RN, CK);
	output Q, QN;
	input D, RN, CK;
	reg notifier;
	wire delayed_D, delayed_CK;

	// Function
	wire int_fwire_N30, int_fwire_QBINT, int_fwire_r;
	wire xcr_0;

	not (int_fwire_r, RN);
	altos_dff_r_err (xcr_0, delayed_CK, delayed_D, int_fwire_r);
	altos_dff_r (int_fwire_N30, notifier, delayed_CK, delayed_D, int_fwire_r, xcr_0);
	buf (Q, int_fwire_N30);
	not (int_fwire_QBINT, int_fwire_N30);
	buf (QN, int_fwire_QBINT);

	// Timing
	specify
		(negedge RN => (Q+:1'b0)) = 0;
		(posedge CK => (Q+:D)) = 0;
		(negedge RN => (QN-:1'b0)) = 0;
		(posedge CK => (QN-:D)) = 0;
		$setuphold (posedge CK, posedge D, 0, 0, notifier,,, delayed_CK, delayed_D);
		$setuphold (posedge CK, negedge D, 0, 0, notifier,,, delayed_CK, delayed_D);
		$recovery (posedge RN, posedge CK, 0, notifier);
		$hold (posedge CK, posedge RN, 0, notifier);
		$width (negedge RN, 0, 0, notifier);
		$width (posedge CK, 0, 0, notifier);
		$width (negedge CK, 0, 0, notifier);
	endspecify
endmodule*/


module DFFRX1 (Q, QN, D, RN, CK);
	output Q, QN;
	input D, RN, CK;

	reg Q=0;
	wire QN;
	always@(posedge CK or negedge RN) begin
		if(!RN) begin
			Q <= 0;
		end
		else begin
			Q <= D;
		end
	end

	assign QN = !Q;
endmodule
/*module DFFRXL (Q, QN, D, RN, CK);
	output Q, QN;
	input D, RN, CK;
	reg notifier;
	wire delayed_D, delayed_CK;

	// Function
	wire int_fwire_N30, int_fwire_QBINT, int_fwire_r;
	wire xcr_0;

	not (int_fwire_r, RN);
	altos_dff_r_err (xcr_0, delayed_CK, delayed_D, int_fwire_r);
	altos_dff_r (int_fwire_N30, notifier, delayed_CK, delayed_D, int_fwire_r, xcr_0);
	buf (Q, int_fwire_N30);
	not (int_fwire_QBINT, int_fwire_N30);
	buf (QN, int_fwire_QBINT);

	// Timing
	specify
		(negedge RN => (Q+:1'b0)) = 0;
		(posedge CK => (Q+:D)) = 0;
		(negedge RN => (QN-:1'b0)) = 0;
		(posedge CK => (QN-:D)) = 0;
		$setuphold (posedge CK, posedge D, 0, 0, notifier,,, delayed_CK, delayed_D);
		$setuphold (posedge CK, negedge D, 0, 0, notifier,,, delayed_CK, delayed_D);
		$recovery (posedge RN, posedge CK, 0, notifier);
		$hold (posedge CK, posedge RN, 0, notifier);
		$width (negedge RN, 0, 0, notifier);
		$width (posedge CK, 0, 0, notifier);
		$width (negedge CK, 0, 0, notifier);
	endspecify
endmodule*/

module DFFRXL (Q, QN, D, RN, CK);
	output Q, QN;
	input D, RN, CK;
	reg Q=0;
	wire QN;

	always@(posedge CK or negedge RN) begin
		if(!RN) begin
			Q <= 0;		
		end
		else begin
			Q <= D;
		end
	end
	assign QN = ~Q;
	
endmodule
/*module DFFSHQX1 (Q, D, SN, CK);
	output Q;
	input D, SN, CK;
	reg notifier;
	wire delayed_D, delayed_CK;

	// Function
	wire int_fwire_N35, int_fwire_s, xcr_0;

	not (int_fwire_s, SN);
	altos_dff_s_err (xcr_0, delayed_CK, delayed_D, int_fwire_s);
	altos_dff_s (int_fwire_N35, notifier, delayed_CK, delayed_D, int_fwire_s, xcr_0);
	buf (Q, int_fwire_N35);

	// Timing
	specify
		(negedge SN => (Q+:1'b1)) = 0;
		(posedge CK => (Q+:D)) = 0;
		$setuphold (posedge CK, posedge D, 0, 0, notifier,,, delayed_CK, delayed_D);
		$setuphold (posedge CK, negedge D, 0, 0, notifier,,, delayed_CK, delayed_D);
		$recovery (posedge SN, posedge CK, 0, notifier);
		$hold (posedge CK, posedge SN, 0, notifier);
		$width (negedge SN, 0, 0, notifier);
		$width (posedge CK, 0, 0, notifier);
		$width (negedge CK, 0, 0, notifier);
	endspecify
endmodule*/

module DFFSHQX1 (Q, D, SN, CK);
	output Q;
	input D, SN, CK;

	// Function
	reg Q = 0;
	always@(posedge CK or negedge SN) begin
		if(!SN) begin
			Q <= 1;		
		end
		else begin
			Q <= D;
		end
	end
endmodule
/*module INVX1 (Y, A);
	output Y;
	input A;

	// Function
	not (Y, A);

	// Timing
	specify
		(A => Y) = 0;
	endspecify
endmodule*/

module INVX1 (Y, A);
	output Y;
	input A;

	// Function
	reg Y=0;
	always@(*) begin
		Y = ~A;
	end
endmodule
/*module INVX2 (Y, A);
	output Y;
	input A;

	// Function
	not (Y, A);

	// Timing
	specify
		(A => Y) = 0;
	endspecify
endmodule*/


module INVX2 (Y, A);
	output Y;
	input A;

	reg Y=0;
	// Function
	always@(*) begin
		Y = ~A;	
	end

endmodule
/*module INVX4 (Y, A);
	output Y;
	input A;

	// Function
	not (Y, A);

	// Timing
	specify
		(A => Y) = 0;
	endspecify
endmodule*/

module INVX4 (Y, A);
	output Y;
	input A;

	// Function
	assign Y = ~A;	
endmodule
/*module INVX8 (Y, A);
	output Y;
	input A;

	// Function
	not (Y, A);

	// Timing
	specify
		(A => Y) = 0;
	endspecify
endmodule*/

module INVX8 (Y, A);
	output Y;
	input A;

	assign Y = ~A;
endmodule
/*module INVXL (Y, A);
	output Y;
	input A;

	// Function
	not (Y, A);

	// Timing
	specify
		(A => Y) = 0;
	endspecify
endmodule*/


module INVXL (Y, A);
	output Y;
	input A;

	// Function
	assign Y = ~A;
endmodule
/*module MX2X1 (Y, A, B, S0);
	output Y;
	input A, B, S0;

	// Function
	wire int_fwire_0, int_fwire_1, S0__bar;

	not (S0__bar, S0);
	and (int_fwire_0, S0__bar, A);
	and (int_fwire_1, S0, B);
	or (Y, int_fwire_1, int_fwire_0);

	// Timing
	specify
		(A => Y) = 0;
		(B => Y) = 0;
		(posedge S0 => (Y:S0)) = 0;
		(negedge S0 => (Y:S0)) = 0;
	endspecify
endmodule*/


module MX2X1 (Y, A, B, S0);
	output Y;
	input A, B, S0;

	// Function
	reg Y=0;
	always@(*) begin
		Y = (~S0&A)|(S0&B);
	end
endmodule
/*module NAND2X1 (Y, A, B);
	output Y;
	input A, B;

	// Function
	wire int_fwire_0;

	and (int_fwire_0, A, B);
	not (Y, int_fwire_0);

	// Timing
	specify
		(A => Y) = 0;
		(B => Y) = 0;
	endspecify
endmodule*/


module NAND2X1 (Y, A, B);
	output Y;
	input A, B;

	// Function
	reg Y=0;
	always@(*) begin
		Y = ~(A&B);
	end
endmodule
/*module NAND2X2 (Y, A, B);
	output Y;
	input A, B;

	// Function
	wire int_fwire_0;

	and (int_fwire_0, A, B);
	not (Y, int_fwire_0);

	// Timing
	specify
		(A => Y) = 0;
		(B => Y) = 0;
	endspecify
endmodule
*/
module NAND2X2 (Y, A, B);
	output Y;
	input A, B;

	// Function
	reg Y=0;

	always@(*) begin
		Y = ~(A&B);
	end
endmodule
/*module NAND2XL (Y, A, B);
	output Y;
	input A, B;

	// Function
	wire int_fwire_0;

	and (int_fwire_0, A, B);
	not (Y, int_fwire_0);

	// Timing
	specify
		(A => Y) = 0;
		(B => Y) = 0;
	endspecify
endmodule*/

module NAND2XL (Y, A, B);
	output Y;
	input A, B;

	// Function
	assign Y = ~(A&B);
endmodule
/*module NAND3X1 (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	wire int_fwire_0;

	and (int_fwire_0, A, B, C);
	not (Y, int_fwire_0);

	// Timing
	specify
		(A => Y) = 0;
		(B => Y) = 0;
		(C => Y) = 0;
	endspecify
endmodule*/


module NAND3X1 (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	reg Y=0;
	always@(*) begin
		Y = ~(A&B&C);
	end
endmodule
/*module NAND4X1 (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	wire int_fwire_0;

	and (int_fwire_0, A, B, C, D);
	not (Y, int_fwire_0);

	// Timing
	specify
		(A => Y) = 0;
		(B => Y) = 0;
		(C => Y) = 0;
		(D => Y) = 0;
	endspecify
endmodule*/


module NAND4X1 (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	reg Y=0;
	always@(*) begin
		Y = ~(A&B&C&D);
	end
endmodule
/*module NOR2X1 (Y, A, B);
	output Y;
	input A, B;

	// Function
	wire int_fwire_0;

	or (int_fwire_0, A, B);
	not (Y, int_fwire_0);

	// Timing
	specify
		(A => Y) = 0;
		(B => Y) = 0;
	endspecify
endmodule*/

module NOR2X1 (Y, A, B);
	output Y;
	input A, B;

	// Function
	reg Y=0;
	always@(*) begin
		Y = ~(A|B);
	end
endmodule
/*module NOR2X2 (Y, A, B);
	output Y;
	input A, B;

	// Function
	wire int_fwire_0;

	or (int_fwire_0, A, B);
	not (Y, int_fwire_0);

	// Timing
	specify
		(A => Y) = 0;
		(B => Y) = 0;
	endspecify
endmodule*/

module NOR2X2 (Y, A, B);
	output Y;
	input A, B;

	// Function
	assign Y = ~(A|B);
endmodule
/*module NOR2XL (Y, A, B);
	output Y;
	input A, B;

	// Function
	wire int_fwire_0;

	or (int_fwire_0, A, B);
	not (Y, int_fwire_0);

	// Timing
	specify
		(A => Y) = 0;
		(B => Y) = 0;
	endspecify
endmodule*/

module NOR2XL (Y, A, B);
	output Y;
	input A, B;

	// Function
	assign Y = ~(A|B);
endmodule
/*module NOR3X1 (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	wire int_fwire_0;

	or (int_fwire_0, A, B, C);
	not (Y, int_fwire_0);

	// Timing
	specify
		(A => Y) = 0;
		(B => Y) = 0;
		(C => Y) = 0;
	endspecify
endmodule*/

module NOR3X1 (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	reg Y=0;
	always@(*) begin
		Y = ~(A|B|C);
	end

endmodule
/*module NOR4X1 (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	wire int_fwire_0;

	or (int_fwire_0, A, B, C, D);
	not (Y, int_fwire_0);

	// Timing
	specify
		(A => Y) = 0;
		(B => Y) = 0;
		(C => Y) = 0;
		(D => Y) = 0;
	endspecify
endmodule*/


module NOR4X1 (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	reg Y=0;
	always@(*) begin
		Y = ~(A|B|C|D);
	end
endmodule
/*module OAI21X1 (Y, A0, A1, B0);
	output Y;
	input A0, A1, B0;

	// Function
	wire int_fwire_0, int_fwire_1;

	or (int_fwire_0, A0, A1);
	and (int_fwire_1, int_fwire_0, B0);
	not (Y, int_fwire_1);

	// Timing
	specify
		(A0 => Y) = 0;
		(A1 => Y) = 0;
		(B0 => Y) = 0;
	endspecify
endmodule*/


module OAI21X1 (Y, A0, A1, B0);
	output Y;
	input A0, A1, B0;

	// Function
	reg Y=0;
	always@(*) begin
		Y = ~((A0|A1)&B0);
	end
endmodule
/*module OAI22X1 (Y, A0, A1, B0, B1);
	output Y;
	input A0, A1, B0, B1;

	// Function
	wire int_fwire_0, int_fwire_1, int_fwire_2;

	or (int_fwire_0, A0, A1);
	or (int_fwire_1, B0, B1);
	and (int_fwire_2, int_fwire_1, int_fwire_0);
	not (Y, int_fwire_2);

	// Timing
	specify
		(A0 => Y) = 0;
		(A1 => Y) = 0;
		(B0 => Y) = 0;
		(B1 => Y) = 0;
	endspecify
endmodule*/


module OAI22X1 (Y, A0, A1, B0, B1);
	output Y;
	input A0, A1, B0, B1;

	// Function
	reg Y=0;
	always@(*) begin
		Y = ~((A0|A1)&(B0|B1));
	end
	
endmodule
/*module OAI33X1 (Y, A0, A1, A2, B0, B1, B2);
	output Y;
	input A0, A1, A2, B0, B1, B2;

	// Function
	wire int_fwire_0, int_fwire_1, int_fwire_2;

	or (int_fwire_0, A0, A1, A2);
	or (int_fwire_1, B0, B1, B2);
	and (int_fwire_2, int_fwire_1, int_fwire_0);
	not (Y, int_fwire_2);

	// Timing
	specify
		(A0 => Y) = 0;
		(A1 => Y) = 0;
		(A2 => Y) = 0;
		(B0 => Y) = 0;
		(B1 => Y) = 0;
		(B2 => Y) = 0;
	endspecify
endmodule*/


module OAI33X1 (Y, A0, A1, A2, B0, B1, B2);
	output Y;
	input A0, A1, A2, B0, B1, B2;

	// Function
	reg Y=0;
	always@(*) begin
		Y = ~((A0|A1|A2)&(B0|B1|B2));
	end
endmodule
/*module OR2X1 (Y, A, B);
	output Y;
	input A, B;

	// Function
	or (Y, A, B);

	// Timing
	specify
		(A => Y) = 0;
		(B => Y) = 0;
	endspecify
endmodule*/


module OR2X1 (Y, A, B);
	output Y;
	input A, B;

	// Function
	reg Y=0;
	always@(*) begin
		Y = A|B;
	end
endmodule
/*module OR2XL (Y, A, B);
	output Y;
	input A, B;

	// Function
	or (Y, A, B);

	// Timing
	specify
		(A => Y) = 0;
		(B => Y) = 0;
	endspecify
endmodule*/

module OR2XL (Y, A, B);
	output Y;
	input A, B;

	// Function
	assign Y = A|B;
endmodule
/*module OR4X1 (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	or (Y, A, B, C, D);

	// Timing
	specify
		(A => Y) = 0;
		(B => Y) = 0;
		(C => Y) = 0;
		(D => Y) = 0;
	endspecify
endmodule*/


module OR4X1 (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	reg Y=0;
	always@(*) begin
		Y = (A|B|C|D);
	end
endmodule
/*module SDFFQX1 (Q, D, SE, SI, CK);
	output Q;
	input D, SE, SI, CK;
	reg notifier;
	wire delayed_D, delayed_SE, delayed_SI, delayed_CK;

	// Function
	wire delayed_SE__bar, int_fwire_0, int_fwire_1;
	wire int_fwire_d, int_fwire_N30, xcr_0;

	not (delayed_SE__bar, delayed_SE);
	and (int_fwire_0, delayed_SE__bar, delayed_D);
	and (int_fwire_1, delayed_SE, delayed_SI);
	or (int_fwire_d, int_fwire_1, int_fwire_0);
	altos_dff_err (xcr_0, delayed_CK, int_fwire_d);
	altos_dff (int_fwire_N30, notifier, delayed_CK, int_fwire_d, xcr_0);
	buf (Q, int_fwire_N30);

	// Timing
	specify
		(posedge CK => (Q+:((SE && SI) || (!SE && D)))) = 0;
		$setuphold (posedge CK, posedge D, 0, 0, notifier,,, delayed_CK, delayed_D);
		$setuphold (posedge CK, negedge D, 0, 0, notifier,,, delayed_CK, delayed_D);
		$setuphold (posedge CK, posedge SE, 0, 0, notifier,,, delayed_CK, delayed_SE);
		$setuphold (posedge CK, negedge SE, 0, 0, notifier,,, delayed_CK, delayed_SE);
		$setuphold (posedge CK, posedge SI, 0, 0, notifier,,, delayed_CK, delayed_SI);
		$setuphold (posedge CK, negedge SI, 0, 0, notifier,,, delayed_CK, delayed_SI);
		$width (posedge CK, 0, 0, notifier);
		$width (negedge CK, 0, 0, notifier);
	endspecify
endmodule*/

module SDFFQX1 (Q, D, SE, SI, CK);
	output Q;
	input D, SE, SI, CK;
	
	reg Q=0;
	always@(posedge CK) begin
		Q <= (SE & SI) | (~SE & D);
	end

endmodule
/*module SDFFRHQX1 (Q, D, SE, SI, RN, CK);
	output Q;
	input D, SE, SI, RN, CK;
	reg notifier;
	wire delayed_D, delayed_SE, delayed_SI, delayed_CK;

	// Function
	wire delayed_SE__bar, int_fwire_0, int_fwire_1;
	wire int_fwire_d, int_fwire_N30, int_fwire_r;
	wire xcr_0;

	not (delayed_SE__bar, delayed_SE);
	and (int_fwire_0, delayed_SE__bar, delayed_D);
	and (int_fwire_1, delayed_SE, delayed_SI);
	or (int_fwire_d, int_fwire_1, int_fwire_0);
	not (int_fwire_r, RN);
	altos_dff_r_err (xcr_0, delayed_CK, int_fwire_d, int_fwire_r);
	altos_dff_r (int_fwire_N30, notifier, delayed_CK, int_fwire_d, int_fwire_r, xcr_0);
	buf (Q, int_fwire_N30);

	// Timing
	specify
		(negedge RN => (Q+:1'b0)) = 0;
		(posedge CK => (Q+:((SE && SI) || (!SE && D)))) = 0;
		$setuphold (posedge CK, posedge D, 0, 0, notifier,,, delayed_CK, delayed_D);
		$setuphold (posedge CK, negedge D, 0, 0, notifier,,, delayed_CK, delayed_D);
		$setuphold (posedge CK, posedge SE, 0, 0, notifier,,, delayed_CK, delayed_SE);
		$setuphold (posedge CK, negedge SE, 0, 0, notifier,,, delayed_CK, delayed_SE);
		$setuphold (posedge CK, posedge SI, 0, 0, notifier,,, delayed_CK, delayed_SI);
		$setuphold (posedge CK, negedge SI, 0, 0, notifier,,, delayed_CK, delayed_SI);
		$recovery (posedge RN, posedge CK, 0, notifier);
		$hold (posedge CK, posedge RN, 0, notifier);
		$width (negedge RN, 0, 0, notifier);
		$width (posedge CK, 0, 0, notifier);
		$width (negedge CK, 0, 0, notifier);
	endspecify
endmodule*/

module SDFFRHQX1 (Q, D, SE, SI, RN, CK);
	output Q;
	input D, SE, SI, RN, CK;

	reg Q=0;

	always@(posedge CK or negedge RN) begin
		if(!RN) begin
			Q <= 0;
		end
		else begin
			Q <= (~SE & D) | (SE & SI);
		end
	end
endmodule
/*module SDFFSXL (Q, QN, D, SE, SI, SN, CK);
	output Q, QN;
	input D, SE, SI, SN, CK;
	reg notifier;
	wire delayed_D, delayed_SE, delayed_SI, delayed_CK;

	// Function
	wire delayed_SE__bar, int_fwire_0, int_fwire_1;
	wire int_fwire_d, int_fwire_N35, int_fwire_QBINT;
	wire int_fwire_s, xcr_0;

	not (delayed_SE__bar, delayed_SE);
	and (int_fwire_0, delayed_SE__bar, delayed_D);
	and (int_fwire_1, delayed_SE, delayed_SI);
	or (int_fwire_d, int_fwire_1, int_fwire_0);
	not (int_fwire_s, SN);
	altos_dff_s_err (xcr_0, delayed_CK, int_fwire_d, int_fwire_s);
	altos_dff_s (int_fwire_N35, notifier, delayed_CK, int_fwire_d, int_fwire_s, xcr_0);
	buf (Q, int_fwire_N35);
	not (int_fwire_QBINT, int_fwire_N35);
	buf (QN, int_fwire_QBINT);

	// Timing
	specify
		(negedge SN => (Q+:1'b1)) = 0;
		(posedge CK => (Q+:((SE && SI) || (!SE && D)))) = 0;
		(negedge SN => (QN-:1'b1)) = 0;
		(posedge CK => (QN-:((SE && SI) || (!SE && D)))) = 0;
		$setuphold (posedge CK, posedge D, 0, 0, notifier,,, delayed_CK, delayed_D);
		$setuphold (posedge CK, negedge D, 0, 0, notifier,,, delayed_CK, delayed_D);
		$setuphold (posedge CK, posedge SE, 0, 0, notifier,,, delayed_CK, delayed_SE);
		$setuphold (posedge CK, negedge SE, 0, 0, notifier,,, delayed_CK, delayed_SE);
		$setuphold (posedge CK, posedge SI, 0, 0, notifier,,, delayed_CK, delayed_SI);
		$setuphold (posedge CK, negedge SI, 0, 0, notifier,,, delayed_CK, delayed_SI);
		$recovery (posedge SN, posedge CK, 0, notifier);
		$hold (posedge CK, posedge SN, 0, notifier);
		$width (negedge SN, 0, 0, notifier);
		$width (posedge CK, 0, 0, notifier);
		$width (negedge CK, 0, 0, notifier);
	endspecify
endmodule*/

module SDFFSRX2 (Q, QN, D, SE, SI, RN, SN, CK);
	output Q, QN;
	input D, SE, SI, SN, CK, RN;

	reg Q = 0;
	wire QN;
	always@(posedge CK or negedge SN) begin
		if(!SN) begin
			Q <= 1;		
		end
    else if (!RN) begin
      Q <= 0;
    end
		else begin
			Q <= (SE & SI) | (~SE & D);
		end
	end
	assign QN = ~Q;
endmodule
/*module SDFFSXL (Q, QN, D, SE, SI, SN, CK);
	output Q, QN;
	input D, SE, SI, SN, CK;
	reg notifier;
	wire delayed_D, delayed_SE, delayed_SI, delayed_CK;

	// Function
	wire delayed_SE__bar, int_fwire_0, int_fwire_1;
	wire int_fwire_d, int_fwire_N35, int_fwire_QBINT;
	wire int_fwire_s, xcr_0;

	not (delayed_SE__bar, delayed_SE);
	and (int_fwire_0, delayed_SE__bar, delayed_D);
	and (int_fwire_1, delayed_SE, delayed_SI);
	or (int_fwire_d, int_fwire_1, int_fwire_0);
	not (int_fwire_s, SN);
	altos_dff_s_err (xcr_0, delayed_CK, int_fwire_d, int_fwire_s);
	altos_dff_s (int_fwire_N35, notifier, delayed_CK, int_fwire_d, int_fwire_s, xcr_0);
	buf (Q, int_fwire_N35);
	not (int_fwire_QBINT, int_fwire_N35);
	buf (QN, int_fwire_QBINT);

	// Timing
	specify
		(negedge SN => (Q+:1'b1)) = 0;
		(posedge CK => (Q+:((SE && SI) || (!SE && D)))) = 0;
		(negedge SN => (QN-:1'b1)) = 0;
		(posedge CK => (QN-:((SE && SI) || (!SE && D)))) = 0;
		$setuphold (posedge CK, posedge D, 0, 0, notifier,,, delayed_CK, delayed_D);
		$setuphold (posedge CK, negedge D, 0, 0, notifier,,, delayed_CK, delayed_D);
		$setuphold (posedge CK, posedge SE, 0, 0, notifier,,, delayed_CK, delayed_SE);
		$setuphold (posedge CK, negedge SE, 0, 0, notifier,,, delayed_CK, delayed_SE);
		$setuphold (posedge CK, posedge SI, 0, 0, notifier,,, delayed_CK, delayed_SI);
		$setuphold (posedge CK, negedge SI, 0, 0, notifier,,, delayed_CK, delayed_SI);
		$recovery (posedge SN, posedge CK, 0, notifier);
		$hold (posedge CK, posedge SN, 0, notifier);
		$width (negedge SN, 0, 0, notifier);
		$width (posedge CK, 0, 0, notifier);
		$width (negedge CK, 0, 0, notifier);
	endspecify
endmodule*/

module SDFFSXL (Q, QN, D, SE, SI, SN, CK);
	output Q, QN;
	input D, SE, SI, SN, CK;

	reg Q = 0;
	wire QN;
	always@(posedge CK or negedge SN) begin
		if(!SN) begin
			Q <= 1;		
		end
		else begin
			Q <= (SE & SI) | (~SE & D);
		end
	end
	assign QN = ~Q;
endmodule
module TLATNX1 (  input D,
                  input GN,
                  output QN,
                  output reg Q=0);

 

   always @ (D or GN)
      if (!GN)
         Q <= D;

 

   assign QN = !Q;
endmodule
/*module TLATX1 (Q, QN, D, G);
	output Q, QN;
	input D, G;
	reg notifier;
	wire delayed_D, delayed_G;

	// Function
	wire int_fwire_N0, int_fwire_QINT;

	altos_latch (int_fwire_QINT, notifier, delayed_G, delayed_D);
	buf (Q, int_fwire_QINT);
	not (int_fwire_N0, int_fwire_QINT);
	buf (QN, int_fwire_N0);

	// Timing
	specify
		(D => Q) = 0;
		(posedge G => (Q+:D)) = 0;
		(D => QN) = 0;
		(posedge G => (QN-:D)) = 0;
		$setuphold (negedge G, posedge D, 0, 0, notifier,,, delayed_G, delayed_D);
		$setuphold (negedge G, negedge D, 0, 0, notifier,,, delayed_G, delayed_D);
		$width (posedge G, 0, 0, notifier);
	endspecify
endmodule*/

module TLATX1 (Q, QN, D, G);
	output Q, QN;
	input D, G;
	
	reg Q = 0;
	always @ (D or G) begin
		if(G) begin
			Q <= D;
		end
	end

	assign QN = !Q;
endmodule
/*module XNOR2X1 (Y, A, B);
	output Y;
	input A, B;

	// Function
	wire int_fwire_0;

	xor (int_fwire_0, A, B);
	not (Y, int_fwire_0);

	// Timing
	specify
		(posedge A => (Y:A)) = 0;
		(negedge A => (Y:A)) = 0;
		(posedge B => (Y:B)) = 0;
		(negedge B => (Y:B)) = 0;
	endspecify
endmodule*/


module XNOR2X1 (Y, A, B);
	output Y;
	input A, B;

	// Function
	reg Y=0;
	always@(*) begin
		Y = ~(A^B);
	end
endmodule
/*module XOR2X1 (Y, A, B);
	output Y;
	input A, B;

	// Function
	xor (Y, A, B);

	// Timing
	specify
		(posedge A => (Y:A)) = 0;
		(negedge A => (Y:A)) = 0;
		(posedge B => (Y:B)) = 0;
		(negedge B => (Y:B)) = 0;
	endspecify
endmodule*/


module XOR2X1 (Y, A, B);
	output Y;
	input A, B;

	// Function
	reg Y=0;
	always@(*) begin
		Y = (A^B);
	end
endmodule
/*module XOR2XL (Y, A, B);
	output Y;
	input A, B;

	// Function
	xor (Y, A, B);

	// Timing
	specify
		(posedge A => (Y:A)) = 0;
		(negedge A => (Y:A)) = 0;
		(posedge B => (Y:B)) = 0;
		(negedge B => (Y:B)) = 0;
	endspecify
endmodule*/

module XOR2XL (Y, A, B);
	output Y;
	input A, B;

	// Function
	assign Y = A^B;
endmodule
/////////////////////////////////////////////////////////////
// Created by: Synopsys DC Expert(TM) in wire load mode
// Version   : R-2020.09-SP4
// Date      : Wed May  4 17:40:46 2022
/////////////////////////////////////////////////////////////


module riscv_core ( clk_i, rst_i, mem_d_data_rd_i, mem_d_accept_i, mem_d_ack_i, 
        mem_d_error_i, mem_d_resp_tag_i, mem_i_accept_i, mem_i_valid_i, 
        mem_i_error_i, mem_i_inst_i, intr_i, reset_vector_i, cpu_id_i, 
        mem_d_addr_o, mem_d_data_wr_o, mem_d_rd_o, mem_d_wr_o, 
        mem_d_cacheable_o, mem_d_req_tag_o, mem_d_invalidate_o, mem_d_flush_o, 
        mem_i_rd_o, mem_i_flush_o, mem_i_invalidate_o, mem_i_pc_o,
        challenge );
  input [31:0] mem_d_data_rd_i;
  input [10:0] mem_d_resp_tag_i;
  input [31:0] mem_i_inst_i;
  input [31:0] reset_vector_i;
  input [31:0] cpu_id_i;
  output [31:0] mem_d_addr_o;
  output [31:0] mem_d_data_wr_o;
  output [3:0] mem_d_wr_o;
  output [10:0] mem_d_req_tag_o;
  output [31:0] mem_i_pc_o;
  input [107:0] challenge;
  input clk_i, rst_i, mem_d_accept_i, mem_d_ack_i, mem_d_error_i,
         mem_i_accept_i, mem_i_valid_i, mem_i_error_i, intr_i;
  output mem_d_rd_o, mem_d_cacheable_o, mem_d_invalidate_o, mem_d_flush_o,
         mem_i_rd_o, mem_i_flush_o, mem_i_invalidate_o;
  parameter wm_select = 1'b1;
  wire   n8572, n8805, n8886, n8561, u_fetch_icache_fetch_q, n8555, n8556,
         u_mmu_N235, net1802, u_mmu_pte_entry_q_1, u_mmu_N236,
         u_mmu_pte_entry_q_2, u_mmu_N237, u_mmu_pte_entry_q_3, u_mmu_N238,
         u_mmu_pte_entry_q_4, u_mmu_N249, u_mmu_N250, n8550, n8549, n8548,
         n8547, n8546, n8545, n8544, n8543, n8445, n8558, u_arb_read_hold_q,
         n8557, u_arb_src_mmu_q, n8539, n8552, u_mmu_virt_addr_q_31,
         u_mmu_virt_addr_q_30, u_mmu_virt_addr_q_29, u_mmu_virt_addr_q_28,
         n8444, u_fetch_N80, \mmu_ifetch_pc_w[31] , u_fetch_N52, u_fetch_N53,
         u_fetch_N54, u_fetch_N55, u_fetch_N56, u_fetch_N57, u_fetch_N58,
         u_fetch_N59, u_fetch_N60, u_fetch_N61, u_fetch_N62, u_fetch_N63,
         u_fetch_N64, u_fetch_N65, u_fetch_N66, u_fetch_N67, u_fetch_N68,
         u_fetch_N69, u_fetch_N70, u_fetch_N71, u_fetch_N72, u_fetch_N73,
         u_fetch_N74, u_fetch_N75, u_fetch_N76, u_fetch_N77, u_fetch_N78,
         u_fetch_N79, u_decode_N320, u_decode_u_regfile_N981, u_muldiv_N262,
         net1913, u_decode_u_regfile_N944, n8520, u_muldiv_invert_res_q,
         u_decode_u_regfile_N988, u_muldiv_N232, net1908,
         u_decode_u_regfile_N982, n8443, u_fetch_active_q, u_fetch_N15,
         u_fetch_branch_valid_q, u_decode_N305, u_decode_u_regfile_N966,
         u_muldiv_N247, u_decode_u_regfile_N929, u_muldiv_N311, net1893,
         u_muldiv_N310, u_muldiv_N309, u_muldiv_N308, u_muldiv_N307,
         u_muldiv_N306, u_muldiv_N305, u_muldiv_N304, u_muldiv_N303,
         u_muldiv_N302, u_muldiv_N301, u_muldiv_N300, u_muldiv_N299,
         u_muldiv_N298, u_muldiv_N297, u_muldiv_N296, net1888, u_muldiv_N295,
         u_muldiv_N294, u_muldiv_N293, u_muldiv_N292, u_muldiv_N291,
         u_muldiv_N290, u_muldiv_N289, u_muldiv_N288, u_muldiv_N287,
         u_muldiv_N286, u_muldiv_N285, u_muldiv_N284, u_muldiv_N283,
         u_muldiv_N282, u_muldiv_N281, u_muldiv_N280, net1883, u_muldiv_N279,
         u_muldiv_N278, u_muldiv_N277, u_muldiv_N276, u_muldiv_N275,
         u_muldiv_N274, u_muldiv_N273, u_muldiv_N272, u_muldiv_N271,
         u_muldiv_N270, u_muldiv_N269, u_muldiv_N268, u_muldiv_N267,
         u_muldiv_N266, u_muldiv_N265, u_muldiv_N263, u_muldiv_N246,
         u_decode_u_regfile_N965, n8300, u_decode_u_regfile_N928,
         u_decode_u_regfile_N945, u_decode_u_regfile_N980, n8332,
         u_decode_u_regfile_N943, u_decode_u_regfile_N979, u_muldiv_N260,
         u_decode_u_regfile_N942, u_decode_u_regfile_N951,
         u_decode_u_regfile_N993, u_muldiv_N237, u_decode_u_regfile_N956,
         u_csr_N3696, u_decode_N321, u_decode_u_regfile_N968,
         u_decode_u_regfile_N975, u_decode_u_regfile_N976,
         u_decode_u_regfile_N978, u_decode_u_regfile_N964,
         u_decode_u_regfile_N989, u_muldiv_N233, u_decode_u_regfile_N952,
         u_decode_u_regfile_N992, u_muldiv_N236, u_decode_u_regfile_N955,
         u_decode_u_regfile_N996, u_decode_u_regfile_N963,
         u_decode_u_regfile_N969, u_decode_u_regfile_N977,
         u_decode_u_regfile_N995, u_decode_u_regfile_N972,
         u_decode_u_regfile_N967, u_decode_u_regfile_N973,
         u_decode_u_regfile_N974, u_decode_u_regfile_N997,
         u_decode_u_regfile_N991, u_muldiv_N235, u_decode_u_regfile_N954,
         u_decode_u_regfile_N971, u_decode_u_regfile_N998,
         u_decode_u_regfile_N990, u_muldiv_N234, u_decode_u_regfile_N953,
         u_decode_u_regfile_N994, u_decode_u_regfile_N970,
         u_decode_u_regfile_N999, u_csr_csr_sr_r_12, u_csr_csr_sr_r_11,
         u_csr_csr_sr_r_8, u_csr_csr_sr_r_7, u_csr_csr_sr_r_5,
         u_csr_csr_sr_r_3, u_csr_csr_sr_r_1, u_csr_N3161, u_csr_N3162,
         u_csr_N3697, n8696, u_muldiv_N264, u_muldiv_div_busy_q, n8536, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, net1903, net1898, u_muldiv_N328, net1918,
         u_muldiv_N329, u_muldiv_N330, u_muldiv_N331, u_muldiv_N332,
         u_muldiv_N333, u_muldiv_N334, u_muldiv_N335, u_muldiv_N336,
         u_muldiv_N337, u_muldiv_N338, u_muldiv_N339, u_muldiv_N340,
         u_muldiv_N341, u_muldiv_N342, u_muldiv_N343, u_muldiv_N344, net1923,
         u_muldiv_N345, u_muldiv_N346, u_muldiv_N347, u_muldiv_N348,
         u_muldiv_N349, u_muldiv_N350, u_muldiv_N351, u_muldiv_N352,
         u_muldiv_N353, u_muldiv_N354, u_muldiv_N355, u_muldiv_N356,
         u_muldiv_N357, u_muldiv_N358, u_muldiv_N359, u_muldiv_N513, n8801,
         net2370, u_decode_N783, u_muldiv_mult_busy_q, u_csr_csr_satp_q_31_,
         n8554, u_mmu_dtlb_req_q, net1782, n8417, u_mmu_dtlb_entry_q_4, n8442,
         net1792, u_mmu_itlb_entry_q_3, u_mmu_itlb_entry_q_4, u_fetch_N157,
         u_fetch_fetch_page_fault_q, net2374, n8538, net2373, net2372, net2371,
         net2368, net2367, net2366, n8513, net2365, n8512, net2364, n8511,
         net2363, net2362, u_decode_N342, net2361, u_decode_N341, net2360,
         u_decode_N340, net2359, u_decode_N339, net2358, u_decode_N338,
         net2352, u_decode_N337, net2351, net2350, net2349, u_decode_N334,
         net2348, u_decode_N333, n8506, u_muldiv_N517, net2347, u_decode_N332,
         n8507, u_muldiv_N516, net2346, u_decode_N331, n8508, u_muldiv_N515,
         net2345, n8509, u_muldiv_N514, net2344, u_decode_N329, n8510, net2343,
         net2342, net2341, net2340, net2339, net2337, net2336, u_decode_N792,
         opcode_instr_w_57, opcode_instr_w_56, opcode_instr_w_55,
         opcode_instr_w_51, opcode_instr_w_48, opcode_instr_w_46,
         opcode_instr_w_45, opcode_instr_w_41, opcode_instr_w_40,
         opcode_instr_w_39, opcode_instr_w_38, opcode_instr_w_37,
         opcode_instr_w_36, opcode_instr_w_35, opcode_instr_w_28,
         opcode_instr_w_26, opcode_instr_w_25, opcode_instr_w_24,
         opcode_instr_w_18, opcode_instr_w_17, opcode_instr_w_16,
         opcode_instr_w_1, u_decode_N791, u_decode_N775, u_decode_N774,
         u_decode_N788, u_decode_N780, u_decode_N769, u_decode_N762,
         u_decode_N756, u_decode_N744, u_decode_N787, u_decode_N768, n17098,
         u_decode_N761, u_decode_N741, u_decode_N789, n8887, u_decode_N781,
         u_decode_N770, u_decode_N740, u_decode_N785, u_decode_N778,
         u_decode_N773, u_decode_N767, u_decode_N738, u_decode_N784,
         u_decode_N777, u_decode_N772, u_decode_N766, u_decode_N760,
         u_decode_N771, u_decode_N765, u_lsu_N103, n8574, n8441, u_mmu_load_q,
         u_lsu_N230, n8647, n8302, n8330, n8336, n8338, u_lsu_N226, u_lsu_N227,
         u_lsu_N228, u_lsu_N229, n8540, n8541, n8542, u_lsu_N98, n8810,
         u_lsu_N231, n8954, n8498, n8496, n8495, n8494, u_lsu_N99, n4705,
         n8255, u_decode_N759, u_decode_N748, u_decode_N737, u_decode_N786,
         u_decode_N779, u_decode_N739, u_decode_N790, u_decode_N782,
         u_csr_N2391, net1878, n8835, n8499, n8537, net1867, net1872,
         u_csr_N3471, u_csr_writeback_en_q, u_csr_N2377, \u_csr_csr_mip_r[11] ,
         u_csr_csr_mip_r_9, u_csr_csr_mip_r_7, u_csr_csr_mip_r_5,
         u_csr_csr_mip_r_3, u_csr_csr_mip_r_1, \u_csr_csr_mip_q[11] ,
         u_csr_csr_mip_q_7, u_csr_csr_mip_q_5, u_csr_csr_mip_q_3,
         u_csr_csr_mip_q_1, \u_csr_csr_mie_r[11] , u_csr_csr_mie_r_9,
         u_csr_csr_mie_r_7, u_csr_csr_mie_r_5, u_csr_csr_mie_r_3,
         u_csr_csr_mie_r_1, \u_csr_csr_mie_q[11] , u_csr_csr_mie_q_9,
         u_csr_csr_mie_q_7, u_csr_csr_mie_q_5, u_csr_csr_mie_q_3,
         u_csr_csr_mie_q_1, u_csr_N2395, u_csr_csr_sr_q_22, u_csr_N2394,
         u_csr_csr_sr_q_21, u_csr_N2393, u_csr_csr_sr_q_20, u_csr_N2392,
         u_csr_csr_sr_q_19, u_csr_N2390, u_csr_N2389, u_csr_N2388, u_csr_N2387,
         u_csr_N2386, u_csr_N2383, u_csr_N2382, u_csr_N2379, u_csr_N2375,
         u_csr_N2373, u_decode_N764, u_decode_N736, u_decode_N758,
         u_decode_N746, u_decode_N745, u_decode_N757, u_decode_valid_q,
         u_decode_N180, u_csr_csr_sr_q_31, u_csr_csr_sr_q_30,
         u_csr_csr_sr_q_29, u_csr_csr_sr_q_28, u_csr_csr_sr_q_27,
         u_csr_csr_sr_q_26, u_csr_csr_sr_q_25, u_csr_csr_sr_q_24,
         u_csr_csr_sr_q_23, n8504, u_mmu_dtlb_valid_q, n8505,
         u_mmu_itlb_valid_q, u_decode_N755, n8955, u_decode_N754,
         u_decode_N753, u_decode_N752, u_decode_N751, u_decode_N750,
         u_decode_N749, u_decode_N747, u_decode_N743, u_decode_N742,
         u_exec_N242, u_exec_N241, u_exec_N240, u_exec_N239, u_exec_N238,
         u_decode_N793, u_decode_N776, u_csr_N3472, net2415, net2416, n8521,
         u_muldiv_div_inst_q, u_csr_csr_scause_r_31, u_csr_csr_scause_q_31,
         u_csr_csr_mcause_r_31, u_csr_csr_mcause_q_31, u_csr_N3676, net2292,
         net2391, u_decode_N301, u_csr_N3694, net2315, net2414, u_decode_N319,
         u_csr_N3693, net2314, net2413, u_decode_N318, u_csr_N3692, net2313,
         net2412, u_decode_N317, u_csr_N3665, n8848, net2281, net2380,
         u_decode_N290, u_csr_N184, u_decode_u_regfile_N100,
         u_decode_u_regfile_N1025, u_decode_u_regfile_N1062,
         u_decode_u_regfile_N1099, u_decode_u_regfile_N1136,
         u_decode_u_regfile_N1173, u_decode_u_regfile_N1210,
         u_decode_u_regfile_N137, u_decode_u_regfile_N174,
         u_decode_u_regfile_N211, u_decode_u_regfile_N248,
         u_decode_u_regfile_N285, u_decode_u_regfile_N322,
         u_decode_u_regfile_N359, u_decode_u_regfile_N396,
         u_decode_u_regfile_N433, u_decode_u_regfile_N470,
         u_decode_u_regfile_N507, u_decode_u_regfile_N544,
         u_decode_u_regfile_N581, u_decode_u_regfile_N618,
         u_decode_u_regfile_N655, u_decode_u_regfile_N692,
         u_decode_u_regfile_N729, u_decode_u_regfile_N766,
         u_decode_u_regfile_N803, u_decode_u_regfile_N840,
         u_decode_u_regfile_N877, u_decode_u_regfile_N914, u_csr_N3666, n8836,
         net2282, net2381, u_decode_N291, u_decode_u_regfile_N101,
         u_decode_u_regfile_N1026, u_decode_u_regfile_N1063,
         u_decode_u_regfile_N1100, u_decode_u_regfile_N1137,
         u_decode_u_regfile_N1174, u_decode_u_regfile_N1211,
         u_decode_u_regfile_N138, u_decode_u_regfile_N175,
         u_decode_u_regfile_N212, u_decode_u_regfile_N249,
         u_decode_u_regfile_N286, u_decode_u_regfile_N323,
         u_decode_u_regfile_N360, u_decode_u_regfile_N397,
         u_decode_u_regfile_N434, u_decode_u_regfile_N471,
         u_decode_u_regfile_N508, u_decode_u_regfile_N545,
         u_decode_u_regfile_N582, u_decode_u_regfile_N619,
         u_decode_u_regfile_N656, u_decode_u_regfile_N693,
         u_decode_u_regfile_N730, u_decode_u_regfile_N767,
         u_decode_u_regfile_N804, u_decode_u_regfile_N841,
         u_decode_u_regfile_N878, u_decode_u_regfile_N915, u_csr_N3667, n8845,
         net2283, net2382, u_decode_u_regfile_N102, u_decode_u_regfile_N1027,
         u_decode_u_regfile_N1064, u_decode_u_regfile_N1101,
         u_decode_u_regfile_N1138, u_decode_u_regfile_N1175,
         u_decode_u_regfile_N1212, u_decode_u_regfile_N139,
         u_decode_u_regfile_N176, u_decode_u_regfile_N213,
         u_decode_u_regfile_N250, u_decode_u_regfile_N287,
         u_decode_u_regfile_N324, u_decode_u_regfile_N361,
         u_decode_u_regfile_N398, u_decode_u_regfile_N435,
         u_decode_u_regfile_N472, u_decode_u_regfile_N509,
         u_decode_u_regfile_N546, u_decode_u_regfile_N583,
         u_decode_u_regfile_N620, u_decode_u_regfile_N657,
         u_decode_u_regfile_N694, u_decode_u_regfile_N731,
         u_decode_u_regfile_N768, u_decode_u_regfile_N805,
         u_decode_u_regfile_N842, u_decode_u_regfile_N879,
         u_decode_u_regfile_N916, u_csr_N3668, net2284, net2383,
         u_decode_u_regfile_N1028, u_decode_u_regfile_N103,
         u_decode_u_regfile_N1065, u_decode_u_regfile_N1102,
         u_decode_u_regfile_N1139, u_decode_u_regfile_N1176,
         u_decode_u_regfile_N1213, u_decode_u_regfile_N140,
         u_decode_u_regfile_N177, u_decode_u_regfile_N214,
         u_decode_u_regfile_N251, u_decode_u_regfile_N288,
         u_decode_u_regfile_N325, u_decode_u_regfile_N362,
         u_decode_u_regfile_N399, u_decode_u_regfile_N436,
         u_decode_u_regfile_N473, u_decode_u_regfile_N510,
         u_decode_u_regfile_N547, u_decode_u_regfile_N584,
         u_decode_u_regfile_N621, u_decode_u_regfile_N658,
         u_decode_u_regfile_N695, u_decode_u_regfile_N732,
         u_decode_u_regfile_N769, u_decode_u_regfile_N806,
         u_decode_u_regfile_N843, u_decode_u_regfile_N880,
         u_decode_u_regfile_N917, u_csr_N3669, net2285, net2384, u_decode_N294,
         u_decode_u_regfile_N1029, u_decode_u_regfile_N104,
         u_decode_u_regfile_N1066, u_decode_u_regfile_N1103,
         u_decode_u_regfile_N1140, u_decode_u_regfile_N1177,
         u_decode_u_regfile_N1214, u_decode_u_regfile_N141,
         u_decode_u_regfile_N178, u_decode_u_regfile_N215,
         u_decode_u_regfile_N252, u_decode_u_regfile_N289,
         u_decode_u_regfile_N326, u_decode_u_regfile_N363,
         u_decode_u_regfile_N400, u_decode_u_regfile_N437,
         u_decode_u_regfile_N474, u_decode_u_regfile_N511,
         u_decode_u_regfile_N548, u_decode_u_regfile_N585,
         u_decode_u_regfile_N622, u_decode_u_regfile_N659,
         u_decode_u_regfile_N696, u_decode_u_regfile_N733,
         u_decode_u_regfile_N770, u_decode_u_regfile_N807,
         u_decode_u_regfile_N844, u_decode_u_regfile_N881,
         u_decode_u_regfile_N918, u_csr_N3670, net2286, net2385, u_decode_N295,
         u_decode_u_regfile_N1030, u_decode_u_regfile_N105,
         u_decode_u_regfile_N1067, u_decode_u_regfile_N1104,
         u_decode_u_regfile_N1141, u_decode_u_regfile_N1178,
         u_decode_u_regfile_N1215, u_decode_u_regfile_N142,
         u_decode_u_regfile_N179, u_decode_u_regfile_N216,
         u_decode_u_regfile_N253, u_decode_u_regfile_N290,
         u_decode_u_regfile_N327, u_decode_u_regfile_N364,
         u_decode_u_regfile_N401, u_decode_u_regfile_N438,
         u_decode_u_regfile_N475, u_decode_u_regfile_N512,
         u_decode_u_regfile_N549, u_decode_u_regfile_N586,
         u_decode_u_regfile_N623, u_decode_u_regfile_N660,
         u_decode_u_regfile_N697, u_decode_u_regfile_N734,
         u_decode_u_regfile_N771, u_decode_u_regfile_N808,
         u_decode_u_regfile_N845, u_decode_u_regfile_N882,
         u_decode_u_regfile_N919, u_csr_N3671, net2287, net2386, u_decode_N296,
         u_csr_N3672, net2288, net2387, u_decode_N297, u_csr_N3673, net2289,
         net2388, u_decode_N298, u_csr_N3674, net2290, net2389, u_decode_N299,
         u_csr_N3675, net2291, net2390, u_decode_N300, u_csr_N3677, net2293,
         net2392, u_decode_N302, u_csr_N3678, net2294, net2393, u_decode_N303,
         u_csr_N3679, net2295, net2394, u_decode_N304, n17100, u_mmu_N241,
         u_csr_N3680, net2296, net2395, u_mmu_N242, u_csr_N3681, net2302,
         net2401, u_decode_N306, u_csr_N3682, net2303, net2402, u_decode_N307,
         u_csr_N3683, net2304, net2403, u_decode_N308, u_csr_N3684, net2305,
         net2404, u_decode_N309, u_csr_N3685, net2306, net2405, u_decode_N310,
         u_csr_N3686, net2307, net2406, u_decode_N311, u_csr_N3687, net2308,
         net2407, u_decode_N312, u_csr_N3688, net2309, net2408, u_decode_N313,
         u_csr_N3689, net2310, net2409, u_decode_N314, u_csr_N3690, net2311,
         net2410, u_decode_N315, u_csr_N3691, net2312, net2411, u_decode_N316,
         n8502, n8501, n8551, n8440, n8439, u_decode_u_regfile_N1016,
         u_decode_u_regfile_N1053, u_decode_u_regfile_N1090,
         u_decode_u_regfile_N1127, u_decode_u_regfile_N1164,
         u_decode_u_regfile_N1201, u_decode_u_regfile_N1238,
         u_decode_u_regfile_N128, u_decode_u_regfile_N165,
         u_decode_u_regfile_N202, u_decode_u_regfile_N239,
         u_decode_u_regfile_N276, u_decode_u_regfile_N313,
         u_decode_u_regfile_N350, u_decode_u_regfile_N387,
         u_decode_u_regfile_N424, u_decode_u_regfile_N461,
         u_decode_u_regfile_N498, u_decode_u_regfile_N535,
         u_decode_u_regfile_N572, u_decode_u_regfile_N609,
         u_decode_u_regfile_N646, u_decode_u_regfile_N683,
         u_decode_u_regfile_N720, u_decode_u_regfile_N757,
         u_decode_u_regfile_N794, u_decode_u_regfile_N831,
         u_decode_u_regfile_N868, u_decode_u_regfile_N905, n8500, u_csr_N3695,
         net2316, u_decode_u_regfile_N1003, u_decode_u_regfile_N1040,
         u_decode_u_regfile_N1077, u_decode_u_regfile_N1114,
         u_decode_u_regfile_N115, u_decode_u_regfile_N1151,
         u_decode_u_regfile_N1188, u_decode_u_regfile_N1225,
         u_decode_u_regfile_N152, u_decode_u_regfile_N189,
         u_decode_u_regfile_N226, u_decode_u_regfile_N263,
         u_decode_u_regfile_N300, u_decode_u_regfile_N337,
         u_decode_u_regfile_N374, u_decode_u_regfile_N411,
         u_decode_u_regfile_N448, u_decode_u_regfile_N485,
         u_decode_u_regfile_N522, u_decode_u_regfile_N559,
         u_decode_u_regfile_N596, u_decode_u_regfile_N633,
         u_decode_u_regfile_N670, u_decode_u_regfile_N707,
         u_decode_u_regfile_N744, u_decode_u_regfile_N781,
         u_decode_u_regfile_N818, u_decode_u_regfile_N855,
         u_decode_u_regfile_N892, u_muldiv_N243, u_decode_u_regfile_N1036,
         u_decode_u_regfile_N1073, u_decode_u_regfile_N111,
         u_decode_u_regfile_N1110, u_decode_u_regfile_N1147,
         u_decode_u_regfile_N1184, u_decode_u_regfile_N1221,
         u_decode_u_regfile_N148, u_decode_u_regfile_N185,
         u_decode_u_regfile_N222, u_decode_u_regfile_N259,
         u_decode_u_regfile_N296, u_decode_u_regfile_N333,
         u_decode_u_regfile_N370, u_decode_u_regfile_N407,
         u_decode_u_regfile_N444, u_decode_u_regfile_N481,
         u_decode_u_regfile_N518, u_decode_u_regfile_N555,
         u_decode_u_regfile_N592, u_decode_u_regfile_N629,
         u_decode_u_regfile_N666, u_decode_u_regfile_N703,
         u_decode_u_regfile_N740, u_decode_u_regfile_N777,
         u_decode_u_regfile_N814, u_decode_u_regfile_N851,
         u_decode_u_regfile_N888, u_decode_u_regfile_N925,
         u_decode_u_regfile_N962, n8310, u_mmu_N246, u_muldiv_N251,
         u_decode_u_regfile_N1007, u_decode_u_regfile_N1044,
         u_decode_u_regfile_N1081, u_decode_u_regfile_N1118,
         u_decode_u_regfile_N1155, u_decode_u_regfile_N119,
         u_decode_u_regfile_N1192, u_decode_u_regfile_N1229,
         u_decode_u_regfile_N156, u_decode_u_regfile_N193,
         u_decode_u_regfile_N230, u_decode_u_regfile_N267,
         u_decode_u_regfile_N304, u_decode_u_regfile_N341,
         u_decode_u_regfile_N378, u_decode_u_regfile_N415,
         u_decode_u_regfile_N452, u_decode_u_regfile_N489,
         u_decode_u_regfile_N526, u_decode_u_regfile_N563,
         u_decode_u_regfile_N600, u_decode_u_regfile_N637,
         u_decode_u_regfile_N674, u_decode_u_regfile_N711,
         u_decode_u_regfile_N748, u_decode_u_regfile_N785,
         u_decode_u_regfile_N822, u_decode_u_regfile_N859,
         u_decode_u_regfile_N896, u_decode_u_regfile_N933, u_muldiv_N238,
         u_decode_u_regfile_N1031, u_decode_u_regfile_N106,
         u_decode_u_regfile_N1068, u_decode_u_regfile_N1105,
         u_decode_u_regfile_N1142, u_decode_u_regfile_N1179,
         u_decode_u_regfile_N1216, u_decode_u_regfile_N143,
         u_decode_u_regfile_N180, u_decode_u_regfile_N217,
         u_decode_u_regfile_N254, u_decode_u_regfile_N291,
         u_decode_u_regfile_N328, u_decode_u_regfile_N365,
         u_decode_u_regfile_N402, u_decode_u_regfile_N439,
         u_decode_u_regfile_N476, u_decode_u_regfile_N513,
         u_decode_u_regfile_N550, u_decode_u_regfile_N587,
         u_decode_u_regfile_N624, u_decode_u_regfile_N661,
         u_decode_u_regfile_N698, u_decode_u_regfile_N735,
         u_decode_u_regfile_N772, u_decode_u_regfile_N809,
         u_decode_u_regfile_N846, u_decode_u_regfile_N883,
         u_decode_u_regfile_N920, u_decode_u_regfile_N957, u_lsu_N200,
         u_lsu_N196, u_muldiv_N242, u_decode_u_regfile_N1035,
         u_decode_u_regfile_N1072, u_decode_u_regfile_N110,
         u_decode_u_regfile_N1109, u_decode_u_regfile_N1146,
         u_decode_u_regfile_N1183, u_decode_u_regfile_N1220,
         u_decode_u_regfile_N147, u_decode_u_regfile_N184,
         u_decode_u_regfile_N221, u_decode_u_regfile_N258,
         u_decode_u_regfile_N295, u_decode_u_regfile_N332,
         u_decode_u_regfile_N369, u_decode_u_regfile_N406,
         u_decode_u_regfile_N443, u_decode_u_regfile_N480,
         u_decode_u_regfile_N517, u_decode_u_regfile_N554,
         u_decode_u_regfile_N591, u_decode_u_regfile_N628,
         u_decode_u_regfile_N665, u_decode_u_regfile_N702,
         u_decode_u_regfile_N739, u_decode_u_regfile_N776,
         u_decode_u_regfile_N813, u_decode_u_regfile_N850,
         u_decode_u_regfile_N887, u_decode_u_regfile_N924,
         u_decode_u_regfile_N961, u_lsu_N204, n8314, u_mmu_N247, u_muldiv_N252,
         u_decode_u_regfile_N1008, u_decode_u_regfile_N1045,
         u_decode_u_regfile_N1082, u_decode_u_regfile_N1119,
         u_decode_u_regfile_N1156, u_decode_u_regfile_N1193,
         u_decode_u_regfile_N120, u_decode_u_regfile_N1230,
         u_decode_u_regfile_N157, u_decode_u_regfile_N194,
         u_decode_u_regfile_N231, u_decode_u_regfile_N268,
         u_decode_u_regfile_N305, u_decode_u_regfile_N342,
         u_decode_u_regfile_N379, u_decode_u_regfile_N416,
         u_decode_u_regfile_N453, u_decode_u_regfile_N490,
         u_decode_u_regfile_N527, u_decode_u_regfile_N564,
         u_decode_u_regfile_N601, u_decode_u_regfile_N638,
         u_decode_u_regfile_N675, u_decode_u_regfile_N712,
         u_decode_u_regfile_N749, u_decode_u_regfile_N786,
         u_decode_u_regfile_N823, u_decode_u_regfile_N860,
         u_decode_u_regfile_N897, u_decode_u_regfile_N934, u_lsu_N197,
         u_lsu_N205, u_lsu_N213, net1847, u_muldiv_N241,
         u_decode_u_regfile_N1034, u_decode_u_regfile_N1071,
         u_decode_u_regfile_N109, u_decode_u_regfile_N1108,
         u_decode_u_regfile_N1145, u_decode_u_regfile_N1182,
         u_decode_u_regfile_N1219, u_decode_u_regfile_N146,
         u_decode_u_regfile_N183, u_decode_u_regfile_N220,
         u_decode_u_regfile_N257, u_decode_u_regfile_N294,
         u_decode_u_regfile_N331, u_decode_u_regfile_N368,
         u_decode_u_regfile_N405, u_decode_u_regfile_N442,
         u_decode_u_regfile_N479, u_decode_u_regfile_N516,
         u_decode_u_regfile_N553, u_decode_u_regfile_N590,
         u_decode_u_regfile_N627, u_decode_u_regfile_N664,
         u_decode_u_regfile_N701, u_decode_u_regfile_N738,
         u_decode_u_regfile_N775, u_decode_u_regfile_N812,
         u_decode_u_regfile_N849, u_decode_u_regfile_N886,
         u_decode_u_regfile_N923, u_decode_u_regfile_N960, n8320, n8438, n8437,
         u_muldiv_N255, u_decode_u_regfile_N1011, u_decode_u_regfile_N1048,
         u_decode_u_regfile_N1085, u_decode_u_regfile_N1122,
         u_decode_u_regfile_N1159, u_decode_u_regfile_N1196,
         u_decode_u_regfile_N123, u_decode_u_regfile_N1233,
         u_decode_u_regfile_N160, u_decode_u_regfile_N197,
         u_decode_u_regfile_N234, u_decode_u_regfile_N271,
         u_decode_u_regfile_N308, u_decode_u_regfile_N345,
         u_decode_u_regfile_N382, u_decode_u_regfile_N419,
         u_decode_u_regfile_N456, u_decode_u_regfile_N493,
         u_decode_u_regfile_N530, u_decode_u_regfile_N567,
         u_decode_u_regfile_N604, u_decode_u_regfile_N641,
         u_decode_u_regfile_N678, u_decode_u_regfile_N715,
         u_decode_u_regfile_N752, u_decode_u_regfile_N789,
         u_decode_u_regfile_N826, u_decode_u_regfile_N863,
         u_decode_u_regfile_N900, u_decode_u_regfile_N937, n8318, n8436, n8435,
         u_muldiv_N254, u_decode_u_regfile_N1010, u_decode_u_regfile_N1047,
         u_decode_u_regfile_N1084, u_decode_u_regfile_N1121,
         u_decode_u_regfile_N1158, u_decode_u_regfile_N1195,
         u_decode_u_regfile_N122, u_decode_u_regfile_N1232,
         u_decode_u_regfile_N159, u_decode_u_regfile_N196,
         u_decode_u_regfile_N233, u_decode_u_regfile_N270,
         u_decode_u_regfile_N307, u_decode_u_regfile_N344,
         u_decode_u_regfile_N381, u_decode_u_regfile_N418,
         u_decode_u_regfile_N455, u_decode_u_regfile_N492,
         u_decode_u_regfile_N529, u_decode_u_regfile_N566,
         u_decode_u_regfile_N603, u_decode_u_regfile_N640,
         u_decode_u_regfile_N677, u_decode_u_regfile_N714,
         u_decode_u_regfile_N751, u_decode_u_regfile_N788,
         u_decode_u_regfile_N825, u_decode_u_regfile_N862,
         u_decode_u_regfile_N899, u_decode_u_regfile_N936, u_lsu_N216, n8304,
         u_mmu_N243, u_muldiv_N248, u_decode_u_regfile_N1004,
         u_decode_u_regfile_N1041, u_decode_u_regfile_N1078,
         u_decode_u_regfile_N1115, u_decode_u_regfile_N1152,
         u_decode_u_regfile_N116, u_decode_u_regfile_N1189,
         u_decode_u_regfile_N1226, u_decode_u_regfile_N153,
         u_decode_u_regfile_N190, u_decode_u_regfile_N227,
         u_decode_u_regfile_N264, u_decode_u_regfile_N301,
         u_decode_u_regfile_N338, u_decode_u_regfile_N375,
         u_decode_u_regfile_N412, u_decode_u_regfile_N449,
         u_decode_u_regfile_N486, u_decode_u_regfile_N523,
         u_decode_u_regfile_N560, u_decode_u_regfile_N597,
         u_decode_u_regfile_N634, u_decode_u_regfile_N671,
         u_decode_u_regfile_N708, u_decode_u_regfile_N745,
         u_decode_u_regfile_N782, u_decode_u_regfile_N819,
         u_decode_u_regfile_N856, u_decode_u_regfile_N893,
         u_decode_u_regfile_N930, n8316, n8434, u_mmu_N248, u_muldiv_N253,
         u_decode_u_regfile_N1009, u_decode_u_regfile_N1046,
         u_decode_u_regfile_N1083, u_decode_u_regfile_N1120,
         u_decode_u_regfile_N1157, u_decode_u_regfile_N1194,
         u_decode_u_regfile_N121, u_decode_u_regfile_N1231,
         u_decode_u_regfile_N158, u_decode_u_regfile_N195,
         u_decode_u_regfile_N232, u_decode_u_regfile_N269,
         u_decode_u_regfile_N306, u_decode_u_regfile_N343,
         u_decode_u_regfile_N380, u_decode_u_regfile_N417,
         u_decode_u_regfile_N454, u_decode_u_regfile_N491,
         u_decode_u_regfile_N528, u_decode_u_regfile_N565,
         u_decode_u_regfile_N602, u_decode_u_regfile_N639,
         u_decode_u_regfile_N676, u_decode_u_regfile_N713,
         u_decode_u_regfile_N750, u_decode_u_regfile_N787,
         u_decode_u_regfile_N824, u_decode_u_regfile_N861,
         u_decode_u_regfile_N898, u_decode_u_regfile_N935, u_muldiv_N239,
         u_decode_u_regfile_N1032, u_decode_u_regfile_N1069,
         u_decode_u_regfile_N107, u_decode_u_regfile_N1106,
         u_decode_u_regfile_N1143, u_decode_u_regfile_N1180,
         u_decode_u_regfile_N1217, u_decode_u_regfile_N144,
         u_decode_u_regfile_N181, u_decode_u_regfile_N218,
         u_decode_u_regfile_N255, u_decode_u_regfile_N292,
         u_decode_u_regfile_N329, u_decode_u_regfile_N366,
         u_decode_u_regfile_N403, u_decode_u_regfile_N440,
         u_decode_u_regfile_N477, u_decode_u_regfile_N514,
         u_decode_u_regfile_N551, u_decode_u_regfile_N588,
         u_decode_u_regfile_N625, u_decode_u_regfile_N662,
         u_decode_u_regfile_N699, u_decode_u_regfile_N736,
         u_decode_u_regfile_N773, u_decode_u_regfile_N810,
         u_decode_u_regfile_N847, u_decode_u_regfile_N884,
         u_decode_u_regfile_N921, u_decode_u_regfile_N958, u_lsu_N201,
         u_lsu_N209, u_lsu_N217, u_lsu_N225, n8326, n8433, n8432,
         u_muldiv_N258, u_decode_u_regfile_N1014, u_decode_u_regfile_N1051,
         u_decode_u_regfile_N1088, u_decode_u_regfile_N1125,
         u_decode_u_regfile_N1162, u_decode_u_regfile_N1199,
         u_decode_u_regfile_N1236, u_decode_u_regfile_N126,
         u_decode_u_regfile_N163, u_decode_u_regfile_N200,
         u_decode_u_regfile_N237, u_decode_u_regfile_N274,
         u_decode_u_regfile_N311, u_decode_u_regfile_N348,
         u_decode_u_regfile_N385, u_decode_u_regfile_N422,
         u_decode_u_regfile_N459, u_decode_u_regfile_N496,
         u_decode_u_regfile_N533, u_decode_u_regfile_N570,
         u_decode_u_regfile_N607, u_decode_u_regfile_N644,
         u_decode_u_regfile_N681, u_decode_u_regfile_N718,
         u_decode_u_regfile_N755, u_decode_u_regfile_N792,
         u_decode_u_regfile_N829, u_decode_u_regfile_N866,
         u_decode_u_regfile_N903, u_decode_u_regfile_N940, u_lsu_N220, n8308,
         n17102, u_mmu_N245, u_muldiv_N250, u_decode_u_regfile_N1006,
         u_decode_u_regfile_N1043, u_decode_u_regfile_N1080,
         u_decode_u_regfile_N1117, u_decode_u_regfile_N1154,
         u_decode_u_regfile_N118, u_decode_u_regfile_N1191,
         u_decode_u_regfile_N1228, u_decode_u_regfile_N155,
         u_decode_u_regfile_N192, u_decode_u_regfile_N229,
         u_decode_u_regfile_N266, u_decode_u_regfile_N303,
         u_decode_u_regfile_N340, u_decode_u_regfile_N377,
         u_decode_u_regfile_N414, u_decode_u_regfile_N451,
         u_decode_u_regfile_N488, u_decode_u_regfile_N525,
         u_decode_u_regfile_N562, u_decode_u_regfile_N599,
         u_decode_u_regfile_N636, u_decode_u_regfile_N673,
         u_decode_u_regfile_N710, u_decode_u_regfile_N747,
         u_decode_u_regfile_N784, u_decode_u_regfile_N821,
         u_decode_u_regfile_N858, u_decode_u_regfile_N895,
         u_decode_u_regfile_N932, u_lsu_N212, n8296, u_mmu_N239, u_muldiv_N244,
         u_decode_u_regfile_N1000, u_decode_u_regfile_N1037,
         u_decode_u_regfile_N1074, u_decode_u_regfile_N1111,
         u_decode_u_regfile_N112, u_decode_u_regfile_N1148,
         u_decode_u_regfile_N1185, u_decode_u_regfile_N1222,
         u_decode_u_regfile_N149, u_decode_u_regfile_N186,
         u_decode_u_regfile_N223, u_decode_u_regfile_N260,
         u_decode_u_regfile_N297, u_decode_u_regfile_N334,
         u_decode_u_regfile_N371, u_decode_u_regfile_N408,
         u_decode_u_regfile_N445, u_decode_u_regfile_N482,
         u_decode_u_regfile_N519, u_decode_u_regfile_N556,
         u_decode_u_regfile_N593, u_decode_u_regfile_N630,
         u_decode_u_regfile_N667, u_decode_u_regfile_N704,
         u_decode_u_regfile_N741, u_decode_u_regfile_N778,
         u_decode_u_regfile_N815, u_decode_u_regfile_N852,
         u_decode_u_regfile_N889, u_decode_u_regfile_N926, u_muldiv_N240,
         u_decode_u_regfile_N1033, u_decode_u_regfile_N1070,
         u_decode_u_regfile_N108, u_decode_u_regfile_N1107,
         u_decode_u_regfile_N1144, u_decode_u_regfile_N1181,
         u_decode_u_regfile_N1218, u_decode_u_regfile_N145,
         u_decode_u_regfile_N182, u_decode_u_regfile_N219,
         u_decode_u_regfile_N256, u_decode_u_regfile_N293,
         u_decode_u_regfile_N330, u_decode_u_regfile_N367,
         u_decode_u_regfile_N404, u_decode_u_regfile_N441,
         u_decode_u_regfile_N478, u_decode_u_regfile_N515,
         u_decode_u_regfile_N552, u_decode_u_regfile_N589,
         u_decode_u_regfile_N626, u_decode_u_regfile_N663,
         u_decode_u_regfile_N700, u_decode_u_regfile_N737,
         u_decode_u_regfile_N774, u_decode_u_regfile_N811,
         u_decode_u_regfile_N848, u_decode_u_regfile_N885,
         u_decode_u_regfile_N922, u_decode_u_regfile_N959, u_lsu_N198,
         u_lsu_N206, u_lsu_N214, u_lsu_N195, u_lsu_N203, n8298, n16237,
         u_mmu_N240, u_muldiv_N245, u_decode_u_regfile_N1001,
         u_decode_u_regfile_N1038, u_decode_u_regfile_N1075,
         u_decode_u_regfile_N1112, u_decode_u_regfile_N113,
         u_decode_u_regfile_N1149, u_decode_u_regfile_N1186,
         u_decode_u_regfile_N1223, u_decode_u_regfile_N150,
         u_decode_u_regfile_N187, u_decode_u_regfile_N224,
         u_decode_u_regfile_N261, u_decode_u_regfile_N298,
         u_decode_u_regfile_N335, u_decode_u_regfile_N372,
         u_decode_u_regfile_N409, u_decode_u_regfile_N446,
         u_decode_u_regfile_N483, u_decode_u_regfile_N520,
         u_decode_u_regfile_N557, u_decode_u_regfile_N594,
         u_decode_u_regfile_N631, u_decode_u_regfile_N668,
         u_decode_u_regfile_N705, u_decode_u_regfile_N742,
         u_decode_u_regfile_N779, u_decode_u_regfile_N816,
         u_decode_u_regfile_N853, u_decode_u_regfile_N890,
         u_decode_u_regfile_N927, n8328, u_muldiv_N259,
         u_decode_u_regfile_N1015, u_decode_u_regfile_N1052,
         u_decode_u_regfile_N1089, u_decode_u_regfile_N1126,
         u_decode_u_regfile_N1163, u_decode_u_regfile_N1200,
         u_decode_u_regfile_N1237, u_decode_u_regfile_N127,
         u_decode_u_regfile_N164, u_decode_u_regfile_N201,
         u_decode_u_regfile_N238, u_decode_u_regfile_N275,
         u_decode_u_regfile_N312, u_decode_u_regfile_N349,
         u_decode_u_regfile_N386, u_decode_u_regfile_N423,
         u_decode_u_regfile_N460, u_decode_u_regfile_N497,
         u_decode_u_regfile_N534, u_decode_u_regfile_N571,
         u_decode_u_regfile_N608, u_decode_u_regfile_N645,
         u_decode_u_regfile_N682, u_decode_u_regfile_N719,
         u_decode_u_regfile_N756, u_decode_u_regfile_N793,
         u_decode_u_regfile_N830, u_decode_u_regfile_N867,
         u_decode_u_regfile_N904, u_decode_u_regfile_N941, u_lsu_N221, n8324,
         n8431, n8430, u_muldiv_N257, u_decode_u_regfile_N1013,
         u_decode_u_regfile_N1050, u_decode_u_regfile_N1087,
         u_decode_u_regfile_N1124, u_decode_u_regfile_N1161,
         u_decode_u_regfile_N1198, u_decode_u_regfile_N1235,
         u_decode_u_regfile_N125, u_decode_u_regfile_N162,
         u_decode_u_regfile_N199, u_decode_u_regfile_N236,
         u_decode_u_regfile_N273, u_decode_u_regfile_N310,
         u_decode_u_regfile_N347, u_decode_u_regfile_N384,
         u_decode_u_regfile_N421, u_decode_u_regfile_N458,
         u_decode_u_regfile_N495, u_decode_u_regfile_N532,
         u_decode_u_regfile_N569, u_decode_u_regfile_N606,
         u_decode_u_regfile_N643, u_decode_u_regfile_N680,
         u_decode_u_regfile_N717, u_decode_u_regfile_N754,
         u_decode_u_regfile_N791, u_decode_u_regfile_N828,
         u_decode_u_regfile_N865, u_decode_u_regfile_N902,
         u_decode_u_regfile_N939, u_lsu_N219, n8322, n8429, n8428,
         u_muldiv_N256, u_decode_u_regfile_N1012, u_decode_u_regfile_N1049,
         u_decode_u_regfile_N1086, u_decode_u_regfile_N1123,
         u_decode_u_regfile_N1160, u_decode_u_regfile_N1197,
         u_decode_u_regfile_N1234, u_decode_u_regfile_N124,
         u_decode_u_regfile_N161, u_decode_u_regfile_N198,
         u_decode_u_regfile_N235, u_decode_u_regfile_N272,
         u_decode_u_regfile_N309, u_decode_u_regfile_N346,
         u_decode_u_regfile_N383, u_decode_u_regfile_N420,
         u_decode_u_regfile_N457, u_decode_u_regfile_N494,
         u_decode_u_regfile_N531, u_decode_u_regfile_N568,
         u_decode_u_regfile_N605, u_decode_u_regfile_N642,
         u_decode_u_regfile_N679, u_decode_u_regfile_N716,
         u_decode_u_regfile_N753, u_decode_u_regfile_N790,
         u_decode_u_regfile_N827, u_decode_u_regfile_N864,
         u_decode_u_regfile_N901, u_decode_u_regfile_N938, n8306, u_mmu_N244,
         u_muldiv_N249, u_decode_u_regfile_N1005, u_decode_u_regfile_N1042,
         u_decode_u_regfile_N1079, u_decode_u_regfile_N1116,
         u_decode_u_regfile_N1153, u_decode_u_regfile_N117,
         u_decode_u_regfile_N1190, u_decode_u_regfile_N1227,
         u_decode_u_regfile_N154, u_decode_u_regfile_N191,
         u_decode_u_regfile_N228, u_decode_u_regfile_N265,
         u_decode_u_regfile_N302, u_decode_u_regfile_N339,
         u_decode_u_regfile_N376, u_decode_u_regfile_N413,
         u_decode_u_regfile_N450, u_decode_u_regfile_N487,
         u_decode_u_regfile_N524, u_decode_u_regfile_N561,
         u_decode_u_regfile_N598, u_decode_u_regfile_N635,
         u_decode_u_regfile_N672, u_decode_u_regfile_N709,
         u_decode_u_regfile_N746, u_decode_u_regfile_N783,
         u_decode_u_regfile_N820, u_decode_u_regfile_N857,
         u_decode_u_regfile_N894, u_decode_u_regfile_N931, u_muldiv_N327,
         u_muldiv_N326, u_lsu_N211, net2317, u_decode_u_regfile_N1019,
         u_decode_u_regfile_N1056, u_decode_u_regfile_N1093,
         u_decode_u_regfile_N1130, u_decode_u_regfile_N1167,
         u_decode_u_regfile_N1204, u_decode_u_regfile_N1241,
         u_decode_u_regfile_N131, u_decode_u_regfile_N168,
         u_decode_u_regfile_N205, u_decode_u_regfile_N242,
         u_decode_u_regfile_N279, u_decode_u_regfile_N316,
         u_decode_u_regfile_N353, u_decode_u_regfile_N390,
         u_decode_u_regfile_N427, u_decode_u_regfile_N464,
         u_decode_u_regfile_N501, u_decode_u_regfile_N538,
         u_decode_u_regfile_N575, u_decode_u_regfile_N612,
         u_decode_u_regfile_N649, u_decode_u_regfile_N686,
         u_decode_u_regfile_N723, u_decode_u_regfile_N760,
         u_decode_u_regfile_N797, u_decode_u_regfile_N834,
         u_decode_u_regfile_N871, u_decode_u_regfile_N908, u_lsu_N199,
         u_lsu_N207, u_lsu_N215, u_lsu_N194, u_lsu_N202, u_lsu_N210,
         u_lsu_N218, u_lsu_N222, u_decode_u_regfile_N1018,
         u_decode_u_regfile_N1055, u_decode_u_regfile_N1092,
         u_decode_u_regfile_N1129, u_decode_u_regfile_N1166,
         u_decode_u_regfile_N1203, u_decode_u_regfile_N1240,
         u_decode_u_regfile_N130, u_decode_u_regfile_N167,
         u_decode_u_regfile_N204, u_decode_u_regfile_N241,
         u_decode_u_regfile_N278, u_decode_u_regfile_N315,
         u_decode_u_regfile_N352, u_decode_u_regfile_N389,
         u_decode_u_regfile_N426, u_decode_u_regfile_N463,
         u_decode_u_regfile_N500, u_decode_u_regfile_N537,
         u_decode_u_regfile_N574, u_decode_u_regfile_N611,
         u_decode_u_regfile_N648, u_decode_u_regfile_N685,
         u_decode_u_regfile_N722, u_decode_u_regfile_N759,
         u_decode_u_regfile_N796, u_decode_u_regfile_N833,
         u_decode_u_regfile_N870, u_decode_u_regfile_N907,
         u_decode_u_regfile_N1017, u_decode_u_regfile_N1054,
         u_decode_u_regfile_N1091, u_decode_u_regfile_N1128,
         u_decode_u_regfile_N1165, u_decode_u_regfile_N1202,
         u_decode_u_regfile_N1239, u_decode_u_regfile_N129,
         u_decode_u_regfile_N166, u_decode_u_regfile_N203,
         u_decode_u_regfile_N240, u_decode_u_regfile_N277,
         u_decode_u_regfile_N314, u_decode_u_regfile_N351,
         u_decode_u_regfile_N388, u_decode_u_regfile_N425,
         u_decode_u_regfile_N462, u_decode_u_regfile_N499,
         u_decode_u_regfile_N536, u_decode_u_regfile_N573,
         u_decode_u_regfile_N610, u_decode_u_regfile_N647,
         u_decode_u_regfile_N684, u_decode_u_regfile_N721,
         u_decode_u_regfile_N758, u_decode_u_regfile_N795,
         u_decode_u_regfile_N832, u_decode_u_regfile_N869,
         u_decode_u_regfile_N906, u_lsu_N223, u_muldiv_N325, u_muldiv_N324,
         u_muldiv_N323, u_muldiv_N322, u_muldiv_N321, u_muldiv_N320,
         u_muldiv_N319, u_muldiv_N318, u_muldiv_N317, u_muldiv_N316,
         u_muldiv_N315, u_muldiv_N314, u_muldiv_N313, u_muldiv_N312,
         u_muldiv_N261, u_decode_u_regfile_N1002, u_decode_u_regfile_N1039,
         u_decode_u_regfile_N1076, u_decode_u_regfile_N1113,
         u_decode_u_regfile_N114, u_decode_u_regfile_N1150,
         u_decode_u_regfile_N1187, u_decode_u_regfile_N1224,
         u_decode_u_regfile_N151, u_decode_u_regfile_N188,
         u_decode_u_regfile_N225, u_decode_u_regfile_N262,
         u_decode_u_regfile_N299, u_decode_u_regfile_N336,
         u_decode_u_regfile_N373, u_decode_u_regfile_N410,
         u_decode_u_regfile_N447, u_decode_u_regfile_N484,
         u_decode_u_regfile_N521, u_decode_u_regfile_N558,
         u_decode_u_regfile_N595, u_decode_u_regfile_N632,
         u_decode_u_regfile_N669, u_decode_u_regfile_N706,
         u_decode_u_regfile_N743, u_decode_u_regfile_N780,
         u_decode_u_regfile_N817, u_decode_u_regfile_N854,
         u_decode_u_regfile_N891, u_lsu_N208, u_lsu_N224, n8553, n8427, n8426,
         n8560, n8425, n8424, n8423, U1_U7_Z_2, U1_U7_Z_3, U1_U7_Z_4,
         U1_U7_Z_5, U1_U7_Z_6, U1_U7_Z_7, U1_U7_Z_8, U1_U7_Z_9, U1_U7_Z_10,
         U1_U7_Z_11, U1_U6_Z_12, U1_U6_Z_13, U1_U6_Z_14, U1_U6_Z_15,
         U1_U6_Z_16, U1_U6_Z_17, U1_U6_Z_18, U1_U6_Z_19, U1_U6_Z_20,
         U1_U6_Z_21, U1_U6_Z_22, U1_U6_Z_23, U1_U6_Z_24, U1_U6_Z_25,
         U1_U6_Z_26, U1_U6_Z_27, U1_U6_Z_28, U1_U6_Z_29, U1_U6_Z_30,
         U1_U6_Z_31, n8559, n17208, n17209, n17210, n17211, n17212, n17213,
         n17214, n17215, n17216, n17217, n17218, n17219, n17220, n17221,
         n17222, n17223, net1857, n17224, net1862, n17225, n17226, n17227,
         n17228, n17229, n17230, n17231, n17232, n17233, n17234, n17235,
         n17236, n17237, n17238, n17239, n17240, n17241, n17242, n17243,
         n17244, n17245, n17246, n17247, n17248, n17249, n17250, n17251,
         n17252, n17253, n17254, n17255, n17256, n17257, n17258, n17259,
         n17260, n17261, n17262, n17263, n17264, n17265, n17266, n17267,
         n17268, n17269, n17270, n17271, n17272, n17273, n17274, n17275,
         n17276, n17277, n17278, n17279, n17280, n17281, n17282, n17283,
         n17284, n17285, n17286, n17287, n17288, n17289, n17290, n17291,
         n17292, n17293, n17294, n17295, n17296, n17297, n17298, n17299,
         n17300, n17301, n17302, n17303, n17304, n17305, n17306, n17307,
         n17308, n17309, n17310, n17311, n17312, n17313, n17314, n17315,
         u_muldiv_N529, u_muldiv_N528, u_muldiv_N530, u_muldiv_N531,
         u_muldiv_N527, u_muldiv_N532, u_muldiv_N523, u_muldiv_N524,
         u_muldiv_N525, u_muldiv_N522, u_muldiv_N526, u_muldiv_N521,
         u_muldiv_N538, u_muldiv_N545, u_muldiv_N546, u_muldiv_N548,
         u_muldiv_N534, u_muldiv_N533, u_muldiv_N539, u_muldiv_N547,
         u_muldiv_N542, u_muldiv_N537, u_muldiv_N543, u_muldiv_N544,
         u_muldiv_N541, u_muldiv_N540, u_muldiv_N549, u_muldiv_N550,
         u_muldiv_N535, u_muldiv_N536, u_muldiv_N552, u_muldiv_N551,
         u_decode_N292, n8518, n8516, n8517, n8519, n8514, n8515,
         u_decode_N763, u_decode_N330, u_decode_N293, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n48,
         n49, n50, n51, n52, n53, n54, n55, n179, n180, n215, n216, n226, n227,
         n229, n255, n256, n257, n300, n309, n318, n330, n340, n343, n358,
         n360, n361, n362, n363, n364, n368, n369, n371, n373, n375, n378,
         n384, n388, n391, n395, n410, n411, n429, n430, n431, n432, n436,
         n437, n438, n440, n441, n451, n457, n458, n459, n461, n462, n463,
         n465, n466, n469, n470, n474, n487, n491, n492, n493, n494, n495,
         n496, n497, n498, n501, n502, n503, n504, n512, n513, n517, n518,
         n519, n520, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n534, n535, n538, n539, n540, n541, n542, n543, n544, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n558, n559, n562,
         n563, n564, n566, n567, n569, n570, n571, n572, n575, n576, n577,
         n581, n582, n583, n584, n585, n586, n587, n596, n602, n606, n611,
         n612, n621, n655, n692, n697, n708, n709, n710, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n764, n799, n805, n817,
         n833, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n883, n884, n885, n887, n889,
         n896, n971, n973, n980, n981, n1009, n1053, n1054, n1057, n1062,
         n1063, n1064, n1065, n1082, n1083, n1085, n1086, n1137, n1138, n1139,
         n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
         n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
         n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
         n1172, n1173, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1224, n1225, n1409, n1439, n1459, n1471, n1511, n1561, n1582,
         n1629, n1630, n1751, n1757, n1758, n1759, n1760, n1761, n1762, n1763,
         n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
         n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783,
         n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793,
         n1794, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
         n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1815, n1816, n1817,
         n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1829,
         n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839,
         n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849,
         n1850, n1851, n1852, n1853, n1854, n1855, n1857, n1858, n1859, n1860,
         n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870,
         n1871, n1872, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884,
         n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1895, n1896, n1898,
         n1899, n1902, n1903, n1913, n1916, n1919, n1920, n1921, n1924, n1925,
         n1926, n1929, n1930, n1931, n1932, n1934, n1935, n1936, n1937, n1938,
         n1939, n1940, n1941, n1943, n1944, n1945, n1946, n1947, n1948, n1949,
         n1950, n1951, n1952, n1953, n1954, n1955, n1957, n1958, n1959, n1960,
         n1961, n1962, n1963, n1964, n1965, n1967, n1968, n1969, n1970, n1971,
         n1972, n1973, n1976, n1977, n1978, n1980, n1981, n1982, n1984, n1985,
         n1988, n1989, n1990, n1992, n1994, n1995, n1996, n1997, n1998, n2000,
         n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010,
         n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020,
         n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030,
         n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2039, n2040, n2041,
         n2042, n2044, n2046, n2047, n2048, n2052, n2054, n2055, n2056, n2057,
         n2065, n2066, n2067, n2069, n2071, n2072, n2073, n2074, n2076, n2078,
         n2079, n2080, n2081, n2082, n2084, n2086, n2087, n2088, n2089, n2090,
         n2092, n2094, n2096, n2097, n2098, n2099, n2101, n2102, n2103, n2104,
         n2105, n2106, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115,
         n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125,
         n2126, n2127, n2128, n2129, n2130, n2131, n2133, n2134, n2136, n2137,
         n2138, n2139, n2140, n2142, n2143, n2144, n2145, n2146, n2147, n2148,
         n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158,
         n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168,
         n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178,
         n2180, n2181, n2183, n2184, n2186, n2187, n2189, n2190, n2192, n2193,
         n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203,
         n2204, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214,
         n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224,
         n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234,
         n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245,
         n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255,
         n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2266,
         n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276,
         n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286,
         n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296,
         n2297, n2298, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307,
         n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317,
         n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327,
         n2328, n2329, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338,
         n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348,
         n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358,
         n2359, n2360, n2361, n2362, n2363, n2365, n2366, n2367, n2368, n2369,
         n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379,
         n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389,
         n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399,
         n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409,
         n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419,
         n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429,
         n2430, n2431, n2432, n2434, n2435, n2436, n2437, n2438, n2439, n2440,
         n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450,
         n2451, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461,
         n2462, n2463, n2464, n2465, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493,
         n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503,
         n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513,
         n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523,
         n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2533, n2534,
         n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544,
         n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554,
         n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2565,
         n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575,
         n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585,
         n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2596,
         n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606,
         n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616,
         n2617, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627,
         n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637,
         n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647,
         n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657,
         n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667,
         n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677,
         n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687,
         n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697,
         n2698, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708,
         n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718,
         n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728,
         n2729, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739,
         n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749,
         n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759,
         n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2769, n2770,
         n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780,
         n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790,
         n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800,
         n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810,
         n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2819, n2820, n2821,
         n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831,
         n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841,
         n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2931, n2932, n2933,
         n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943,
         n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953,
         n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963,
         n2964, n2965, n2966, n2968, n2969, n2970, n2971, n2972, n2973, n2974,
         n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984,
         n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994,
         n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004,
         n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014,
         n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024,
         n3025, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035,
         n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045,
         n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055,
         n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n10607,
         n10608, n13840, n13841, n13843, n13844, n13845, n13846, n13847,
         n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856,
         n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864,
         n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13872,
         n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880,
         n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888,
         n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896,
         n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13904,
         n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912,
         n13913, n13914, n13915, n13916, n13917, n13918, n13919, n13920,
         n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928,
         n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936,
         n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13944,
         n13945, n13946, n13947, n13948, n13949, n13950, n13951, n13952,
         n13953, n13954, n13955, n13956, n13957, n13958, n13959, n13960,
         n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968,
         n13969, n13970, n13971, n13972, n13973, n13974, n13975, n13976,
         n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13984,
         n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13992,
         n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000,
         n14001, n14002, n14003, n14004, n14005, n14006, n14007, n14008,
         n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016,
         n14017, n14018, n14019, n14020, n14021, n14022, n14023, n14024,
         n14025, n14026, n14027, n14028, n14029, n14030, n14031, n14032,
         n14033, n14034, n14035, n14036, n14037, n14038, n14039, n14040,
         n14041, n14042, n14043, n14044, n14045, n14046, n14047, n14048,
         n14049, n14050, n14051, n14052, n14053, n14054, n14055, n14056,
         n14057, n14058, n14059, n14060, n14061, n14062, n14063, n14064,
         n14065, n14066, n14067, n14068, n14069, n14070, n14071, n14072,
         n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080,
         n14081, n14082, n14083, n14084, n14085, n14086, n14087, n14088,
         n14089, n14090, n14091, n14092, n14093, n14094, n14095, n14096,
         n14097, n14098, n14099, n14100, n14101, n14102, n14103, n14104,
         n14105, n14106, n14107, n14108, n14109, n14110, n14111, n14112,
         n14113, n14114, n14115, n14116, n14117, n14118, n14119, n14120,
         n14121, n14122, n14123, n14124, n14125, n14126, n14127, n14128,
         n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136,
         n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144,
         n14145, n14146, n14147, n14148, n14149, n14150, n14151, n14152,
         n14153, n14154, n14155, n14156, n14157, n14158, n14159, n14160,
         n14161, n14162, n14163, n14164, n14165, n14167, n14168, n14169,
         n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177,
         n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185,
         n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193,
         n14194, n14195, n14196, n14197, n14202, n14203, n14210, n14211,
         n14218, n14219, n14227, n14228, n14234, n14235, n14243, n14244,
         n14250, n14251, n14258, n14259, n14266, n14267, n14275, n14276,
         n14282, n14283, n14291, n14292, n14298, n14299, n14307, n14308,
         n14314, n14315, n14323, n14324, n14330, n14331, n14339, n14340,
         n14346, n14347, n14355, n14356, n14362, n14363, n14371, n14372,
         n14378, n14379, n14387, n14388, n14394, n14395, n14403, n14404,
         n14410, n14411, n14419, n14420, n14426, n14427, n14436, n14437,
         n14443, n14444, n14449, n14457, n14458, n14459, n14460, n14461,
         n14462, n14463, n14464, n14465, n14466, n14467, n14468, n14469,
         n14470, n14471, n14472, n14473, n14474, n14481, n14482, n14483,
         n14484, n14485, n14486, n14487, n14488, n14495, n14496, n14497,
         n14498, n14499, n14500, n14501, n14502, n14509, n14510, n14511,
         n14512, n14513, n14514, n14515, n14516, n14523, n14524, n14525,
         n14526, n14527, n14528, n14529, n14530, n14537, n14538, n14539,
         n14540, n14541, n14542, n14543, n14544, n14551, n14552, n14553,
         n14554, n14555, n14556, n14557, n14558, n14565, n14566, n14567,
         n14568, n14569, n14570, n14571, n14572, n14579, n14580, n14581,
         n14582, n14583, n14584, n14585, n14586, n14593, n14594, n14595,
         n14596, n14597, n14598, n14599, n14600, n14607, n14608, n14609,
         n14610, n14611, n14612, n14613, n14614, n14621, n14622, n14623,
         n14624, n14625, n14626, n14627, n14628, n14635, n14636, n14637,
         n14638, n14639, n14640, n14641, n14642, n14649, n14650, n14651,
         n14652, n14653, n14654, n14655, n14656, n14663, n14664, n14665,
         n14666, n14667, n14668, n14669, n14670, n14677, n14678, n14679,
         n14680, n14681, n14682, n14683, n14684, n14691, n14692, n14693,
         n14694, n14695, n14696, n14697, n14698, n14705, n14706, n14707,
         n14708, n14709, n14710, n14711, n14712, n14719, n14720, n14721,
         n14722, n14723, n14724, n14725, n14726, n14733, n14734, n14735,
         n14736, n14737, n14738, n14739, n14740, n14747, n14748, n14749,
         n14750, n14751, n14752, n14753, n14754, n14761, n14762, n14763,
         n14764, n14765, n14766, n14767, n14768, n14775, n14776, n14777,
         n14778, n14779, n14780, n14781, n14782, n14789, n14790, n14791,
         n14792, n14793, n14794, n14795, n14796, n14803, n14804, n14805,
         n14806, n14807, n14808, n14809, n14810, n14817, n14818, n14819,
         n14820, n14821, n14822, n14823, n14824, n14831, n14832, n14833,
         n14834, n14835, n14836, n14837, n14838, n14845, n14846, n14847,
         n14848, n14849, n14850, n14851, n14852, n14853, n14854, n14855,
         n14856, n14857, n14864, n14865, n14866, n14867, n14868, n14869,
         n14870, n14871, n14872, n14878, n14879, n14880, n14881, n14882,
         n14890, n14891, n14892, n15219, n15220, n15221, n15318, n15319,
         n15320, n15400, n15401, n15402, n15403, n15404, n15405, n15406,
         n15407, n15408, n15409, n15410, n15411, n15412, n15413, n15414,
         n15415, n15416, n15417, n15418, n15420, n15421, n15422, n15423,
         n15424, n15425, n15426, n15433, n15436, n15437, n15438, n15439,
         n15441, n15442, n15443, n15444, n15445, n15447, n15448, n15449,
         n15450, n15453, n15456, n15458, n15460, n15461, n15462, n15463,
         n15464, n15465, n15466, n15467, n15468, n15469, n15470, n15471,
         n15473, n15474, n15475, n15476, n15481, n15482, n15483, n15484,
         n15487, n15488, n15489, n15490, n15491, n15492, n15493, n15494,
         n15495, n15496, n15497, n15498, n15499, n15500, n15501, n15502,
         n15503, n15504, n15505, n15508, n15509, n15510, n15511, n15512,
         n15513, n15514, n15515, n15516, n15517, n15518, n15519, n15520,
         n15521, n15522, n15523, n15524, n15525, n15526, n15527, n15528,
         n15529, n15530, n15531, n15532, n15533, n15534, n15535, n15539,
         n15544, n15545, n15546, n15547, n15548, n15549, n15550, n15551,
         n15552, n15553, n15554, n15555, n15556, n15557, n15558, n15561,
         n15562, n15563, n15564, n15565, n15566, n15567, n15568, n15569,
         n15571, n15572, n15573, n15574, n15575, n15580, n15581, n15582,
         n15583, n15584, n15585, n15586, n15587, n15588, n15591, n15592,
         n15593, n15594, n15595, n15596, n15597, n15598, n15599, n15600,
         n15601, n15602, n15603, n15604, n15605, n15606, n15607, n15608,
         n15609, n15610, n15613, n15614, n15615, n15616, n15617, n15618,
         n15619, n15620, n15621, n15622, n15623, n15624, n15625, n15626,
         n15627, n15628, n15629, n15630, n15631, n15632, n15633, n15634,
         n15635, n15636, n15637, n15638, n15641, n15646, n15647, n15648,
         n15649, n15650, n15651, n15652, n15653, n15654, n15655, n15656,
         n15657, n15658, n15659, n15660, n15661, n15662, n15663, n15666,
         n15668, n15672, n15673, n15674, n15675, n15676, n15677, n15678,
         n15679, n15680, n15681, n15682, n15683, n15684, n15685, n15686,
         n15687, n15688, n15689, n15690, n15691, n15692, n15695, n15700,
         n15701, n15702, n15703, n15704, n15705, n15706, n15707, n15708,
         n15709, n15710, n15711, n15712, n15713, n15716, n15717, n15718,
         n15719, n15720, n15721, n15722, n15723, n15724, n15725, n15726,
         n15727, n15728, n15729, n15730, n15731, n15732, n15733, n15734,
         n15735, n15736, n15737, n15738, n15739, n15740, n15741, n15742,
         n15743, n15744, n15745, n15746, n15747, n15748, n15749, n15750,
         n15751, n15752, n15753, n15756, n15761, n15762, n15763, n15764,
         n15765, n15766, n15767, n15768, n15769, n15770, n15771, n15772,
         n15773, n15774, n15777, n15779, n15782, n15783, n15784, n15788,
         n15789, n15790, n15791, n15792, n15793, n15794, n15795, n15797,
         n15798, n15799, n15800, n15801, n15802, n15803, n15804, n15805,
         n15807, n15808, n15809, n15810, n15811, n15812, n15813, n15815,
         n15818, n15819, n15820, n15821, n15822, n15823, n15824, n15826,
         n15827, n15828, n15829, n15832, n15834, n15836, n15837, n15838,
         n15839, n15840, n15841, n15842, n15843, n15844, n15845, n15846,
         n15847, n15848, n15849, n15850, n15851, n15852, n15853, n15854,
         n15855, n15856, n15857, n15858, n15860, n15861, n15862, n15863,
         n15864, n15871, n15872, n15873, n15874, n15875, n15876, n15877,
         n15878, n15879, n15880, n15881, n15882, n15883, n15884, n15885,
         n15886, n15887, n15888, n15889, n15890, n15891, n15892, n15893,
         n15896, n15897, n15898, n15899, n15900, n15901, n15904, n15905,
         n15906, n15907, n15909, n15912, n15913, n15914, n15915, n15916,
         n15917, n15918, n15919, n15920, n15921, n15922, n15923, n15924,
         n15925, n15926, n15927, n15928, n15929, n15932, n15938, n15939,
         n15940, n15941, n15942, n15943, n15944, n15945, n15948, n15949,
         n15950, n15953, n15954, n15955, n15956, n15957, n15958, n15961,
         n15962, n15963, n15964, n15965, n15966, n15967, n15968, n15969,
         n15970, n15971, n15972, n15973, n15974, n15975, n15976, n15977,
         n15978, n15979, n15980, n15981, n15982, n15983, n15984, n15985,
         n15986, n15987, n15988, n15990, n15991, n15992, n15993, n16000,
         n16001, n16002, n16003, n16004, n16005, n16006, n16007, n16008,
         n16009, n16010, n16011, n16012, n16013, n16014, n16015, n16016,
         n16017, n16018, n16019, n16020, n16021, n16022, n16023, n16024,
         n16025, n16028, n16029, n16030, n16031, n16032, n16033, n16036,
         n16037, n16038, n16039, n16040, n16041, n16042, n16043, n16044,
         n16045, n16046, n16047, n16048, n16049, n16050, n16051, n16052,
         n16053, n16054, n16055, n16056, n16057, n16058, n16059, n16060,
         n16061, n16062, n16063, n16064, n16065, n16070, n16071, n16074,
         n16075, n16076, n16077, n16078, n16079, n16080, n16081, n16082,
         n16084, n16085, n16086, n16087, n16088, n16089, n16090, n16091,
         n16092, n16093, n16094, n16095, n16096, n16097, n16098, n16099,
         n16100, n16101, n16104, n16105, n16106, n16107, n16108, n16109,
         n16110, n16111, n16113, n16114, n16115, n16116, n16117, n16118,
         n16119, n16120, n16121, n16122, n16123, n16124, n16125, n16126,
         n16127, n16128, n16129, n16130, n16131, n16132, n16137, n16140,
         n16141, n16142, n16143, n16144, n16145, n16146, n16147, n16148,
         n16149, n16150, n16151, n16152, n16153, n16154, n16155, n16156,
         n16158, n16159, n16160, n16161, n16162, n16163, n16164, n16165,
         n16166, n16167, n16168, n16171, n16172, n16173, n16174, n16175,
         n16176, n16177, n16178, n16179, n16180, n16181, n16182, n16183,
         n16184, n16185, n16186, n16187, n16188, n16189, n16190, n16191,
         n16192, n16194, n16195, n16196, n16197, n16198, n16199, n16200,
         n16201, n16202, n16203, n16210, n16211, n16212, n16213, n16214,
         n16215, n16216, n16217, n16218, n16219, n16220, n16221, n16222,
         n16223, n16224, n16225, n16226, n16227, n16228, n16229, n16230,
         n16231, n16232, n16233, n16234, n16235, n16236, n16240, n16241,
         n16242, n16243, n16244, n16245, n16246, n16247, n16248, n16249,
         n16250, n16251, n16252, n16253, n16254, n16255, n16256, n16257,
         n16259, n16260, n16261, n16262, n16263, n16264, n16265, n16266,
         n16267, n16268, n16275, n16276, n16277, n16278, n16279, n16280,
         n16281, n16282, n16283, n16284, n16285, n16286, n16287, n16288,
         n16289, n16290, n16291, n16292, n16293, n16294, n16295, n16296,
         n16297, n16298, n16299, n16300, n16301, n16304, n16305, n16306,
         n16307, n16308, n16309, n16310, n16311, n16312, n16313, n16314,
         n16315, n16316, n16317, n16318, n16319, n16320, n16321, n16322,
         n16323, n16324, n16325, n16326, n16327, n16332, n16335, n16336,
         n16337, n16338, n16339, n16340, n16341, n16342, n16343, n16344,
         n16345, n16346, n16347, n16348, n16349, n16350, n16351, n16352,
         n16353, n16354, n16355, n16356, n16357, n16358, n16359, n16360,
         n16363, n16364, n16365, n16366, n16367, n16368, n16369, n16370,
         n16371, n16372, n16373, n16374, n16375, n16376, n16377, n16378,
         n16379, n16380, n16381, n16382, n16383, n16384, n16385, n16390,
         n16393, n16394, n16395, n16396, n16397, n16398, n16399, n16400,
         n16401, n16402, n16403, n16404, n16405, n16406, n16407, n16408,
         n16409, n16410, n16411, n16412, n16413, n16416, n16417, n16418,
         n16419, n16420, n16421, n16422, n16423, n16424, n16425, n16426,
         n16427, n16428, n16429, n16430, n16431, n16432, n16433, n16434,
         n16435, n16436, n16437, n16438, n16443, n16446, n16447, n16448,
         n16449, n16450, n16451, n16452, n16453, n16454, n16455, n16456,
         n16457, n16458, n16459, n16460, n16461, n16462, n16463, n16464,
         n16465, n16466, n16467, n16468, n16471, n16472, n16473, n16474,
         n16475, n16476, n16477, n16478, n16479, n16480, n16481, n16482,
         n16483, n16484, n16485, n16486, n16487, n16488, n16489, n16490,
         n16491, n16492, n16493, n16498, n16501, n16502, n16503, n16504,
         n16505, n16506, n16507, n16508, n16509, n16510, n16511, n16512,
         n16513, n16514, n16515, n16516, n16517, n16518, n16519, n16520,
         n16521, n16522, n16525, n16526, n16527, n16528, n16529, n16530,
         n16532, n16533, n16534, n16535, n16536, n16537, n16538, n16539,
         n16540, n16541, n16542, n16544, n16545, n16546, n16547, n16554,
         n16555, n16556, n16557, n16558, n16559, n16560, n16561, n16562,
         n16563, n16566, n16567, n16568, n16569, n16570, n16571, n16572,
         n16573, n16574, n16575, n16576, n16577, n16578, n16579, n16582,
         n16583, n16584, n16585, n16586, n16587, n16588, n16589, n16590,
         n16591, n16592, n16593, n16594, n16595, n16596, n16597, n16598,
         n16599, n16600, n16601, n16602, n16603, n16604, n16605, n16606,
         n16607, n16608, n16616, n16617, n16618, n16619, n16621, n16622,
         n16623, n16624, n16625, n16626, n16627, n16628, n16629, n16630,
         n16631, n16632, n16633, n16634, n16635, n16636, n16637, n16640,
         n16641, n16642, n16645, n16646, n16647, n16648, n16649, n16650,
         n16651, n16652, n16653, n16656, n16657, n16658, n16659, n16660,
         n16661, n16662, n16663, n16665, n16666, n16667, n16668, n16669,
         n16671, n16672, n16673, n16674, n16675, n16682, n16683, n16684,
         n16685, n16686, n16687, n16688, n16689, n16690, n16691, n16692,
         n16693, n16694, n16695, n16696, n16697, n16698, n16701, n16702,
         n16703, n16704, n16705, n16706, n16707, n16708, n16709, n16710,
         n16711, n16712, n16713, n16714, n16715, n16716, n16717, n16718,
         n16719, n16721, n16722, n16723, n16724, n16725, n16726, n16727,
         n16728, n16729, n16736, n16737, n16738, n16739, n16740, n16741,
         n16742, n16743, n16744, n16745, n16746, n16747, n16748, n16749,
         n16750, n16751, n16752, n16755, n16756, n16757, n16758, n16759,
         n16760, n16761, n16762, n16763, n16764, n16765, n16766, n16767,
         n16768, n16769, n16771, n16772, n16773, n16774, n16775, n16776,
         n16778, n16779, n16780, n16781, n16782, n16789, n16790, n16791,
         n16792, n16793, n16794, n16795, n16796, n16797, n16798, n16799,
         n16800, n16801, n16802, n16803, n16804, n16805, n16808, n16809,
         n16810, n16811, n16812, n16813, n16814, n16815, n16817, n16818,
         n16819, n16820, n16821, n16822, n16823, n16824, n16825, n16826,
         n16828, n16829, n16830, n16831, n16832, n16833, n16834, n16841,
         n16842, n16843, n16844, n16845, n16846, n16847, n16848, n16849,
         n16850, n16851, n16852, n16853, n16854, n16855, n16856, n16857,
         n16860, n16861, n16862, n16863, n16864, n16865, n16866, n16867,
         n16868, n16869, n16870, n16871, n16872, n16873, n16874, n16875,
         n16876, n16878, n16879, n16880, n16881, n16888, n16889, n16890,
         n16891, n16892, n16893, n16894, n16895, n16896, n16897, n16898,
         n16899, n16900, n16901, n16902, n16903, n16904, n16905, n16906,
         n16907, n16908, n16909, n16910, n16911, n16912, n16915, n16916,
         n16917, n16918, n16919, n16920, n16921, n16922, n16923, n16924,
         n16925, n16926, n16927, n16929, n16930, n16931, n16932, n16933,
         n16934, n16936, n16937, n16938, n16939, n16940, n16941, n16942,
         n16949, n16950, n16951, n16952, n16953, n16954, n16955, n16956,
         n16957, n16958, n16959, n16960, n16961, n16962, n16963, n16966,
         n16967, n16968, n16969, n16970, n16971, n16972, n16973, n16974,
         n16975, n16976, n16977, n16978, n16979, n16980, n16981, n16982,
         n16983, n16984, n16985, n16986, n16987, n16988, n16989, n16990,
         n16991, n16992, n16993, n16994, n16995, n16996, n16997, n16998,
         n16999, n17000, n17001, n17002, n17004, n17005, n17006, n17007,
         n17014, n17015, n17016, n17017, n17018, n17019, n17020, n17021,
         n17022, n17023, n17024, n17025, n17027, n17028, n17029, n17030,
         n17031, n17032, n17033, n17034, n17035, n17036, n17037, n17038,
         n17039, n17040, n17041, n17042, n17043, n17044, n17050, n17052,
         n17054, n17055, n17056, n17057, n17058, n17060, n17061, n17062,
         n17063, n17064, n17065, n17066, n17067, n17068, n17070, n17071,
         n17072, n17073, n17080, n17081, n17082, n17083, n17084, n17085,
         n17086, n17087, n17088, n17089, n17090, n17091, n17092, n17093,
         n17094, n17095, n17096, n17097, n17099, n17101, n17103, n17104,
         n17105, n17106, n17107, n17108, n17109, n17112, n17113, n17114,
         n17115, n17116, n17117, n17118, n17119, n17120, n17121, n17122,
         n17123, n17124, n17125, n17126, n17127, n17128, n17129, n17130,
         n17131, n17132, n17133, n17134, n17135, n17136, n17137, n17138,
         n17139, n17140, n17143, n17144, n17145, n17146, n17153, n17154,
         n17155, n17156, n17157, n17158, n17159, n17160, n17164, n17165,
         n17166, n17167, n17168, n17169, n17170, n17171, n17172, n17173,
         n17174, n17175, n17176, n17177, n17178, n17179, n17180, n17181,
         n17182, n17183, n17186, n17187, n17188, n17189, n17190, n17191,
         n17192, n17193, n17196, n17197, n17198, n17199, n17200, n17201,
         n17203, n17204, n17205, n17206, n17207, n17316, n17317, n17318,
         n17319, n17320, n17321, n17322, n17324, n17325, n17326, n17327,
         n17328, n17331, n17332, n17333, n17334, n17340, n17341, n17342,
         n17343, n17344, n17345, n17348, n17349, n17350, n17351, n17352,
         n17353, n17354, n17355, n17356, n17357, n17358, n17359, n17360,
         n17361, n17362, n17363, n17364, n17365, n17366, n17367, n17368,
         n17369, n17370, n17371, n17372, n17373, n17375, n17376, n17378,
         n17379, n17380, n17381, n17382, n17383, n17384, n17385, n17386,
         n17387, n17388, n17389, n17390, n17391, n17392, n17393, n17394,
         n17395, n17396, n17397, n17398, n17399, n17400, n17401, n17402,
         n17403, n17404, n17405, n17406, n17407, n17413, n17414, n17415,
         n17416, n17417, n17425, n17426, n17427, n17444, n17446, n17447,
         n17448, n17449, n17450, n17451, n17452, n17453, n17454, n17455,
         n17456, n17457, n17458, n17459, n17460, n17461, n17462, n17463,
         n17464, n17465, n17466, n17467, n17468, n17469, n17470, n17471,
         n17472, n17473, n17474, n17475, n17476, n17477, n17478, n17479,
         n17480, n17481, n17482, n17483, n17484, n17485, n17486, n17487,
         n17488, n17489, n17490, n17491, n17492, n17493, n17494, n17495,
         n17496, n17497, n17498, n17499, n17500, n17501, n17502, n17503,
         n17504, n17505, n17506, n17507, n17508, n17509, n17510, n17511,
         n17512, n17513, n17514, n17515, n17516, n17517, n17518, n17519,
         n17520, n17521, n17522, n17523, n17524, n17525, n17526, n17527,
         n17528, n17529, n17530, n17531, n17532, n17533, n17534, n17539,
         n17540, n17541, n17542, n17543, n17544, n17545, n17546, n17547,
         n17548, n17549, n17550, n17551, n17552, n17553, n17554, n17560,
         n17561, n17562, n17563, n17564, n17565, n17566, n17567, n17568,
         n17569, n17570, n17571, n17572, n17573, n17577, n17578, n17584,
         n17585, n17768, n17769, n17770, n17771, n17781, n17782, n17796,
         n17808, n17809, n17810, n17811, n17812, n17813, n17814, n17815,
         n17824, n17833, n17834, n17835, n17836, n17845, n17854, n17855,
         n17856, n17857, n17858, n17859, n17868, n17869, n17880, n17883,
         n17896, n17898, n17899, n17900, n17909, n17910, n17937, n17938,
         n17943, n17944, n17949, n18000, n18002, n18003, n18009, n18011,
         n18016, n18018, n18023, n18025, n18030, n18032, n18037, n18039,
         n18044, n18046, n18051, n18053, n18058, n18060, n18065, n18067,
         n18072, n18074, n18079, n18081, n18086, n18089, n18095, n18097,
         n18102, n18104, n18109, n18111, n18116, n18118, n18123, n18125,
         n18130, n18132, n18137, n18139, n18144, n18146, n18151, n18153,
         n18158, n18160, n18165, n18167, n18172, n18174, n18179, n18181,
         n18186, n18188, n18193, n18195, n18200, n18202, n18207, n18209,
         n18214, n18216, n18221, n18223, n18228, n18229, n18234, n18235,
         n18240, n18241, n18246, n18247, n18252, n18253, n18258, n18259,
         n18264, n18265, n18270, n18271, n18276, n18277, n18282, n18283,
         n18288, n18289, n18294, n18295, n18296, n18297, n18299, n18303,
         n18305, n18306, n18313, n18314, n18319, n18320, n18325, n18326,
         n18331, n18332, n18337, n18338, n18343, n18344, n18349, n18350,
         n18355, n18356, n18361, n18362, n18367, n18368, n18373, n18374,
         n18379, n18380, n18385, n18386, n18391, n18392, n18397, n18398,
         n18403, n18404, n18409, n18410, n18415, n18416, n18421, n18422,
         n18427, n18428, n18433, n18434, n18439, n18440, n18445, n18446,
         n18451, n18452, n18457, n18458, n18463, n18464, n18469, n18470,
         n18475, n18476, n18481, n18482, n18487, n18488, n18493, n18494,
         n18499, n18501, n18507, n18508, n18513, n18514, n18519, n18520,
         n18525, n18526, n18531, n18532, n18537, n18538, n18543, n18544,
         n18549, n18550, n18555, n18556, n18561, n18562, n18567, n18568,
         n18573, n18574, n18579, n18580, n18585, n18586, n18591, n18592,
         n18597, n18598, n18603, n18604, n18609, n18610, n18615, n18616,
         n18621, n18622, n18627, n18628, n18633, n18634, n18639, n18640,
         n18645, n18646, n18651, n18652, n18657, n18658, n18663, n18664,
         n18669, n18670, n18675, n18676, n18681, n18682, n18687, n18688,
         n18689, n18691, n18695, n18696, n18697, n18703, n18704, n18709,
         n18710, n18715, n18716, n18721, n18722, n18727, n18728, n18733,
         n18734, n18739, n18740, n18745, n18746, n18751, n18752, n18757,
         n18758, n18763, n18764, n18769, n18770, n18775, n18776, n18781,
         n18782, n18787, n18788, n18793, n18794, n18799, n18800, n18805,
         n18806, n18811, n18812, n18817, n18818, n18823, n18824, n18829,
         n18830, n18835, n18836, n18841, n18842, n18847, n18848, n18853,
         n18854, n18859, n18860, n18865, n18866, n18871, n18872, n18877,
         n18878, n18883, n18884, n18885, n18887, n18891, n18893, n18899,
         n18900, n18905, n18906, n18911, n18912, n18917, n18918, n18923,
         n18924, n18929, n18930, n18935, n18936, n18941, n18942, n18947,
         n18948, n18953, n18954, n18959, n18960, n18965, n18966, n18971,
         n18972, n18977, n18978, n18983, n18984, n18989, n18990, n18995,
         n18996, n19001, n19002, n19007, n19008, n19013, n19014, n19019,
         n19020, n19025, n19026, n19031, n19032, n19037, n19038, n19043,
         n19044, n19049, n19050, n19055, n19056, n19061, n19062, n19067,
         n19068, n19073, n19074, n19079, n19080, n19081, n19083, n19087,
         n19088, n19089, n19095, n19096, n19101, n19102, n19107, n19108,
         n19113, n19114, n19119, n19120, n19125, n19126, n19131, n19132,
         n19137, n19138, n19143, n19144, n19149, n19150, n19155, n19156,
         n19161, n19162, n19167, n19168, n19173, n19174, n19179, n19180,
         n19185, n19186, n19191, n19192, n19197, n19198, n19203, n19204,
         n19209, n19210, n19215, n19216, n19221, n19222, n19227, n19228,
         n19233, n19234, n19239, n19240, n19245, n19246, n19251, n19252,
         n19257, n19258, n19263, n19264, n19269, n19270, n19275, n19276,
         n19277, n19279, n19283, n19285, n19291, n19292, n19297, n19298,
         n19303, n19304, n19309, n19310, n19315, n19316, n19321, n19322,
         n19327, n19328, n19333, n19334, n19339, n19340, n19345, n19346,
         n19351, n19352, n19357, n19358, n19363, n19364, n19369, n19370,
         n19375, n19376, n19381, n19382, n19387, n19388, n19393, n19394,
         n19399, n19400, n19405, n19406, n19411, n19412, n19417, n19418,
         n19423, n19424, n19429, n19430, n19435, n19436, n19441, n19442,
         n19447, n19448, n19453, n19454, n19459, n19460, n19465, n19466,
         n19471, n19472, n19473, n19475, n19479, n19481, n19482, n19489,
         n19490, n19495, n19496, n19501, n19502, n19507, n19508, n19513,
         n19514, n19519, n19520, n19525, n19526, n19531, n19532, n19537,
         n19538, n19543, n19544, n19549, n19550, n19555, n19556, n19561,
         n19562, n19567, n19568, n19573, n19574, n19579, n19580, n19585,
         n19586, n19591, n19592, n19597, n19598, n19603, n19604, n19609,
         n19610, n19615, n19616, n19621, n19622, n19627, n19628, n19633,
         n19634, n19639, n19640, n19645, n19646, n19651, n19652, n19657,
         n19658, n19663, n19664, n19669, n19670, n19671, n19676, n19678,
         n19679, n19686, n19687, n19692, n19693, n19698, n19699, n19704,
         n19705, n19710, n19711, n19716, n19717, n19722, n19723, n19728,
         n19729, n19734, n19735, n19740, n19741, n19746, n19747, n19752,
         n19753, n19758, n19759, n19764, n19765, n19770, n19771, n19776,
         n19777, n19782, n19783, n19788, n19789, n19794, n19795, n19800,
         n19801, n19806, n19807, n19812, n19813, n19818, n19819, n19824,
         n19825, n19830, n19831, n19836, n19837, n19842, n19843, n19848,
         n19849, n19854, n19855, n19860, n19861, n19866, n19867, n19868,
         n19873, n19875, n19876, n19883, n19884, n19889, n19890, n19895,
         n19896, n19901, n19902, n19907, n19908, n19913, n19914, n19919,
         n19920, n19925, n19926, n19931, n19932, n19937, n19938, n19943,
         n19944, n19949, n19950, n19955, n19956, n19961, n19962, n19967,
         n19968, n19973, n19974, n19979, n19980, n19985, n19986, n19991,
         n19992, n19997, n19998, n20003, n20004, n20009, n20010, n20015,
         n20016, n20021, n20022, n20027, n20028, n20033, n20034, n20039,
         n20040, n20045, n20046, n20051, n20052, n20057, n20058, n20063,
         n20064, n20069, n20071, n20072, n20079, n20080, n20085, n20086,
         n20091, n20092, n20097, n20098, n20103, n20104, n20109, n20110,
         n20115, n20116, n20121, n20122, n20127, n20128, n20133, n20134,
         n20139, n20140, n20145, n20146, n20151, n20152, n20157, n20158,
         n20163, n20164, n20169, n20170, n20175, n20176, n20181, n20182,
         n20187, n20188, n20193, n20194, n20199, n20200, n20205, n20206,
         n20211, n20212, n20217, n20218, n20223, n20224, n20229, n20230,
         n20235, n20236, n20241, n20242, n20247, n20248, n20253, n20254,
         n20259, n20260, n20265, n20267, n20268, n20275, n20276, n20281,
         n20282, n20287, n20288, n20293, n20294, n20299, n20300, n20305,
         n20306, n20311, n20312, n20317, n20318, n20323, n20324, n20329,
         n20330, n20335, n20336, n20341, n20342, n20347, n20348, n20353,
         n20354, n20359, n20360, n20365, n20366, n20371, n20372, n20377,
         n20378, n20383, n20384, n20389, n20390, n20395, n20396, n20401,
         n20402, n20407, n20408, n20413, n20414, n20419, n20420, n20425,
         n20426, n20431, n20432, n20437, n20438, n20443, n20444, n20449,
         n20450, n20455, n20456, n20461, n20464, n20471, n20472, n20477,
         n20478, n20483, n20484, n20489, n20490, n20495, n20496, n20501,
         n20502, n20507, n20508, n20513, n20514, n20519, n20520, n20525,
         n20526, n20531, n20532, n20537, n20538, n20543, n20544, n20549,
         n20550, n20555, n20556, n20561, n20562, n20567, n20568, n20573,
         n20574, n20579, n20580, n20585, n20586, n20591, n20592, n20597,
         n20598, n20603, n20604, n20609, n20610, n20615, n20616, n20621,
         n20622, n20627, n20628, n20633, n20634, n20639, n20640, n20645,
         n20646, n20651, n20652, n20657, n20659, n20660, n20667, n20668,
         n20673, n20674, n20679, n20680, n20685, n20686, n20691, n20692,
         n20697, n20698, n20703, n20704, n20709, n20710, n20715, n20716,
         n20721, n20722, n20727, n20728, n20733, n20734, n20739, n20740,
         n20745, n20746, n20751, n20752, n20757, n20758, n20763, n20764,
         n20769, n20770, n20775, n20776, n20781, n20782, n20787, n20788,
         n20793, n20794, n20799, n20800, n20805, n20806, n20811, n20812,
         n20817, n20818, n20823, n20824, n20829, n20830, n20835, n20836,
         n20841, n20842, n20847, n20848, n20853, n20856, n20863, n20864,
         n20869, n20870, n20875, n20876, n20881, n20882, n20887, n20888,
         n20893, n20894, n20899, n20900, n20905, n20906, n20911, n20912,
         n20917, n20918, n20923, n20924, n20929, n20930, n20935, n20936,
         n20941, n20942, n20947, n20948, n20953, n20954, n20959, n20960,
         n20965, n20966, n20971, n20972, n20977, n20978, n20983, n20984,
         n20989, n20990, n20995, n20996, n21001, n21002, n21007, n21008,
         n21013, n21014, n21019, n21020, n21025, n21026, n21031, n21032,
         n21037, n21038, n21043, n21044, n21049, n21051, n21052, n21059,
         n21060, n21065, n21066, n21071, n21072, n21077, n21078, n21083,
         n21084, n21089, n21090, n21095, n21096, n21101, n21102, n21107,
         n21108, n21113, n21114, n21119, n21120, n21125, n21126, n21131,
         n21132, n21137, n21138, n21143, n21144, n21149, n21150, n21155,
         n21156, n21161, n21162, n21167, n21168, n21173, n21174, n21179,
         n21180, n21185, n21186, n21191, n21192, n21197, n21198, n21203,
         n21204, n21209, n21210, n21215, n21216, n21221, n21222, n21227,
         n21228, n21233, n21234, n21239, n21240, n21241, n21246, n21249,
         n21256, n21257, n21262, n21263, n21268, n21269, n21274, n21275,
         n21280, n21281, n21286, n21287, n21292, n21293, n21298, n21299,
         n21304, n21305, n21310, n21311, n21316, n21317, n21322, n21323,
         n21328, n21329, n21334, n21335, n21340, n21341, n21346, n21347,
         n21352, n21353, n21358, n21359, n21364, n21365, n21370, n21371,
         n21376, n21377, n21382, n21383, n21388, n21389, n21394, n21395,
         n21400, n21401, n21406, n21407, n21412, n21413, n21418, n21419,
         n21424, n21425, n21430, n21431, n21436, n21437, n21438, n21443,
         n21445, n21446, n21453, n21454, n21459, n21460, n21465, n21466,
         n21471, n21472, n21477, n21478, n21483, n21484, n21489, n21490,
         n21495, n21496, n21501, n21502, n21507, n21508, n21513, n21514,
         n21519, n21520, n21525, n21526, n21531, n21532, n21537, n21538,
         n21543, n21544, n21549, n21550, n21555, n21556, n21561, n21562,
         n21567, n21568, n21573, n21574, n21579, n21580, n21585, n21586,
         n21591, n21592, n21597, n21598, n21603, n21604, n21609, n21610,
         n21615, n21616, n21621, n21622, n21627, n21628, n21633, n21634,
         n21639, n21641, n21642, n21649, n21650, n21655, n21656, n21661,
         n21662, n21667, n21668, n21673, n21674, n21679, n21680, n21685,
         n21686, n21691, n21692, n21697, n21698, n21703, n21704, n21709,
         n21710, n21715, n21716, n21721, n21722, n21727, n21728, n21733,
         n21734, n21739, n21740, n21745, n21746, n21751, n21752, n21757,
         n21758, n21763, n21764, n21769, n21770, n21775, n21776, n21781,
         n21782, n21787, n21788, n21793, n21794, n21799, n21800, n21805,
         n21806, n21811, n21812, n21817, n21818, n21823, n21824, n21829,
         n21830, n21835, n21837, n21838, n21845, n21846, n21851, n21852,
         n21857, n21858, n21863, n21864, n21869, n21870, n21875, n21876,
         n21881, n21882, n21887, n21888, n21893, n21894, n21899, n21900,
         n21905, n21906, n21911, n21912, n21917, n21918, n21923, n21924,
         n21929, n21930, n21935, n21936, n21941, n21942, n21947, n21948,
         n21953, n21954, n21959, n21960, n21965, n21966, n21971, n21972,
         n21977, n21978, n21983, n21984, n21989, n21990, n21995, n21996,
         n22001, n22002, n22007, n22008, n22013, n22014, n22019, n22020,
         n22025, n22026, n22031, n22033, n22034, n22041, n22042, n22047,
         n22048, n22053, n22054, n22059, n22060, n22065, n22066, n22071,
         n22072, n22077, n22078, n22083, n22084, n22089, n22090, n22095,
         n22096, n22101, n22102, n22107, n22108, n22113, n22114, n22119,
         n22120, n22125, n22126, n22131, n22132, n22137, n22138, n22143,
         n22144, n22149, n22150, n22155, n22156, n22161, n22162, n22167,
         n22168, n22173, n22174, n22179, n22180, n22185, n22186, n22191,
         n22192, n22197, n22198, n22203, n22204, n22209, n22210, n22215,
         n22216, n22221, n22222, n22227, n22229, n22230, n22237, n22238,
         n22243, n22244, n22249, n22250, n22255, n22256, n22261, n22262,
         n22267, n22268, n22273, n22274, n22279, n22280, n22285, n22286,
         n22291, n22292, n22297, n22298, n22303, n22304, n22309, n22310,
         n22315, n22316, n22321, n22322, n22327, n22328, n22333, n22334,
         n22339, n22340, n22345, n22346, n22351, n22352, n22357, n22358,
         n22363, n22364, n22369, n22370, n22375, n22376, n22381, n22382,
         n22387, n22388, n22393, n22394, n22399, n22400, n22405, n22406,
         n22411, n22412, n22417, n22418, n22423, n22425, n22426, n22433,
         n22434, n22439, n22440, n22445, n22446, n22451, n22452, n22457,
         n22458, n22463, n22464, n22469, n22470, n22475, n22476, n22481,
         n22482, n22487, n22488, n22493, n22494, n22499, n22500, n22505,
         n22506, n22511, n22512, n22517, n22518, n22523, n22524, n22529,
         n22530, n22535, n22536, n22541, n22542, n22547, n22548, n22553,
         n22554, n22559, n22560, n22565, n22566, n22571, n22572, n22577,
         n22578, n22583, n22584, n22589, n22590, n22595, n22596, n22601,
         n22602, n22607, n22608, n22613, n22614, n22619, n22622, n22629,
         n22630, n22635, n22636, n22641, n22642, n22647, n22648, n22653,
         n22654, n22659, n22660, n22665, n22667, n22668, n22675, n22676,
         n22681, n22682, n22687, n22688, n22693, n22694, n22699, n22700,
         n22705, n22706, n22711, n22712, n22717, n22718, n22723, n22724,
         n22729, n22730, n22735, n22736, n22741, n22742, n22747, n22748,
         n22753, n22754, n22759, n22760, n22765, n22766, n22771, n22772,
         n22777, n22778, n22783, n22784, n22789, n22790, n22795, n22796,
         n22801, n22802, n22807, n22808, n22813, n22814, n22819, n22820,
         n22825, n22826, n22831, n22832, n22837, n22838, n22843, n22844,
         n22849, n22850, n22855, n22856, n22861, n22862, n22867, n22868,
         n22873, n22874, n22879, n22880, n22885, n22887, n22888, n22895,
         n22896, n22901, n22902, n22907, n22908, n22913, n22914, n22919,
         n22920, n22925, n22926, n22931, n22932, n22937, n22938, n22943,
         n22944, n22949, n22950, n22955, n22956, n22961, n22962, n22967,
         n22968, n22973, n22974, n22979, n22980, n22985, n22986, n22991,
         n22992, n22997, n22998, n23003, n23004, n23009, n23010, n23015,
         n23016, n23021, n23022, n23027, n23028, n23033, n23034, n23039,
         n23040, n23045, n23046, n23051, n23052, n23057, n23058, n23063,
         n23064, n23069, n23070, n23075, n23076, n23081, n23082, n23087,
         n23088, n23093, n23094, n23099, n23100, n23105, n23107, n23108,
         n23115, n23116, n23121, n23122, n23127, n23128, n23133, n23134,
         n23139, n23140, n23145, n23146, n23151, n23152, n23157, n23158,
         n23163, n23164, n23169, n23170, n23175, n23176, n23181, n23182,
         n23187, n23188, n23193, n23194, n23199, n23200, n23205, n23206,
         n23211, n23212, n23217, n23218, n23223, n23224, n23229, n23230,
         n23235, n23236, n23241, n23242, n23247, n23248, n23253, n23254,
         n23259, n23260, n23265, n23266, n23271, n23272, n23277, n23278,
         n23283, n23284, n23289, n23290, n23295, n23296, n23301, n23302,
         n23307, n23308, n23313, n23314, n23319, n23321, n23322, n23329,
         n23330, n23335, n23336, n23341, n23342, n23347, n23348, n23353,
         n23354, n23359, n23360, n23365, n23366, n23371, n23372, n23377,
         n23378, n23383, n23384, n23389, n23390, n23395, n23396, n23401,
         n23402, n23407, n23408, n23413, n23414, n23419, n23420, n23425,
         n23426, n23431, n23432, n23437, n23438, n23443, n23444, n23449,
         n23450, n23455, n23456, n23461, n23462, n23467, n23468, n23473,
         n23474, n23479, n23480, n23485, n23486, n23491, n23492, n23497,
         n23498, n23503, n23504, n23509, n23510, n23515, n23516, n23521,
         n23522, n23527, n23528, n23533, n23534, n23539, n23541, n23542,
         n23549, n23550, n23555, n23556, n23561, n23562, n23567, n23568,
         n23573, n23574, n23579, n23580, n23585, n23586, n23591, n23592,
         n23597, n23598, n23603, n23604, n23609, n23610, n23615, n23616,
         n23621, n23622, n23627, n23628, n23633, n23634, n23639, n23640,
         n23645, n23646, n23651, n23652, n23657, n23658, n23663, n23664,
         n23669, n23670, n23675, n23676, n23681, n23682, n23687, n23688,
         n23693, n23694, n23699, n23700, n23705, n23706, n23711, n23712,
         n23717, n23718, n23723, n23724, n23729, n23730, n23735, n23736,
         n23741, n23742, n23747, n23748, n23753, n23754, n23759, n23761,
         n23762, n23769, n23770, n23775, n23776, n23781, n23782, n23787,
         n23788, n23793, n23794, n23799, n23800, n23805, n23806, n23811,
         n23812, n23817, n23818, n23823, n23824, n23829, n23830, n23835,
         n23836, n23841, n23842, n23847, n23848, n23853, n23854, n23859,
         n23860, n23865, n23866, n23871, n23872, n23877, n23878, n23883,
         n23884, n23889, n23890, n23895, n23896, n23901, n23902, n23907,
         n23908, n23913, n23914, n23919, n23920, n23925, n23926, n23931,
         n23932, n23937, n23938, n23943, n23944, n23949, n23950, n23955,
         n23956, n23961, n23962, n23967, n23968, n23973, n23974, n23979,
         n23980, n23985, n23986, n23991, n23992, n23997, n23998, n24003,
         n24004, n24009, n24010, n24015, n24016, n24021, n24022, n24027,
         n24028, n24033, n24034, n24039, n24040, n24045, n24046, n24051,
         n24052, n24057, n24058, n24063, n24064, n24069, n24070, n24075,
         n24076, n24081, n24082, n24087, n24088, n24093, n24094, n24099,
         n24100, n24101, n24102, n24104, n24108, n24109, n24110, n24112,
         n24113, n24114, n24115, n24117, n24119, n24120, n24121, n24122,
         n24123, n24125, n24129, n24134, n24135, n24136, n24140, n24144,
         n24145, n24149, n24153, n24154, n24158, n24161, n24162, n24164,
         n24165, n24166, n24167, n24170, n24175, n24179, n24180, n24184,
         n24188, n24190, n24191, n24192, n24193, n24196, n24200, n24203,
         n24207, n24210, n24212, n24213, n24214, n24217, n24219, n24220,
         n24221, n24224, n24225, n24226, n24227, n24228, n24229, n24231,
         n24232, n24233, n24234, n24235, n24237, n24239, n24243, n24247,
         n24252, n24256, n24260, n24263, n24267, n24270, n24271, n24272,
         n24273, n24274, n24275, n24278, n24279, n24280, n24283, n24285,
         n24286, n24287, n24290, n24291, n24292, n24293, n24294, n24295,
         n24296, n24298, n24299, n24300, n24301, n24302, n24306, n24312,
         n24316, n24319, n24323, n24328, n24333, n24336, n24337, n24341,
         n24347, n24348, n24349, n24350, n24353, n24355, n24356, n24357,
         n24361, n24365, n24366, n24367, n24376, n24378, n24379, n24381,
         n24382, n24383, n24384, n24385, n24386, n24387, n24388, n24389,
         n24397, n24403, n24405, n24406, n24407, n24409, n24410, n24411,
         n24412, n24413, n24414, n24415, n24416, n24419, n24420, n24421,
         n24422, n24425, n24426, n24429, n24430, n24431, n24432, n24433,
         n24434, n24435, n24436, n24437, n24438, n24440, n24441, n24442,
         n24443, n24444, n24445, n24446, n24447, n24448, n24449, n24450,
         n24451, n24452, n24453, n24454, n24455, n24456, n24457, n24458,
         n24459, n24460, n24461, n24462, n24463, n24464, n24469, n24473,
         n24474, n24488, n24502, n24504, n24508, n24511, n24512, n24513,
         n24514, n24515, n24516, n24517, n24518, n24519, n24520, n24522,
         n24523, n24524, n24525, n24526, n24527, n24528, n24529, n24530,
         n24533, n24535, n24538, n24539, n24552, n24555, n24556, n24557,
         n24564, n24565, n24566, n24570, n24571, n24572, n24573, n24574,
         n24839, n24842, n24845, n24847, n24848, n24849, n24850, n24851,
         n24852, n24853, n24854, n24855, n24856, n24861, n24862, n24863,
         n24864, n24865, n24866, n24867, n24868, n24871, n24872, n24873,
         n24874, n24876, n24877, n24878, n24879, n24880, n24881, n24884,
         n24885, n24886, n24887, n24889, n24890, n24892, n24893, n24894,
         n24895, n24898, n24899, n24900, n24901, n24902, n24903, n24904,
         n24905, n24906, n24907, n24908, n24909, n24910, n24911, n24912,
         n24913, n24914, n24915, n24916, n24917, n24918, n24919, n24920,
         n24921, n24922, n24923, n24924, n24925, n24926, n24927, n24928,
         n24929, n24930, n24931, n24932, n24933, n24934, n24935, n24936,
         n24937, n24938, n24940, n24941, n24942, n24943, n24944, n24945,
         n24946, n24947, n24948, n24949, n24950, n24951, n24952, n24953,
         n24954, n24955, n24956, n24957, n24958, n24959, n24960, n24961,
         n24962, n24963, n24964, n24965, n24966, n24967, n24968, n24969,
         n24970, n24971, n24972, n24973, n24974, n24975, n24976, n24977,
         n24978, n24979, n24980, n24981, n24982, n24983, n24984, n24985,
         n24986, n24987, n24988, n24989, n24990, n24991, n24992, n24993,
         n24994, n24995, n24996, n24997, n24998, n24999, n25000, n25001,
         n25002, n25003, n25004, n25005, n25006, n25007, n25008, n25009,
         n25010, n25011, n25012, n25013, n25014, n25015, n25016, n25017,
         n25018, n25019, n25020, n25021, n25022, n25023, n25024, n25025,
         n25026, n25027, n25028, n25029, n25030, n25031, n25032, n25033,
         n25034, n25035, n25036, n25037, n25038, n25039, n25040, n25041,
         n25042, n25043, n25044, n25045, n25046, n25047, n25048, n25049,
         n25050, n25051, n25052, n25053, n25054, n25055, n25057, n25058,
         n25059, n25060, n25061, n25062, n25063, n25064, n25065, n25066,
         n25067, n25068, n25069, n25070, n25071, n25072, n25073, n25074,
         n25075, n25076, n25077, n25078, n25079, n25080, n25081, n25082,
         n25083, n25084, n25085, n25086, n25087, n25088, n25089, n25090,
         n25091, n25092, n25093, n25094, n25095, n25096, n25097, n25098,
         n25099, n25100, n25101, n25102, n25103, n25104, n25105, n25106,
         n25107, n25108, n25109, n25110, n25111, n25112, n25113, n25114,
         n25115, n25116, n25117, n25118, n25119, n25120, n25121, n25122,
         n25123, n25124, n25125, n25126, n25127, n25128, n25129, n25130,
         n25131, n25132, n25133, n25134, n25135, n25136, n25137, n25138,
         n25139, n25140, n25141, n25142, n25143, n25144, n25145, n25146,
         n25147, n25148, n25149, n25150, n25151, n25152, n25153, n25154,
         n25155, n25156, n25157, n25158, n25159, n25160, n25161, n25162,
         n25163, n25164, n25165, n25166, n25167, n25168, n25169, n25170,
         n25171, n25172, n25173, n25174, n25175, n25176, n25177, n25178,
         n25179, n25180, n25181, n25182, n25183, n25184, n25185, n25186,
         n25187, n25188, n25189, n25190, n25191, n25192, n25193, n25194,
         n25195, n25196, n25197, n25198, n25199, n25200, n25201, n25202,
         n25203, n25204, n25205, n25206, n25207, n25208, n25209, n25210,
         n25211, n25212, n25213, n25214, n25215, n25216, n25217, n25218,
         n25219, n25220, n25221, n25222, n25223, n25224, n25225, n25226,
         n25227, n25228, n25229, n25230, n25231, n25232, n25233, n25234,
         n25235, n25236, n25237, n25238, n25239, n25240, n25241, n25242,
         n25243, n25244, n25245, n25246, n25247, n25248, n25249, n25250,
         n25251, n25252, n25253, n25254, n25255, n25256, n25257, n25258,
         n25259, n25260, n25261, n25262, n25263, n25264, n25265, n25266,
         n25267, n25268, n25269, n25270, n25271, n25272, n25273, n25274,
         n25275, n25276, n25277, n25278, n25279, n25280, n25281, n25282,
         n25283, n25284, n25285, n25286, n25287, n25288, n25289, n25290,
         n25291, n25292, n25293, n25294, n25295, n25296, n25297, n25298,
         n25299, n25300, n25301, n25302, n25303, n25304, n25305, n25306,
         n25307, n25308, n25309, n25310, n25311, n25312, n25313, n25314,
         n25315, n25316, n25317, n25318, n25319, n25320, n25321, n25322,
         n25323, n25325, n25326, n25327, n25328, n25329, n25330, n25331,
         n25332, n25333, n25334, n25335, n25336, n25337, n25338, n25339,
         n25340, n25342, n25343, n25344, n25345, n25346, n25347, n25348,
         n25349, n25350, n25351, n25352, n25353, n25354, n25355, n25356,
         n25357, n25358, n25359, n25360, n25361, n25362, n25364, n25365,
         n25367, n25368, n25369, n25370, n25371, n25372, n25373, n25374,
         n25375, n25376, n25377, n25378, n25379, n25380, n25381, n25382,
         n25383, n25384, n25385, n25386, n25387, n25388, n25389, n25390,
         n25391, n25392, n25393, n25394, n25395, n25396, n25397, n25398,
         n25399, n25401, n25402, n25403, n25404, n25405, n25406, n25407,
         n25408, n25409, n25410, n25411, n25412, n25413, n25414, n25415,
         n25416, n25417, n25419, n25420, n25421, n25422, n25423, n25424,
         n25425, n25426, n25427, n25428, n25429, n25430, n25431, n25432,
         n25433, n25434, n25435, n25436, n25437, n25438, n25439, n25440,
         n25441, n25443, n25444, n25445, n25446, n25447, n25448, n25449,
         n25450, n25451, n25452, n25453, n25454, n25455, n25456, n25457,
         n25458, n25459, n25460, n25461, n25463, n25464, n25465, n25466,
         n25467, n25468, n25469, n25470, n25471, n25472, n25473, n25474,
         n25475, n25476, n25477, n25478, n25479, n25480, n25482, n25483,
         n25484, n25486, n25487, n25488, n25489, n25490, n25491, n25492,
         n25493, n25494, n25495, n25496, n25497, n25498, n25499, n25500,
         n25501, n25502, n25503, n25504, n25506, n25507, n25508, n25510,
         n25511, n25512, n25513, n25514, n25515, n25516, n25517, n25518,
         n25519, n25520, n25521, n25522, n25523, n25524, n25525, n25526,
         n25527, n25528, n25530, n25531, n25532, n25534, n25535, n25536,
         n25537, n25538, n25539, n25540, n25541, n25542, n25543, n25544,
         n25545, n25548, n25549, n25550, n25551, n25552, n25553, n25555,
         n25556, n25557, n25558, n25560, n25561, n25562, n25563, n25564,
         n25565, n25566, n25567, n25568, n25569, n25570, n25571, n25572,
         n25573, n25574, n25575, n25576, n25577, n25578, n25579, n25580,
         n25581, n25582, n25583, n25584, n25585, n25586, n25587, n25588,
         n25589, n25590, n25591, n25592, n25593, n25594, n25595, n25596,
         n25597, n25598, n25599, n25600, n25601, n25602, n25603, n25604,
         n25605, n25606, n25607, n25608, n25609, n25610, n25611, n25612,
         n25613, n25614, n25615, n25616, n25617, n25618, n25619, n25620,
         n25621, n25622, n25623, n25624, n25625, n25626, n25627, n25628,
         n25629, n25630, n25631, n25632, n25635, n25637, n25638, n25639,
         n25640, n25643, n25644, n25645, n25646, n25647, n25648, n25649,
         n25650, n25651, n25652, n25653, n25654, n25677, n25678, n25679,
         n25680, n25681, n25683, n25684, n25685, n25686, n25696, n25697,
         n25698, n25699, n25741, n25742, n25743, n25744, n25786, n25788,
         n25789, n25790, n25791, n25792, n25795, n25796, n25797, n25798,
         n25807, n25808, n25811, n25812, n25813, n25814, n25819, n25820,
         n25821, n25822, n25823, n25824, n25829, n25830, n25831, n25832,
         n25833, n25834, n25839, n25840, n25841, n25842, n25843, n25844,
         n25849, n25850, n25851, n25852, n25853, n25854, n25855, n25856,
         n25857, n25858, n25859, n25860, n25861, n25862, n25864, n25865,
         n25866, n25867, n25868, n25869, n25870, n25871, n25872, n25873,
         n25874, n25875, n25876, n25877, n25878, n25885, n25886, n25887,
         n25888, n25895, n25896, n25897, n25898, n25899, n25900, n25901,
         n25902, n25903, n25904, n25905, n25906, n25907, n25908, n25909,
         n25914, n25915, n25916, n25917, n25918, n25919, n25926, n25927,
         n25928, n25929, n25936, n25937, n25938, n25939, n25946, n25947,
         n25948, n25949, n25954, n25955, n25956, n25957, n25958, n25959,
         n25966, n25967, n25968, n25969, n25976, n25977, n25978, n25979,
         n25986, n25987, n25988, n25989, n25996, n25997, n25998, n25999,
         n26004, n26005, n26006, n26007, n26008, n26009, n26010, n26011,
         n26012, n26013, n26014, n26015, n26016, n26017, n26018, n26019,
         n26020, n26025, n26026, n26027, n26028, n26029, n26030, n26037,
         n26038, n26039, n26040, n26047, n26048, n26049, n26050, n26055,
         n26056, n26057, n26058, n26059, n26060, n26067, n26068, n26069,
         n26070, n26077, n26078, n26079, n26080, n26087, n26088, n26089,
         n26090, n26097, n26098, n26099, n26100, n26105, n26106, n26107,
         n26108, n26109, n26110, n26115, n26116, n26117, n26118, n26119,
         n26120, n26121, n26122, n26123, n26124, n26125, n26126, n26127,
         n26128, n26129, n26130, n26131, n26132, n26133, n26134, n26135,
         n26138, n26139, n26140, n26159, n26160, n26161, n26162, n26164,
         n26165, n26166, n26173, n26174, n26175, n26206, n26207, n26208,
         n26241, n26242, n26244, n26245, n26246, n26249, n26250, n26251,
         n26252, n26253, n26254, n26255, n26256, n26257, n26258, n26261,
         n26262, n26263, n26264, n26265, n26266, n26267, n26268, n26269,
         n26270, n26272, n26277, n26278, n26279, n26280, n26281, n26282,
         n26283, n26285, n26286, n26287, n26289, n26290, n26291, n26292,
         n26293, n26294, n26295, n26296, n26297, n26298, n26299, n26304,
         n26306, n26307, n26312, n26313, n26314, n26315, n26318, n26319,
         n26320, n26321, n26323, n26324, n26325, n26326, n26327, n26328,
         n26329, n26331, n26335, n26360, n26361, n26373, n26456, n26714,
         n26855, n26856, n26905, n26906, n26907, n26908, n26909, n26910,
         n26911, n26912, n26913, n26914, n26916, n26917, n26920, n26928,
         n26931, n26932, n26933, n26934, n26935, n26936, n26937, n26939,
         n26940, n26941, n26942, n26943, n26944, n26946, n26947, n26949,
         n26950, n26951, n26952, n26953, n26954, n26955, n26957, n26958,
         n26959, n26960, n26961, n26962, n26963, n26964, n26965, n26966,
         n26967, n26968, n26969, n26970, n26971, n26972, n26973, n26974,
         n26976, n26977, n26978, n26979, n26980, n26981, n26982, n26983,
         n26984, n26985, n26986, n26988, n26989, n26990, n26991, n26992,
         n26993, n26994, n26995, n26997, n26998, n27018, n27019, n27022,
         n27031, n27064, n27095, n27096, n27100, n27101, n27102, n27104,
         n27122, n27123, n27124, n27125, n27126, n27127, n27128, n27135,
         n27136, n27137, n27168, n27169, n27170, n27201, n27202, n27203,
         n27205, n27206, n27207, n27208, n27226, n27227, n27228, n27229,
         n27230, n27231, n27232, n27239, n27240, n27241, n27272, n27273,
         n27274, n27305, n27306, n27307, n27308, n27309, n27310, n27311,
         n27312, n27313, n27314, n27315, n27316, n27317, n27318, n27319,
         n27320, n27321, n27322, n27323, n27324, n27325, n27326, n27327,
         n27328, n27329, n27330, n27331, n27332, n27335, n27336, n27338,
         n27339, n27340, n27342, n27343, n27344, n27345, n27346, n27347,
         n27349, n27350, n27351, n27352, n27353, n27355, n27356, n27357,
         n27358, n27359, n27360, n27361, n27362, n27363, n27364, n27367,
         n27368, n27369, n27370, n27371, n27373, n27374, n27376, n27377,
         n27378, n27379, n27380, n27381, n27382, n27383, n27384, n27385,
         n27386, n27387, n27388, n27389, n27390, n27391, n27392, n27393,
         n27394, n27395, n27398, n27399, n27400, n27401, n27402, n27403,
         n27407, n27420, n27421, n27422, n27423, n27424, n27425, n27426,
         n27427, n27428, n27429, n27430, n27431, n27432, n27433, n27434,
         n27435, n27436, n27461, n27462, n27463, n27464, n27465, n27477,
         n27560, n27960, n27961, n27964, n28010, n28011, n28012, n28013,
         n28014, n28015, n28031, n28032, n28034, n28035, n28045, n28056,
         n28057, n28058, n28059, n28060, n28061, n28062, n28064, n28065,
         n28066, n28067, n28068, n28069, n28070, n28071, n28072, n28091,
         n28092, n28093, n28094, n28095, n28096, n28097, n28098, n28100,
         n28101, n28102, n28103, n28104, n28105, n28106, n28107, n28108,
         n28109, n28110, n28111, n28112, n28113, n28114, n28115, n28116,
         n28117, n28118, n28119, n28120, n28121, n28122, n28123, n28124,
         n28125, n28126, n28127, n28128, n28129, n28130, n28131, n28132,
         n28133, n28134, n28135, n28136, n28137, n28138, n28139, n28140,
         n28141, n28142, n28143, n28144, n28145, n28146, n28147, n28148,
         n28149, n28151, n28153, n28154, n28155, n28156, n28157, n28158,
         n28161, n28162, n28163, n28164, n28165, n28166, n28169, n28170,
         n28171, n28172, n28174, n28175, n28176, n28177, n28178, n28179,
         n28180, n28181, n28182, n28183, n28184, n28185, n28186, n28187,
         n28188, n28189, n28190, n28191, n28192, n28193, n28194, n28195,
         n28196, n28202, n28203, n28204, n28205, n28206, n28207, n28208,
         n28209, n28210, n28211, n28212, n28213, n28214, n28215, n28220,
         n28221, n28222, n28223, n28224, n28225, n28227, n28228, n28229,
         n28230, n28231, n28232, n28233, n28234, n28235, n28236, n28237,
         n28238, n28239, n28240, n28241, n28243, n28244, n28245, n28246,
         n28247, n28249, n28252, n28256, n28259, n28262, n28263, n28264,
         n28268, n28270, n28272, n28273, n28276, n28278, n28280, n28281,
         n28284, n28286, n28288, n28289, n28292, n28294, n28296, n28297,
         n28300, n28302, n28304, n28305, n28308, n28310, n28312, n28313,
         n28316, n28318, n28320, n28321, n28324, n28326, n28328, n28329,
         n28332, n28334, n28336, n28337, n28340, n28342, n28344, n28345,
         n28348, n28350, n28352, n28353, n28356, n28358, n28360, n28361,
         n28364, n28366, n28368, n28369, n28372, n28374, n28376, n28377,
         n28380, n28382, n28384, n28385, n28388, n28390, n28392, n28393,
         n28396, n28398, n28400, n28401, n28404, n28406, n28408, n28409,
         n28412, n28414, n28416, n28417, n28420, n28422, n28424, n28425,
         n28428, n28430, n28432, n28433, n28436, n28438, n28440, n28441,
         n28444, n28446, n28448, n28449, n28452, n28454, n28456, n28457,
         n28460, n28462, n28464, n28465, n28468, n28470, n28472, n28473,
         n28476, n28478, n28480, n28481, n28484, n28486, n28488, n28489,
         n28492, n28494, n28496, n28497, n28500, n28502, n28504, n28505,
         n28508, n28510, n28512, n28515, n28516, n28517, n28518, n28519,
         n28520, n28521, n28522, n28523, n28524, n28525, n28526, n28527,
         n28528, n28529, n28530, n28531, n28532, n28533, n28536, n28537,
         n28538, n28539, n28540, n28541, n28542, n28543, n28544, n28545,
         n28546, n28547, n28549, n28550, n28551, n28558, n28560, n28561,
         n28562, n28563, n28567, n28578, n28579, n28582, n28607, n28608,
         n28610, n28611, n28612, n28613, n28616, n28617, n28618, n28619,
         n28620, n28621, n28624, n28625, n28626, n28627, n28628, n28629,
         n28632, n28633, n28636, n28734, n28735, n28736, n28737, n28738,
         n28739, n28740, n28741, n28742, n28743, n28744, n28745, n28765,
         n28776, n28777, n28778, n28779, n28780, n28781, n28782, n28783,
         n28784, n28785, n28786, n28787, n28788, n28789, n28790, n28791,
         n28796, n28797, n28813, n28814, n28815, n28816, n28817, n28818,
         n28819, n28820, n28821, n28822, n28823, n28824, n28825, n28826,
         n28827, n28828, n28829, n28830, n28831, n28832, n28833, n28834,
         n28835, n28836, n28837, n28838, n28839, n28840, n28841, n28842,
         n28843, n28844, n28845, n28846, n28847, n28848, n28905, n28907,
         n28908, n28909, n28910, n28911, n28913, n28932, n28933, n28934,
         n28941, n28942, n28943, n28944, n28945, n28946, n28947, n28948,
         n28949, n28953, n28982, n28996, n29013, n29026, n29027, n29028,
         n29029, n29030, n29031, n29032, n29033, n29034, n29035, n29036,
         n29037, n29040, n29041, n29042, n29043, n29044, n29045, n29046,
         n29047, n29048, n29049, n29053, n29054, n29055, n29056, n29057,
         n29058, n29059, n29060, n29061, n29062, n29063, n29064, n29067,
         n29068, n29069, n29070, n29071, n29072, n29073, n29074, n29075,
         n29076, n29079, n29080, n29081, n29082, n29083, n29084, n29085,
         n29086, n29087, n29088, n29089, n29090, n29093, n29094, n29095,
         n29096, n29097, n29098, n29099, n29100, n29101, n29102, n29103,
         n29104, n29105, n29106, n29107, n29108, n29109, n29110, n29111,
         n29112, n29113, n29114, n29115, n29116, n29117, n29118, n29119,
         n29120, n29122, n29123, n29124, n29125, n29126, n29127, n29128,
         n29129, n29130, n29132, n29133, n29134, n29135, n29136, n29137,
         n29138, n29139, n29140, n29141, n29144, n29145, n29146, n29147,
         n29148, n29149, n29151, n29152, n29153, n29156, n29157, n29158,
         n29159, n29160, n29161, n29162, n29163, n29164, n29167, n29168,
         n29169, n29170, n29171, n29172, n29173, n29174, n29176, n29177,
         n29178, n29179, n29180, n29181, n29182, n29183, n29184, n29187,
         n29188, n29189, n29190, n29191, n29192, n29193, n29194, n29197,
         n29198, n29199, n29200, n29201, n29202, n29203, n29204, n29205,
         n29207, n29208, n29209, n29210, n29211, n29212, n29213, n29214,
         n29215, n29216, n29217, n29218, n29219, n29220, n29221, n29222,
         n29223, n29224, n29225, n29226, n29227, n29228, n29229, n29230,
         n29231, n29232, n29233, n29234, n29235, n29236, n29237, n29238,
         n29239, n29240, n29241, n29242, n29243, n29244, n29245, n29246,
         n29247, n29248, n29249, n29250, n29251, n29252, n29253, n29254,
         n29255, n29256, n29257, n29258, n29259, n29260, n29261, n29262,
         n29263, n29264, n29265, n29266, n29267, n29268, n29269, n29270,
         n29271, n29272, n29273, n29274, n29275, n29276, n29277, n29278,
         n29279, n29280, n29281, n29282, n29283, n29284, n29285, n29286,
         n29287, n29288, n29289, n29290, n29291, n29292, n29293, n29294,
         n29295, n29298, n29299, n29300, n29301, n29302, n29303, n29304,
         n29305, n29306, n29308, n29309, n29310, n29311, n29312, n29313,
         n29314, n29315, n29316, n29317, n29318, n29320, n29321, n29322,
         n29323, n29324, n29325, n29326, n29327, n29328, n29329, n29330,
         n29332, n29333, n29334, n29335, n29336, n29337, n29338, n29339,
         n29340, n29341, n29343, n29344, n29345, n29346, n29347, n29348,
         n29349, n29350, n29351, n29352, n29354, n29371, n29372, n29373,
         n29374, n29375, n29376, n29377, n29378, n29379, n29380, n29381,
         n29382, n29383, n29384, n29385, n29386, n29387, n29388, n29389,
         n29390, n29391, n29392, n29393, n29394, n29395, n29396, n29397,
         n29398, n29399, n29400, n29401, n29402, n29403, n29404, n29405,
         n29406, n29407, n29408, n29409, n29410, n29411, n29412, n29413,
         n29414, n29415, n29416, n29417, n29418, n29419, n29420, n29421,
         n29422, n29424, n29425, n29426, n29427, n29428, n29429, n29430,
         n29431, n29432, n29433, n29434, n29435, n29436, n29437, n29438,
         n29440, n29441, n29442, n29443, n29444, n29445, n29446, n29447,
         n29448, n29449, n29450, n29451, n29452, n29453, n29454, n29456,
         n29457, n29458, n29459, n29460, n29461, n29462, n29463, n29464,
         n29465, n29466, n29467, n29468, n29469, n29470, n29472, n29473,
         n29474, n29475, n29476, n29477, n29478, n29479, n29480, n29481,
         n29482, n29483, n29484, n29485, n29486, n29488, n29489, n29490,
         n29491, n29492, n29493, n29494, n29495, n29496, n29497, n29498,
         n29499, n29500, n29501, n29502, n29503, n29504, n29505, n29506,
         n29507, n29508, n29509, n29510, n29511, n29512, n29513, n29514,
         n29515, n29516, n29517, n29518, n29519, n29520, n29521, n29522,
         n29523, n29524, n29525, n29526, n29527, n29528, n29529, n29530,
         n29531, n29532, n29533, n29534, n29535, n29536, n29537, n29538,
         n29539, n29544, n29545, n29546, n29547, n29549, n29550, n29551,
         n29552, n29553, n29554, n29555, n29556, n29557, n29558, n29559,
         n29560, n29561, n29562, n29563, n29564, n29567, n29568, n29569,
         n29570, n29571, n29574, n29575, n29576, n29577, n29578, n29579,
         n29580, n29581, n29582, n29583, n29584, n29585, n29586, n29587,
         n29588, n29589, n29590, n29591, n29592, n29593, n29594, n29595,
         n29596, n29597, n29598, n29599, n29600, n29601, n29602, n29603,
         n29604, n29605, n29606, n29607, n29608, n29609, n29610, n29611,
         n29612, n29613, n29614, n29615, n29620, n29621, n29622, n29623,
         n29627, n29628, n29629, n29630, n29631, n29632, n29633, n29634,
         n29640, n29643, n29644, n29645, n29646, n29647, n29649, n29650,
         n29651, n29652, n29653, n29654, n29655, n29657, n29664, n29665,
         n29669, n29670, n29671, n29673, n29674, n29675, n29677, n29680,
         n29681, n29682, n29690, n29691, n29692, n29701, n29702, n29703,
         n29704, n29712, n29713, n29714, n29722, n29723, n29724, n29725,
         n29733, n29734, n29735, n29743, n29744, n29745, n29746, n29754,
         n29755, n29756, n29764, n29765, n29766, n29767, n29776, n29777,
         n29786, n29787, n29788, n29929, n29930, n29931, n29939, n29940,
         n29941, n29942, n29961, n29963, n29964, n29965, n29966, n29967,
         n29968, n29971, n29972, n29973, n29974, n29975, n29976, n29977,
         n29978, n29979, n29980, n29981, n29982, n29983, n29984, n29985,
         n29986, n29987, n29988, n29989, n29990, n29991, n29992, n29993,
         n29994, n29995, n29996, n29997, n29998, n30003, n30004, n30005,
         n30007, n30008, n30009, n30010, n30011, n30012, n30013, n30014,
         n30015, n30016, n30017, n30018, n30019, n30020, n30021, n30023,
         n30024, n30025, n30026, n30027, n30028, n30031, n30032, n30033,
         n30034, n30037, n30038, n30039, n30040, n30041, n30042, n30043,
         n30044, n30045, n30047, n30048, n30049, n30050, n30051, n30053,
         n30054, n30055, n30056, n30057, n30061, n30062, n30063, n30064,
         n30067, n30068, n30069, n30070, n30071, n30072, n30073, n30074,
         n30075, n30076, n30077, n30078, n30079, n30080, n30081, n30082,
         n30085, n30086, n30087, n30088, n30093, n30094, n30095, n30096,
         n30097, n30098, n30099, n30100, n30105, n30106, n30109, n30110,
         n30111, n30112, n30113, n30114, n30117, n30118, n30123, n30124,
         n30125, n30126, n30127, n30128, n30129, n30130, n30131, n30132,
         n30271, n30272, n30273, n30274, n30317, n30318, n30319, n30327,
         n30328, n30329, n30330, n30403, n30413, n30414, n30426, n30429,
         n30435, n30436, n30445, n30455, n30456, n30469, n30470, n30471,
         n30479, n30480, n30481, n30482, n30493, n30494, n30495, n30504,
         n30505, n30513, n30514, n30515, n30523, n30524, n30525, n30526,
         n30544, n30545, n30546, n30547, n30548, n30549, n30558, n30559,
         n30560, n30561, n30569, n30570, n30571, n30572, n30573, n30574,
         n30575, n30583, n30584, n30585, n30586, n30594, n30595, n30596,
         n30604, n30605, n30606, n30607, n30616, n30617, n30618, n30619,
         n30620, n30621, n30622, n30623, n30624, n30632, n30633, n30634,
         n30635, n30636, n30637, n30708, n30709, n30710, n30711, n30771,
         n30772, n30773, n30774, n30775, n30776, n30820, n30821, n30822,
         n30823, n30824, n30825, n31124, n31128, n31129, n31132, n31133,
         n31134, n31135, n31136, n31137, n31138, n31139, n31144, n31145,
         n31146, n31147, n31148, n31149, n31150, n31151, n31152, n31153,
         n31154, n31155, n31156, n31158, n31159, n31160, n31161, n31162,
         n31163, n31164, n31165, n31176, n31177, n31178, n31179, n31182,
         n31183, n31184, n31185, n31186, n31187, n31198, n31199, n31200,
         n31201, n31204, n31205, n31206, n31207, n31208, n31209, n31220,
         n31221, n31222, n31223, n31226, n31227, n31228, n31229, n31230,
         n31231, n31242, n31243, n31244, n31245, n31248, n31249, n31250,
         n31251, n31252, n31253, n31264, n31265, n31266, n31267, n31268,
         n31269, n31270, n31271, n31272, n31273, n31274, n31275, n31276,
         n31277, n31278, n31279, n31280, n31281, n31282, n31283, n31289,
         n31302, n31303, n31308, n31309, n31316, n31317, n31322, n31323,
         n31330, n31331, n31337, n31338, n31343, n31344, n31351, n31352,
         n31357, n31358, n31363, n31364, n31371, n31372, n31377, n31378,
         n31383, n31384, n31391, n31393, n31394, n31395, n31400, n31401,
         n31408, n31409, n31410, n31411, n31412, n31423, n31424, n31444,
         n31445, n31450, n31451, n31460, n31461, n31462, n31463, n31464,
         n31465, n31653, n31654, n31786, n31787, n31921, n31922, n31923,
         n32007, n32008, n32009, n32010, n32011, n32196, n32197, n32198,
         n32199, n32333, n32335, n32467, n32468, n32471, n32472, n32473,
         n32474, n32475, n32476, n32477, n32610, n32743, n32744, n33270,
         n33271, n33539, n33540, n33541, n33542, n33543, n33676, n33677,
         n33678, n33679, n33680, n33681, n34080, n34081, n34082, n34083,
         n34084, n34085, n34086, n34087, n34221, n34356, n34489, n34490,
         n34491, n34492, n34625, n34758, n34759, n34760, n34761, n35026,
         n35027, n35028, n35029, n35030, n35031, n35165, n35166, n35167,
         n35168, n35303, n35304, n35305, n35306, n35307, n35308, n35309,
         n35310, n35311, n35312, n35891, n35892, n35893, n35894, n35895,
         n35896, n35897, n35898, n35899, n35900, n35901, n35902, n35903,
         n35904, n35905, n35906, n35922, n35938, n35945, n35952, n35956,
         n35957, n35958, n35959, n35970, n35981, n35982, n35983, n35987,
         n35988, n35989, n35990, n35991, n35997, n35999, n36000, n36001,
         n36002, n36006, n36009, n36163, n36175, n36176, n36177, n36178,
         n36180, n36191, n36197, n36198, n36199, n36200, n36202, n36207,
         n36208, n36209, n36210, n36211, n36212, n36217, n36219, n36220,
         n36221, n36227, n36228, n36237, n36238, n36239, n36240, n36244,
         n36247, n36248, n36249, n36250, n36251, n36340, n36341, n36342,
         n36343, n36344, \clk_gate_u_mmu_dtlb_entry_q_reg/n2 ,
         \clk_gate_u_mmu_dtlb_entry_q_reg_0/n2 ,
         \clk_gate_u_mmu_itlb_entry_q_reg/n2 ,
         \clk_gate_u_mmu_itlb_entry_q_reg_0/n2 ,
         \clk_gate_u_mmu_pte_entry_q_reg/n2 ,
         \clk_gate_u_mmu_pte_addr_q_reg/n2 ,
         \clk_gate_u_mmu_pte_addr_q_reg_0/n2 ,
         \clk_gate_u_mmu_virt_addr_q_reg/n2 ,
         \clk_gate_u_mmu_lsu_in_addr_q_reg/n2 ,
         \clk_gate_u_mmu_lsu_in_addr_q_reg_0/n2 ,
         \clk_gate_u_lsu_mem_cacheable_q_reg/n2 ,
         \clk_gate_u_lsu_mem_addr_q_reg/n2 ,
         \clk_gate_u_lsu_mem_addr_q_reg_0/n2 ,
         \clk_gate_u_lsu_mem_data_wr_q_reg/n2 ,
         \clk_gate_u_lsu_mem_data_wr_q_reg_0/n2 ,
         \clk_gate_u_csr_writeback_value_q_reg/n2 ,
         \clk_gate_u_csr_writeback_value_q_reg_0/n2 ,
         \clk_gate_u_csr_writeback_idx_q_reg/n2 ,
         \clk_gate_u_csr_pc_m_q_reg/n2 , \clk_gate_u_csr_csr_sr_q_reg/n2 ,
         \clk_gate_u_muldiv_divisor_q_reg/n2 ,
         \clk_gate_u_muldiv_divisor_q_reg_0/n2 ,
         \clk_gate_u_muldiv_divisor_q_reg_1/n2 ,
         \clk_gate_u_muldiv_divisor_q_reg_2/n2 ,
         \clk_gate_u_muldiv_q_mask_q_reg/n2 ,
         \clk_gate_u_muldiv_dividend_q_reg/n2 ,
         \clk_gate_u_muldiv_dividend_q_reg_0/n2 ,
         \clk_gate_u_muldiv_quotient_q_reg/n2 ,
         \clk_gate_u_muldiv_quotient_q_reg_0/n2 ,
         \clk_gate_u_decode_opcode_instr_q_reg/n2 ,
         \clk_gate_u_decode_opcode_instr_q_reg_0/n2 ,
         \clk_gate_u_decode_opcode_instr_q_reg_1/n2 ,
         \clk_gate_u_decode_opcode_instr_q_reg_2/n2 ,
         \clk_gate_u_decode_inst_q_reg/n2 , \clk_gate_u_decode_pc_q_reg/n2 ,
         \clk_gate_u_decode_pc_q_reg_0/n2 ,
         \clk_gate_u_decode_u_regfile_reg_r21_q_reg/n2 ,
         \clk_gate_u_decode_u_regfile_reg_r21_q_reg_0/n2 ,
         \clk_gate_u_decode_u_regfile_reg_r20_q_reg/n2 ,
         \clk_gate_u_decode_u_regfile_reg_r20_q_reg_0/n2 ,
         \clk_gate_u_decode_u_regfile_reg_r19_q_reg/n2 ,
         \clk_gate_u_decode_u_regfile_reg_r19_q_reg_0/n2 ,
         \clk_gate_u_decode_u_regfile_reg_r18_q_reg/n2 ,
         \clk_gate_u_decode_u_regfile_reg_r18_q_reg_0/n2 ,
         \clk_gate_u_decode_u_regfile_reg_r17_q_reg/n2 ,
         \clk_gate_u_decode_u_regfile_reg_r17_q_reg_0/n2 ,
         \clk_gate_u_decode_u_regfile_reg_r16_q_reg/n2 ,
         \clk_gate_u_decode_u_regfile_reg_r16_q_reg_0/n2 ,
         \clk_gate_u_decode_u_regfile_reg_r15_q_reg/n2 ,
         \clk_gate_u_decode_u_regfile_reg_r15_q_reg_0/n2 ,
         \clk_gate_u_decode_u_regfile_reg_r14_q_reg/n2 ,
         \clk_gate_u_decode_u_regfile_reg_r14_q_reg_0/n2 ,
         \clk_gate_u_decode_u_regfile_reg_r13_q_reg/n2 ,
         \clk_gate_u_decode_u_regfile_reg_r13_q_reg_0/n2 ,
         \clk_gate_u_decode_u_regfile_reg_r12_q_reg/n2 ,
         \clk_gate_u_decode_u_regfile_reg_r12_q_reg_0/n2 ,
         \clk_gate_u_decode_u_regfile_reg_r11_q_reg/n2 ,
         \clk_gate_u_decode_u_regfile_reg_r11_q_reg_0/n2 ,
         \clk_gate_u_decode_u_regfile_reg_r10_q_reg/n2 ,
         \clk_gate_u_decode_u_regfile_reg_r10_q_reg_0/n2 ,
         \clk_gate_u_decode_u_regfile_reg_r9_q_reg/n2 ,
         \clk_gate_u_decode_u_regfile_reg_r9_q_reg_0/n2 ,
         \clk_gate_u_decode_u_regfile_reg_r8_q_reg/n2 ,
         \clk_gate_u_decode_u_regfile_reg_r8_q_reg_0/n2 ,
         \clk_gate_u_decode_u_regfile_reg_r7_q_reg/n2 ,
         \clk_gate_u_decode_u_regfile_reg_r7_q_reg_0/n2 ,
         \clk_gate_u_decode_u_regfile_reg_r6_q_reg/n2 ,
         \clk_gate_u_decode_u_regfile_reg_r6_q_reg_0/n2 ,
         \clk_gate_u_decode_u_regfile_reg_r5_q_reg/n2 ,
         \clk_gate_u_decode_u_regfile_reg_r5_q_reg_0/n2 ,
         \clk_gate_u_decode_u_regfile_reg_r4_q_reg/n2 ,
         \clk_gate_u_decode_u_regfile_reg_r4_q_reg_0/n2 ,
         \clk_gate_u_decode_u_regfile_reg_r3_q_reg/n2 ,
         \clk_gate_u_decode_u_regfile_reg_r3_q_reg_0/n2 ,
         \clk_gate_u_decode_u_regfile_reg_r2_q_reg/n2 ,
         \clk_gate_u_decode_u_regfile_reg_r2_q_reg_0/n2 ,
         \clk_gate_u_decode_u_regfile_reg_r1_q_reg/n2 ,
         \clk_gate_u_decode_u_regfile_reg_r1_q_reg_0/n2 ,
         \clk_gate_u_decode_u_regfile_reg_r31_q_reg/n2 ,
         \clk_gate_u_decode_u_regfile_reg_r31_q_reg_0/n2 ,
         \clk_gate_u_decode_u_regfile_reg_r26_q_reg/n2 ,
         \clk_gate_u_decode_u_regfile_reg_r26_q_reg_0/n2 ,
         \clk_gate_u_decode_u_regfile_reg_r27_q_reg/n2 ,
         \clk_gate_u_decode_u_regfile_reg_r27_q_reg_0/n2 ,
         \clk_gate_u_decode_u_regfile_reg_r25_q_reg/n2 ,
         \clk_gate_u_decode_u_regfile_reg_r25_q_reg_0/n2 ,
         \clk_gate_u_decode_u_regfile_reg_r28_q_reg/n2 ,
         \clk_gate_u_decode_u_regfile_reg_r28_q_reg_0/n2 ,
         \clk_gate_u_decode_u_regfile_reg_r24_q_reg/n2 ,
         \clk_gate_u_decode_u_regfile_reg_r24_q_reg_0/n2 ,
         \clk_gate_u_decode_u_regfile_reg_r29_q_reg/n2 ,
         \clk_gate_u_decode_u_regfile_reg_r29_q_reg_0/n2 ,
         \clk_gate_u_decode_u_regfile_reg_r23_q_reg/n2 ,
         \clk_gate_u_decode_u_regfile_reg_r23_q_reg_0/n2 ,
         \clk_gate_u_decode_u_regfile_reg_r30_q_reg/n2 ,
         \clk_gate_u_decode_u_regfile_reg_r30_q_reg_0/n2 ,
         \clk_gate_u_decode_u_regfile_reg_r22_q_reg/n2 ,
         \clk_gate_u_decode_u_regfile_reg_r22_q_reg_0/n2 ,
         \clk_gate_u_fetch_pc_d_q_reg/n2 , \clk_gate_u_fetch_pc_d_q_reg_0/n2 ,
         \clk_gate_u_fetch_branch_pc_q_reg/n2 ,
         \clk_gate_u_fetch_branch_pc_q_reg_0/n2 ,
         \clk_gate_u_fetch_fetch_pc_q_reg/n2 ,
         \clk_gate_u_fetch_fetch_pc_q_reg_0/n2 ,
         \clk_gate_u_fetch_skid_buffer_q_reg/n2 ,
         \clk_gate_u_fetch_skid_buffer_q_reg_0/n2 ,
         \clk_gate_u_fetch_skid_buffer_q_reg_1/n2 ,
         \clk_gate_u_fetch_skid_buffer_q_reg_2/n2 , n36346, n36347, n36348,
         n36349, n36350, n36351, n36352, n36353, n36354, n36355, n36356,
         n36357, n36358, n36359, n36360, n36361, n36362, n36363, n36364,
         n36365, n36366, n36367, n36368, n36369, n36370, n36371, n36372,
         n36373, n36374, n36375, n36376, n36377, n36378, n36379, n36380,
         n36381, n36382, n36383, n36384, n36385, n36386, n36387, n36388,
         n36389, n36390, n36391, n36392, n36393, n36394, n36395, n36396,
         n36397, n36398, n36399, n36400, n36401, n36402, n36403, n36404,
         n36405, n36406, n36407, n36408, n36409, n36410, n36411, n36412,
         n36413, n36414, n36415, n36416, n36417, n36418, n36419, n36420,
         n36421, n36422, n36423, n36424, n36425, n36426, n36427, n36428,
         n36429, n36430, n36431, n36432, n36433, n36434, n36435, n36436,
         n36437, n36438, n36439, n36440, n36441, n36442, n36443, n36444,
         n36445, n36446, n36447, n36448, n36449, n36450, n36451, n36452,
         n36453, n36454, n36455, n36456, n36457, n36458, n36459, n36460,
         n36461, n36462, n36463, n36464, n36465, n36466, n36467, n36468,
         n36469, n36470, n36471, n36472, n36473, n36474, n36475, n36476,
         n36477, n36478, n36479, n36480, n36481, n36482, n36483, n36484,
         n36485, n36486, n36487, n36488, n36489, n36490, n36491, n36492,
         n36493, n36494, n36495, n36496, n36497, n36498, n36499, n36500,
         n36501, n36502, n36503, n36504, n36505, n36506, n36507, n36508,
         n36509, n36510, n36511, n36512, n36513, n36514, n36515, n36516,
         n36517, n36518, n36519, n36520, n36521, n36522, n36523, n36524,
         n36525, n36526, n36527, n36528, n36529, n36530, n36531, n36532,
         n36533, n36534, n36535, n36536, n36537, n36538, n36539, n36540,
         n36541, n36542, n36543, n36544, n36545, n36546, n36547, n36548,
         n36549, n36550, n36551, n36552, n36553, n36554, n36555, n36556,
         n36557, n36558, n36559, n36560, n36561, n36562, n36563, n36564,
         n36565, n36566, n36567, n36568, n36569, n36570, n36571, n36572,
         n36573, n36574, n36575, n36576, n36577, n36578, n36579, n36580,
         n36581, n36582, n36583, n36584, n36585, n36586, n36587, n36588,
         n36589, n36590, n36591, n36592, n36593, n36594, n36595, n36596,
         n36597, n36598, n36599, n36600, n36601, n36602, n36603, n36604,
         n36605, n36606, n36607, n36608, n36609, n36610, n36611, n36612,
         n36613, n36614, n36615, n36616, n36617, n36618, n36619, n36620,
         n36621, n36622, n36623, n36624, n36625, n36626, n36627, n36628,
         n36629, n36630, n36631, n36632, n36633, n36634, n36635, n36636,
         n36637, n36638, n36639, n36640, n36641, n36642, n36643, n36644,
         n36645, n36646, n36647, n36648, n36649, n36650, n36651, n36652,
         n36653, n36654, n36655, n36656, n36657, n36658, n36659, n36660,
         n36661, n36662, n36663, n36664, n36665, n36666, n36667, n36668,
         n36669, n36670, n36671, n36672, n36673, n36674, n36675, n36676,
         n36677, n36678, n36679, n36680, n36681, n36682, n36683, n36684,
         n36685, n36686, n36687, n36688, n36689, n36690, n36691, n36692,
         n36693, n36694, n36695, n36696, n36697, n36698, n36699, n36700,
         n36701, n36702, n36703, n36704, n36705, n36706, n36707, n36708,
         n36709, n36710, n36711, n36712, n36713, n36714, n36715, n36716,
         n36717, n36718, n36719, n36720, n36721, n36722, n36723, n36724,
         n36725, n36726, n36727, n36728, n36729, n36730, n36731, n36732,
         n36733, n36734, n36735, n36736, n36737, n36738, n36739, n36740,
         n36741, n36742, n36743, n36744, n36745, n36746, n36747, n36748,
         n36749, n36750, n36751, n36752, n36753, n36754, n36755, n36756,
         n36757, n36758, n36759, n36760, n36761, n36762, n36763, n36764,
         n36765, n36766, n36767, n36768, n36769, n36770, n36771, n36772,
         n36773, n36774, n36775, n36776, n36777, n36778, n36779, n36780,
         n36781, n36782, n36783, n36784, n36785, n36786, n36787, n36788,
         n36789, n36790, n36791, n36792, n36793, n36794, n36795, n36796,
         n36797, n36798, n36799, n36800, n36801, n36802, n36803, n36804,
         n36805, n36806, n36807, n36808, n36809, n36810, n36811, n36812,
         n36813, n36814, n36815, n36816, n36817, n36818, n36819, n36820,
         n36821, n36822, n36823, n36824, n36825, n36826, n36827, n36828,
         n36829, n36830, n36831, n36832, n36833, n36834, n36835, n36836,
         n36837, n36838, n36839, n36840, n36841, n36842, n36843, n36844,
         n36845, n36846, n36847, n36848, n36849, n36850, n36851, n36852,
         n36853, n36854, n36855, n36856, n36857, n36858, n36859, n36860,
         n36861, n36862, n36863, n36864, n36865, n36866, n36867, n36868,
         n36869, n36870, n36871, n36872, n36873, n36874, n36875, n36876,
         n36877, n36878, n36879, n36880, n36881, n36882, n36883, n36884,
         n36885, n36886, n36887, n36888, n36889, n36890, n36891, n36892,
         n36893, n36894, n36895, n36896, n36897, n36898, n36899, n36900,
         n36901, n36902, n36903, n36904, n36905, n36906, n36907, n36908,
         n36909, n36910, n36911, n36912, n36913, n36914, n36915, n36916,
         n36917, n36918, n36919, n36920, n36921, n36922, n36923, n36924,
         n36925, n36926, n36927, n36928, n36929, n36930, n36931, n36932,
         n36933, n36934, n36935, n36936, n36937, n36938, n36939, n36940,
         n36941, n36942, n36943, n36944, n36945, n36946, n36947, n36948,
         n36949, n36950, n36951, n36952, n36953, n36954, n36955, n36956,
         n36957, n36958, n36959, n36960, n36961, n36962, n36963, n36964,
         n36965, n36966, n36967, n36968, n36969, n36970, n36971, n36972,
         n36973, n36974, n36975, n36976, n36977, n36978, n36979, n36980,
         n36981, n36982, n36983, n36984, n36985, n36986, n36987, n36988,
         n36989, n36990, n36991, n36992, n36993, n36994, n36995, n36996,
         n36997, n36998, n36999, n37000, n37001, n37002, n37003, n37004,
         n37005, n37006, n37007, n37008, n37009, n37010, n37011, n37012,
         n37013, n37014, n37015, n37016, n37017, n37018, n37019, n37020,
         n37021, n37022, n37023, n37024, n37025, n37026, n37027, n37028,
         n37029, n37030, n37031, n37032, n37033, n37034, n37035, n37036,
         n37037, n37038, n37039, n37040, n37041, n37042, n37043, n37044,
         n37045, n37046, n37047, n37048, n37049, n37050, n37051, n37052,
         n37053, n37054, n37055, n37056, n37057, n37058, n37059, n37060,
         n37061, n37062, n37063, n37064, n37065, n37066, n37067, n37068,
         n37069, n37070, n37071, n37072, n37073, n37074, n37075, n37076,
         n37077, n37078, n37079, n37080, n37081, n37082, n37083, n37084,
         n37085, n37086, n37087, n37088, n37089, n37090, n37091, n37092,
         n37093, n37094, n37095, n37096, n37097, n37098, n37099, n37100,
         n37101, n37102, n37103, n37104, n37105, n37106, n37107, n37108,
         n37109, n37110, n37111, n37112, n37113, n37114, n37115, n37116,
         n37117, n37118, n37119, n37120, n37121, n37122, n37123, n37124,
         n37125, n37126, n37127, n37128, n37129, n37130, n37131, n37132,
         n37133, n37134, n37135, n37136, n37137, n37138, n37139, n37140,
         n37141, n37142, n37143, n37144, n37145, n37146, n37147, n37148,
         n37149, n37150, n37151, n37152, n37153, n37154, n37155, n37156,
         n37157, n37158, n37159, n37160, n37161, n37162, n37163, n37164,
         n37165, n37166, n37167, n37168, n37169, n37170, n37171, n37172,
         n37173, n37174, n37175, n37176, n37177, n37178, n37179, n37180,
         n37181, n37182, n37183, n37184, n37185, n37186, n37187, n37188,
         n37189, n37190, n37191, n37192, n37193, n37194, n37195, n37196,
         n37197, n37198, n37199, n37200, n37201, n37202, n37203, n37204,
         n37205, n37206, n37207, n37208, n37209, n37210, n37211, n37212,
         n37213, n37214, n37215, n37216, n37217, n37218, n37219, n37220,
         n37221, n37222, n37223, n37224, n37225, n37226, n37227, n37228,
         n37229, n37230, n37231, n37232, n37233, n37234, n37235, n37236,
         n37237, n37238, n37239, n37240, n37241, n37242, n37243, n37244,
         n37245, n37246, n37247, n37248, n37249, n37250, n37251, n37252,
         n37253, n37254, n37255, n37256, n37257, n37258, n37259, n37260,
         n37261, n37262, n37263, n37264, n37265, n37266, n37267, n37268,
         n37269, n37270, n37271, n37272, n37273, n37274, n37275, n37276,
         n37277, n37278, n37279, n37280, n37281, n37282, n37283, n37284,
         n37285, n37286, n37287, n37288, n37289, n37290, n37291, n37292,
         n37293, n37294, n37295, n37296, n37297, n37298, n37299, n37300,
         n37301, n37302, n37303, n37304, n37305, n37306, n37307, n37308,
         n37309, n37310, n37311, n37312, n37313, n37314, n37315, n37316,
         n37317, n37318, n37319, n37320, n37321, n37322, n37323, n37324,
         n37325, n37326, n37327, n37328, n37329, n37330, n37331, n37332,
         n37333, n37334, n37335, n37336, n37337, n37338, n37339, n37340,
         n37341, n37342, n37343, n37344, n37345, n37346, n37347, n37348,
         n37349, n37350, n37351, n37352, n37353, n37354, n37355, n37356,
         n37357, n37358, n37359, n37360, n37361, n37362, n37363, n37364,
         n37365, n37366, n37367, n37368, n37369, n37370, n37371, n37372,
         n37373, n37374, n37375, n37376, n37377, n37378, n37379, n37380,
         n37381, n37382, n37383, n37384, n37385, n37386, n37387, n37388,
         n37389, n37390, n37391, n37392, n37393, n37394, n37395, n37396,
         n37397, n37398, n37399, n37400, n37401, n37402, n37403, n37404,
         n37405, n37406, n37407, n37408, n37409, n37410, n37411, n37412,
         n37413, n37414, n37415, n37416, n37417, n37418, n37419, n37420,
         n37421, n37422, n37423, n37424, n37425, n37426, n37427, n37428,
         n37429, n37430, n37431, n37432, n37433, n37434, n37435, n37436,
         n37437, n37438, n37439, n37440, n37441, n37442, n37443, n37444,
         n37445, n37446, n37447, n37448, n37449, n37450, n37451, n37452,
         n37453, n37454, n37455, n37456, n37457, n37458, n37459, n37460,
         n37461, n37462, n37463, n37464, n37465, n37466, n37467, n37468,
         n37469, n37470, n37471, n37472, n37473, n37474, n37475, n37476,
         n37477, n37478, n37479, n37480, n37481, n37482, n37483, n37484,
         n37485, n37486, n37487, n37488, n37489, n37490, n37491, n37492,
         n37493, n37494, n37495, n37496, n37497, n37498, n37499, n37500,
         n37501, n37502, n37503, n37504, n37505, n37506, n37507, n37508,
         n37509, n37510, n37511, n37512, n37513, n37514, n37515, n37516,
         n37517, n37518, n37519, n37520, n37521, n37522, n37523, n37524,
         n37525, n37526, n37527, n37528, n37529, n37530, n37531, n37532,
         n37533, n37534, n37535, n37536, n37537, n37538, n37539, n37540,
         n37541, n37542, n37543, n37544, n37545, n37546, n37547, n37548,
         n37549, n37550, n37551, n37552, n37553, n37554, n37555, n37556,
         n37557, n37558, n37559, n37560, n37561, n37562, n37563, n37564,
         n37565, n37566, n37567, n37568, n37569, n37570, n37571, n37572,
         n37573, n37574, n37575, n37576, n37577, n37578, n37579, n37580,
         n37581, n37582, n37583, n37584, n37585, n37586, n37587, n37588,
         n37589, n37590, n37591, n37592, n37593, n37594, n37595, n37596,
         n37597, n37598, n37599, n37600, n37601, n37602, n37603, n37604,
         n37605, n37606, n37607, n37608, n37609, n37610, n37611, n37612,
         n37613, n37614, n37615, n37616, n37617, n37618, n37619, n37620,
         n37621, n37622, n37623, n37624, n37625, n37626, n37627, n37628,
         n37629, n37630, n37631, n37632, n37633, n37634, n37635, n37636,
         n37637, n37638, n37639, n37640, n37641, n37642, n37643, n37644,
         n37645, n37646, n37647, n37648, n37649, n37650, n37651, n37652,
         n37653, n37654, n37655, n37656, n37657, n37658, n37659, n37660,
         n37661, n37662, n37663, n37664, n37665, n37666, n37667, n37668,
         n37669, n37670, n37671, n37672, n37673, n37674, n37675, n37676,
         n37677, n37678, n37679, n37680, n37681, n37682, n37683, n37684,
         n37685, n37686, n37687, n37688, n37689, n37690, n37691, n37692,
         n37693, n37694, n37695, n37696, n37697, n37698, n37699, n37700,
         n37701, n37702, n37703, n37704, n37705, n37706, n37707, n37708,
         n37709, n37710, n37711, n37712, n37713, n37714, n37715, n37716,
         n37717, n37718, n37719, n37720, n37721, n37722, n37723, n37724,
         n37725, n37726, n37727, n37728, n37729, n37730, n37731, n37732,
         n37733, n37734, n37735, n37736, n37737, n37738, n37739, n37740,
         n37741, n37742, n37743, n37744, n37745, n37746, n37747, n37748,
         n37749, n37750, n37751, n37752, n37753, n37754, n37755, n37756,
         n37757, n37758, n37759, n37760, n37761, n37762, n37763, n37764,
         n37765, n37766, n37767, n37768, n37769, n37770, n37771, n37772,
         n37773, n37774, n37775, n37776, n37777, n37778, n37779, n37780,
         n37781, n37782, n37783, n37784, n37785, n37786, n37787, n37788,
         n37789, n37790, n37791, n37792, n37793, n37794, n37795, n37796,
         n37797, n37798, n37799, n37800, n37801, n37802, n37803, n37804,
         n37805, n37806, n37807, n37808, n37809, n37810, n37811, n37812,
         n37813, n37814, n37815, n37816, n37817, n37818, n37819, n37820,
         n37821, n37822, n37823, n37824, n37825, n37826, n37827, n37828,
         n37829, n37830, n37831, n37832, n37833, n37834, n37835, n37836,
         n37837, n37838, n37839, n37840, n37841, n37842, n37843, n37844,
         n37845, n37846, n37847, n37848, n37849, n37850, n37851, n37852,
         n37853, n37854, n37855, n37856, n37857, n37858, n37859, n37860,
         n37861, n37862, n37863, n37864, n37865, n37866, n37867, n37868,
         n37869, n37870, n37871, n37872, n37873, n37874, n37875, n37876,
         n37877, n37878, n37879, n37880, n37881, n37882, n37883, n37884,
         n37885, n37886, n37887, n37888, n37889, n37890, n37891, n37892,
         n37893, n37894, n37895, n37896, n37897, n37898, n37899, n37900,
         n37901, n37902, n37903, n37904, n37905, n37906, n37907, n37908,
         n37909, n37910, n37911, n37912, n37913, n37914, n37915, n37916,
         n37917, n37918, n37919, n37920, n37921, n37922, n37923, n37924,
         n37925, n37926, n37927, n37928, n37929, n37930, n37931, n37932,
         n37933, n37934, n37935, n37936, n37937, n37938, n37939, n37940,
         n37941, n37942, n37943, n37944, n37945, n37946, n37947, n37948,
         n37949, n37950, n37951, n37952, n37953, n37954, n37955, n37956,
         n37957, n37958, n37959, n37960, n37961, n37962, n37963, n37964,
         n37965, n37966, n37967, n37968, n37969, n37970, n37971, n37972,
         n37973, n37974, n37975, n37976, n37977, n37978, n37979, n37980,
         n37981, n37982, n37983, n37984, n37985, n37986, n37987, n37988,
         n37989, n37990, n37991, n37992, n37993, n37994, n37995, n37996,
         n37997, n37998, n37999, n38000, n38001, n38002, n38003, n38004,
         n38005, n38006, n38007, n38008, n38009, n38010, n38011, n38012,
         n38013, n38014, n38015, n38016, n38017, n38018, n38019, n38020,
         n38021, n38022, n38023, n38024, n38025, n38026, n38027, n38028,
         n38029, n38030, n38031, n38032, n38033, n38034, n38035, n38036,
         n38037, n38038, n38039, n38040, n38041, n38042, n38043, n38044,
         n38045, n38046, n38047, n38048, n38049, n38050, n38051, n38052,
         n38053, n38054, n38055, n38056, n38057, n38058, n38059, n38060,
         n38061, n38062, n38063, n38064, n38065, n38066, n38067, n38068,
         n38069, n38070, n38071, n38072, n38073, n38074, n38075, n38076,
         n38077, n38078, n38079, n38080, n38081, n38082, n38083, n38084,
         n38085, n38086, n38087, n38088, n38089, n38090, n38091, n38092,
         n38093, n38094, n38095, n38096, n38097, n38098, n38099, n38100,
         n38101, n38102, n38103, n38104, n38105, n38106, n38107, n38108,
         n38109, n38110, n38111, n38112, n38113, n38114, n38115, n38116,
         n38117, n38118, n38119, n38120, n38121, n38122, n38123, n38124,
         n38125, n38126, n38127, n38128, n38129, n38130, n38131, n38132,
         n38133, n38134, n38135, n38136, n38137, n38138, n38139, n38140,
         n38141, n38142, n38143, n38144, n38145, n38146, n38147, n38148,
         n38149, n38150, n38151, n38152, n38153, n38154, n38155, n38156,
         n38157, n38158, n38159, n38160, n38161, n38162, n38163, n38164,
         n38165, n38166, n38167, n38168, n38169, n38170, n38171, n38172,
         n38173, n38174, n38175, n38176, n38177, n38178, n38179, n38180,
         n38181, n38182, n38183, n38184, n38185, n38186, n38187, n38188,
         n38189, n38190, n38191, n38192, n38193, n38194, n38195, n38196,
         n38197, n38198, n38199, n38200, n38201, n38202, n38203, n38204,
         n38205, n38206, n38207, n38208, n38209, n38210, n38211, n38212,
         n38213, n38214, n38215, n38216, n38217, n38218, n38219, n38220,
         n38221, n38222, n38223, n38224, n38225, n38226, n38227, n38228,
         n38229, n38230, n38231, n38232, n38233, n38234, n38235, n38236,
         n38237, n38238, n38239, n38240, n38241, n38242, n38243, n38244,
         n38245, n38246, n38247, n38248, n38249, n38250, n38251, n38252,
         n38253, n38254, n38255, n38256, n38257, n38258, n38259, n38260,
         n38261, n38262, n38263, n38264, n38265, n38266, n38267, n38268,
         n38269, n38270, n38271, n38272, n38273, n38274, n38275, n38276,
         n38277, n38278, n38279, n38280, n38281, n38282, n38283, n38284,
         n38285, n38286, n38287, n38288, n38289, n38290, n38291, n38292,
         n38293, n38294, n38295, n38296, n38297, n38298, n38299, n38300,
         n38301, n38302, n38303, n38304, n38305, n38306, n38307, n38308,
         n38309, n38310, n38311, n38312, n38313, n38314, n38315, n38316,
         n38317, n38318, n38319, n38320, n38321, n38322, n38323, n38324,
         n38325, n38326, n38327, n38328, n38329, n38330, n38331, n38332,
         n38333, n38334, n38335, n38336, n38337, n38338, n38339, n38340,
         n38341, n38342, n38343, n38344, n38345, n38346, n38347, n38348,
         n38349, n38350, n38351, n38352, n38353, n38354, n38355, n38356,
         n38357, n38358, n38359, n38360, n38361, n38362, n38363, n38364,
         n38365, n38366, n38367, n38368, n38369, n38370, n38371, n38372,
         n38373, n38374, n38375, n38376, n38377, n38378, n38379, n38380,
         n38381, n38382, n38383, n38384, n38385, n38386, n38387, n38388,
         n38389, n38390, n38391, n38392, n38393, n38394, n38395, n38396,
         n38397, n38398, n38399, n38400, n38401, n38402, n38403, n38404,
         n38405, n38406, n38407, n38408, n38409, n38410, n38411, n38412,
         n38413, n38414, n38415, n38416, n38417, n38418, n38419, n38420,
         n38421, n38422, n38423, n38424, n38425, n38426, n38427, n38428,
         n38429, n38430, n38431, n38432, n38433, n38434, n38435, n38436,
         n38437, n38438, n38439, n38440, n38441, n38442, n38443, n38444,
         n38445, n38446, n38447, n38448, n38449, n38450, n38451, n38452,
         n38453, n38454, n38455, n38456, n38457, n38458, n38459, n38460,
         n38461, n38462, n38463, n38464, n38465, n38466, n38467, n38468,
         n38469, n38470, n38471, n38472, n38473, n38474, n38475, n38476,
         n38477, n38478, n38479, n38480, n38481, n38482, n38483, n38484,
         n38485, n38486, n38487, n38488, n38489, n38490, n38491, n38492,
         n38493, n38494, n38495, n38496, n38497, n38498, n38499, n38500,
         n38501, n38502, n38503, n38504, n38505, n38506, n38507, n38508,
         n38509, n38510, n38511, n38512, n38513, n38514, n38515, n38516,
         n38517, n38518, n38519, n38520, n38521, n38522, n38523, n38524,
         n38525, n38526, n38527, n38528, n38529, n38530, n38531, n38532,
         n38533, n38534, n38535, n38536, n38537, n38538, n38539, n38540,
         n38541, n38542, n38543, n38544, n38545, n38546, n38547, n38548,
         n38549, n38550, n38551, n38552, n38553, n38554, n38555, n38556,
         n38557, n38558, n38559, n38560, n38561, n38562, n38563, n38564,
         n38565, n38566, n38567, n38568, n38569, n38570, n38571, n38572,
         n38573, n38574, n38575, n38576, n38577, n38578, n38579, n38580,
         n38581, n38582, n38583, n38584, n38585, n38586, n38587, n38588,
         n38589, n38590, n38591, n38592, n38593, n38594, n38595, n38596,
         n38597, n38598, n38599, n38600, n38601, n38602, n38603, n38604,
         n38605, n38606, n38607, n38608, n38609, n38610, n38611, n38612,
         n38613, n38614, n38615, n38616, n38617, n38618, n38619, n38620,
         n38621, n38622, n38623, n38624, n38625, n38626, n38627, n38628,
         n38629, n38630, n38631, n38632, n38633, n38634, n38635, n38636,
         n38637, n38638, n38639, n38640, n38641, n38642, n38643, n38644,
         n38645, n38646, n38647, n38648, n38649, n38650, n38651, n38652,
         n38653, n38654, n38655, n38656, n38657, n38658, n38659, n38660,
         n38661, n38662, n38663, n38664, n38665, n38666, n38667, n38668,
         n38669, n38670, n38671, n38672, n38673, n38674, n38675, n38676,
         n38677, n38678, n38679, n38680, n38681, n38682, n38683, n38684,
         n38685, n38686, n38687, n38688, n38689, n38690, n38691, n38692,
         n38693, n38694, n38695, n38696, n38697, n38698, n38699, n38700,
         n38701, n38702, n38703, n38704, n38705, n38706, n38707, n38708,
         n38709, n38710, n38711, n38712, n38713, n38714, n38715, n38716,
         n38717, n38718, n38719, n38720, n38721, n38722, n38723, n38724,
         n38725, n38726, n38727, n38728, n38729, n38730, n38731, n38732,
         n38733, n38734, n38735, n38736, n38737, n38738, n38739, n38740,
         n38741, n38742, n38743, n38744, n38745, n38746, n38747, n38748,
         n38749, n38750, n38751, n38752, n38753, n38754, n38755, n38756,
         n38757, n38758, n38759, n38760, n38761, n38762, n38763, n38764,
         n38765, n38766, n38767, n38768, n38769, n38770, n38771, n38772,
         n38773, n38774, n38775, n38776, n38777, n38778, n38779, n38780,
         n38781, n38782, n38783, n38784, n38785, n38786, n38787, n38788,
         n38789, n38790, n38791, n38792, n38793, n38794, n38795, n38796,
         n38797, n38798, n38799, n38800, n38801, n38802, n38803, n38804,
         n38805, n38806, n38807, n38808, n38809, n38810, n38811, n38812,
         n38813, n38814, n38815, n38816, n38817, n38818, n38819, n38820,
         n38821, n38822, n38823, n38824, n38825, n38826, n38827, n38828,
         n38829, n38830, n38831, n38832, n38833, n38834, n38835, n38836,
         n38837, n38838, n38839, n38840, n38841, n38842, n38843, n38844,
         n38845, n38846, n38847, n38848, n38849, n38850, n38851, n38852,
         n38853, n38854, n38855, n38856, n38857, n38858, n38859, n38860,
         n38861, n38862, n38863, n38864, n38865, n38866, n38867, n38868,
         n38869, n38870, n38871, n38872, n38873, n38874, n38875, n38876,
         n38877, n38878, n38879, n38880, n38881, n38882, n38883, n38884,
         n38885, n38886, n38887, n38888, n38889, n38890, n38891, n38892,
         n38893, n38894, n38895, n38896, n38897, n38898, n38899, n38900,
         n38901, n38902, n38903, n38904, n38905, n38906, n38907, n38908,
         n38909, n38910, n38911, n38912, n38913, n38914, n38915, n38916,
         n38917, n38918, n38919, n38920, n38921, n38922, n38923, n38924,
         n38925, n38926, n38927, n38928, n38929, n38930, n38931, n38932,
         n38933, n38934, n38935, n38936, n38937, n38938, n38939, n38940,
         n38941, n38942, n38943, n38944, n38945, n38946, n38947, n38948,
         n38949, n38950, n38951, n38952, n38953, n38954, n38955, n38956,
         n38957, n38958, n38959, n38960, n38961, n38962, n38963, n38964,
         n38965, n38966, n38967, n38968, n38969, n38970, n38971, n38972,
         n38973, n38974, n38975, n38976, n38977, n38978, n38979, n38980,
         n38981, n38982, n38983, n38984, n38985, n38986, n38987, n38988,
         n38989, n38990, n38991, n38992, n38993, n38994, n38995, n38996,
         n38997, n38998, n38999, n39000, n39001, n39002, n39003, n39004,
         n39005, n39006, n39007, n39008, n39009, n39010, n39011, n39012,
         n39013, n39014, n39015, n39016, n39017, n39018, n39019, n39020,
         n39021, n39022, n39023, n39024, n39025, n39026, n39027, n39028,
         n39029, n39030, n39031, n39032, n39033, n39034, n39035, n39036,
         n39037, n39038, n39039, n39040, n39041, n39042, n39043, n39044,
         n39045, n39046, n39047, n39048, n39049, n39050, n39051, n39052,
         n39053, n39054, n39055, n39056, n39057, n39058, n39059, n39060,
         n39061, n39062, n39063, n39064, n39065, n39066, n39067, n39068,
         n39069, n39070, n39071, n39072, n39073, n39074, n39075, n39076,
         n39077, n39078, n39079, n39080, n39081, n39082, n39083, n39084,
         n39085, n39086, n39087, n39088, n39089, n39090, n39091, n39092,
         n39093, n39094, n39095, n39096, n39097, n39098, n39099, n39100,
         n39101, n39102, n39103, n39104, n39105, n39106, n39107, n39108,
         n39109, n39110, n39111, n39112, n39113, n39114, n39115, n39116,
         n39117, n39118, n39119, n39120, n39121, n39122, n39123, n39124,
         n39125, n39126, n39127, n39128, n39129, n39130, n39131, n39132,
         n39133, n39134, n39135, n39136, n39137, n39138, n39139, n39140,
         n39141, n39142, n39143, n39144, n39145, n39146, n39147, n39148,
         n39149, n39150, n39151, n39152, n39153, n39154, n39155, n39156,
         n39157, n39158, n39159, n39160, n39161, n39162, n39163, n39164,
         n39165, n39166, n39167, n39168, n39169, n39170, n39171, n39172,
         n39173, n39174, n39175, n39176, n39177, n39178, n39179, n39180,
         n39181, n39182, n39183, n39184, n39185, n39186, n39187, n39188,
         n39189, n39190, n39191, n39192, n39193, n39194, n39195, n39196,
         n39197, n39198, n39199, n39200, n39201, n39202, n39203, n39204,
         n39205, n39206, n39207, n39208, n39209, n39210, n39211, n39212,
         n39213, n39214, n39215, n39216, n39217, n39218, n39219, n39220,
         n39221, n39222, n39223, n39224, n39225, n39226, n39227, n39228,
         n39229, n39230, n39231, n39232, n39233, n39234, n39235, n39236,
         n39237, n39238, n39239, n39240, n39241, n39242, n39243, n39244,
         n39245, n39246, n39247, n39248, n39249, n39250, n39251, n39252,
         n39253, n39254, n39255, n39256, n39257, n39258, n39259, n39260,
         n39261, n39262, n39263, n39264, n39265, n39266, n39267, n39268,
         n39269, n39270, n39271, n39272, n39273, n39274, n39275, n39276,
         n39277, n39278, n39279, n39280, n39281, n39282, n39283, n39284,
         n39285, n39286, n39287, n39288, n39289, n39290, n39291, n39292,
         n39293, n39294, n39295, n39296, n39297, n39298, n39299, n39300,
         n39301, n39302, n39303, n39304, n39305, n39306, n39307, n39308,
         n39309, n39310, n39311, n39312, n39313, n39314, n39315, n39316,
         n39317, n39318, n39319, n39320, n39321, n39322, n39323, n39324,
         n39325, n39326, n39327, n39328, n39329, n39330, n39331, n39332,
         n39333, n39334, n39335, n39336, n39337, n39338, n39339, n39340,
         n39341, n39342, n39343, n39344, n39345, n39346, n39347, n39348,
         n39349, n39350, n39351, n39352, n39353, n39354, n39355, n39356,
         n39357, n39358, n39359, n39360, n39361, n39362, n39363, n39364,
         n39365, n39366, n39367, n39368, n39369, n39370, n39371, n39372,
         n39373, n39374, n39375, n39376, n39377, n39378, n39379, n39380,
         n39381, n39382, n39383, n39384, n39385, n39386, n39387, n39388,
         n39389, n39390, n39391, n39392, n39393, n39394, n39395, n39396,
         n39397, n39398, n39399, n39400, n39401, n39402, n39403, n39404,
         n39405, n39406, n39407, n39408, n39409, n39410, n39411, n39412,
         n39413, n39414, n39415, n39416, n39417, n39418, n39419, n39420,
         n39421, n39422, n39423, n39424, n39425, n39426, n39427, n39428,
         n39429, n39430, n39431, n39432, n39433, n39434, n39435, n39436,
         n39437, n39438, n39439, n39440, n39441, n39442, n39443, n39444,
         n39445, n39446, n39447, n39448, n39449, n39450, n39451, n39452,
         n39453, n39454, n39455, n39456, n39457, n39458, n39459, n39460,
         n39461, n39462, n39463, n39464, n39465, n39466, n39467, n39468,
         n39469, n39470, n39471, n39472, n39473, n39474, n39475, n39476,
         n39477, n39478, n39479, n39480, n39481, n39482, n39483, n39484,
         n39485, n39486, n39487, n39488, n39489, n39490, n39491, n39492,
         n39493, n39494, n39495, n39496, n39497, n39498, n39499, n39500,
         n39501, n39502, n39503, n39504, n39505, n39506, n39507, n39508,
         n39509, n39510, n39511, n39512, n39513, n39514, n39515, n39516,
         n39517, n39518, n39519, n39520, n39521, n39522, n39523, n39524,
         n39525, n39526, n39527, n39528, n39529, n39530, n39531, n39532,
         n39533, n39534, n39535, n39536, n39537, n39538, n39539, n39540,
         n39541, n39542, n39543, n39544, n39545, n39546, n39547, n39548,
         n39549, n39550, n39551, n39552, n39553, n39554, n39555, n39556,
         n39557, n39558, n39559, n39560, n39561, n39562, n39563, n39564,
         n39565, n39566, n39567, n39568, n39569, n39570, n39571, n39572,
         n39573, n39574, n39575, n39576, n39577, n39578, n39579, n39580,
         n39581, n39582, n39583, n39584, n39585, n39586, n39587, n39588,
         n39589, n39590, n39591, n39592, n39593, n39594, n39595, n39596,
         n39597, n39598, n39599, n39600, n39601, n39602, n39603, n39604,
         n39605, n39606, n39607, n39608, n39609, n39610, n39611, n39612,
         n39613, n39614, n39615, n39616, n39617, n39618, n39619, n39620,
         n39621, n39622, n39623, n39624, n39625, n39626, n39627, n39628,
         n39629, n39630, n39631, n39632, n39633, n39634, n39635, n39636,
         n39637, n39638, n39639, n39640, n39641, n39642, n39643, n39644,
         n39645, n39646, n39647, n39648, n39649, n39650, n39651, n39652,
         n39653, n39654, n39655, n39656, n39657, n39658, n39659, n39660,
         n39661, n39662, n39663, n39664, n39665, n39666, n39667, n39668,
         n39669, n39670, n39671, n39672, n39673, n39674, n39675, n39676,
         n39677, n39678, n39679, n39680, n39681, n39682, n39683, n39684,
         n39685, n39686, n39687, n39688, n39689, n39690, n39691, n39692,
         n39693, n39694, n39695, n39696, n39697, n39698, n39699, n39700,
         n39701, n39702, n39703, n39704, n39705, n39706, n39707, n39708,
         n39709, n39710, n39711, n39712, n39713, n39714, n39715, n39716,
         n39717, n39718, n39719, n39720, n39721, n39722, n39723, n39724,
         n39725, n39726, n39727, n39728, n39729, n39730, n39731, n39732,
         n39733, n39734, n39735, n39736, n39737, n39738, n39739, n39740,
         n39741, n39742, n39743, n39744, n39745, n39746, n39747, n39748,
         n39749, n39750, n39751, n39752, n39753, n39754, n39755, n39756,
         n39757, n39758, n39759, n39760, n39761, n39762, n39763, n39764,
         n39765, n39766, n39767, n39768, n39769, n39770, n39771, n39772,
         n39773, n39774, n39775, n39776, n39777, n39778, n39779, n39780,
         n39781, n39782, n39783, n39784, n39785, n39786, n39787, n39788,
         n39789, n39790, n39791, n39792, n39793, n39794, n39795, n39796,
         n39797, n39798, n39799, n39800, n39801, n39802, n39803, n39804,
         n39805, n39806, n39807, n39808, n39809, n39810, n39811, n39812,
         n39813, n39814, n39815, n39816, n39817, n39818, n39819, n39820,
         n39821, n39822, n39823, n39824, n39825, n39826, n39827, n39828,
         n39829, n39830, n39831, n39832, n39833, n39834, n39835, n39836,
         n39837, n39838, n39839, n39840, n39841, n39842, n39843, n39844,
         n39845, n39846, n39847, n39848, n39849, n39850, n39851, n39852,
         n39853, n39854, n39855, n39856, n39857, n39858, n39859, n39860,
         n39861, n39862, n39863, n39864, n39865, n39866, n39867, n39868,
         n39869, n39870, n39871, n39872, n39873, n39874, n39875, n39876,
         n39877, n39878, n39879, n39880, n39881, n39882, n39883, n39884,
         n39885, n39886, n39887, n39888, n39889, n39890, n39891, n39892,
         n39893, n39894, n39895, n39896, n39897, n39898, n39899, n39900,
         n39901, n39902, n39903, n39904, n39905, n39906, n39907, n39908,
         n39909, n39910, n39911, n39912, n39913, n39914, n39915, n39916,
         n39917, n39918, n39919, n39920, n39921, n39922, n39923, n39924,
         n39925, n39926, n39927, n39928, n39929, n39930, n39931, n39932,
         n39933, n39934, n39935, n39936, n39937, n39938, n39939, n39940,
         n39941, n39942, n39943, n39944, n39945, n39946, n39947, n39948,
         n39949, n39950, n39951, n39952, n39953, n39954, n39955, n39956,
         n39957, n39958, n39959, n39960, n39961, n39962, n39963, n39964,
         n39965, n39966, n39967, n39968, n39969, n39970, n39971, n39972,
         n39973, n39974, n39975, n39976, n39977, n39978, n39979, n39980,
         n39981, n39982, n39983, n39984, n39985, n39986, n39987, n39988,
         n39989, n39990, n39991, n39992, n39993, n39994, n39995, n39996,
         n39997, n39998, n39999, n40000, n40001, n40002, n40003, n40004,
         n40005, n40006, n40007, n40008, n40009, n40010, n40011, n40012,
         n40013, n40014, n40015, n40016, n40017, n40018, n40019, n40020,
         n40021, n40022, n40023, n40024, n40025, n40026, n40027, n40028,
         n40029, n40030, n40031, n40032, n40033, n40034, n40035, n40036,
         n40037, n40038, n40039, n40040, n40041, n40042, n40043, n40044,
         n40045, n40046, n40047, n40048, n40049, n40050, n40051, n40052,
         n40053, n40054, n40055, n40056, n40057, n40058, n40059, n40060,
         n40061, n40062, n40063, n40064, n40065, n40066, n40067, n40068,
         n40069, n40070, n40071, n40072, n40073, n40074, n40075, n40076,
         n40077, n40078, n40079, n40080, n40081, n40082, n40083, n40084,
         n40085, n40086, n40087, n40088, n40089, n40090, n40091, n40092,
         n40093, n40094, n40095, n40096, n40097, n40098, n40099, n40100,
         n40101, n40102, n40103, n40104, n40105, n40106, n40107, n40108,
         n40109, n40110, n40111, n40112, n40113, n40114, n40115, n40116,
         n40117, n40118, n40119, n40120, n40121, n40122, n40123, n40124,
         n40125, n40126, n40127, n40128, n40129, n40130, n40131, n40132,
         n40133, n40134, n40135, n40136, n40137, n40138, n40139, n40140,
         n40141, n40142, n40143, n40144, n40145, n40146, n40147, n40148,
         n40149, n40150, n40151, n40152, n40153, n40154, n40155, n40156,
         n40157, n40158, n40159, n40160, n40161, n40162, n40163, n40164,
         n40165, n40166, n40167, n40168, n40169, n40170, n40171, n40172,
         n40173, n40174, n40175, n40176, n40177, n40178, n40179, n40180,
         n40181, n40182, n40183, n40184, n40185, n40186, n40187, n40188,
         n40189, n40190, n40191, n40192, n40193, n40194, n40195, n40196,
         n40197, n40198, n40199, n40200, n40201, n40202, n40203, n40204,
         n40205, n40206, n40207, n40208, n40209, n40210, n40211, n40212,
         n40213, n40214, n40215, n40216, n40217, n40218, n40219, n40220,
         n40221, n40222, n40223, n40224, n40225, n40226, n40227, n40228,
         n40229, n40230, n40231, n40232, n40233, n40234, n40235, n40236,
         n40237, n40238, n40239, n40240, n40241, n40242, n40243, n40244,
         n40245, n40246, n40247, n40248, n40249, n40250, n40251, n40252,
         n40253, n40254, n40255, n40256, n40257, n40258, n40259, n40260,
         n40261, n40262, n40263, n40264, n40265, n40266, n40267, n40268,
         n40269, n40270, n40271, n40272, n40273, n40274, n40275, n40276,
         n40277, n40278, n40279, n40280, n40281, n40282, n40283, n40284,
         n40285, n40286, n40287, n40288, n40289, n40290, n40291, n40292,
         n40293, n40294, n40295, n40296, n40297, n40298, n40299, n40300,
         n40301, n40302, n40303, n40304, n40305, n40306, n40307, n40308,
         n40309, n40310, n40311, n40312, n40313, n40314, n40315, n40316,
         n40317, n40318, n40319, n40320, n40321, n40322, n40323, n40324,
         n40325, n40326, n40327, n40328, n40329, n40330, n40331, n40332,
         n40333, n40334, n40335, n40336, n40337, n40338, n40339, n40340,
         n40341, n40342, n40343, n40344, n40345, n40346, n40347, n40348,
         n40349, n40350, n40351, n40352, n40353, n40354, n40355, n40356,
         n40357, n40358, n40359, n40360, n40361, n40362, n40363, n40364,
         n40365, n40366, n40367, n40368, n40369, n40370, n40371, n40372,
         n40373, n40374, n40375, n40376, n40377, n40378, n40379, n40380,
         n40381, n40382, n40383, n40384, n40385, n40386, n40387, n40388,
         n40389, n40390, n40391, n40392, n40393, n40394, n40395, n40396,
         n40397, n40398, n40399, n40400, n40401, n40402, n40403, n40404,
         n40405, n40406, n40407, n40408, n40409, n40410, n40411, n40412,
         n40413, n40414, n40415, n40416, n40417, n40418, n40419, n40420,
         n40421, n40422, n40423, n40424, n40425, n40426, n40427, n40428,
         n40429, n40430, n40431, n40432, n40433, n40434, n40435, n40436,
         n40437, n40438, n40439, n40440, n40441, n40442, n40443, n40444,
         n40445, n40446, n40447, n40448, n40449, n40450, n40451, n40452,
         n40453, n40454, n40455, n40456, n40457, n40458, n40459, n40460,
         n40461, n40462, n40463, n40464, n40465, n40466, n40467, n40468,
         n40469, n40470, n40471, n40472, n40473, n40474, n40475, n40476,
         n40477, n40478, n40479, n40480, n40481, n40482, n40483, n40484,
         n40485, n40486, n40487, n40488, n40489, n40490, n40491, n40492,
         n40493, n40494, n40495, n40496, n40497, n40498, n40499, n40500,
         n40501, n40502, n40503, n40504, n40505, n40506, n40507, n40508,
         n40509, n40510, n40511, n40512, n40513, n40514, n40515, n40516,
         n40517, n40518, n40519, n40520, n40521, n40522, n40523, n40524,
         n40525, n40526, n40527, n40528, n40529, n40530, n40531, n40532,
         n40533, n40534, n40535, n40536, n40537, n40538, n40539, n40540,
         n40541, n40542, n40543, n40544, n40545, n40546, n40547, n40548,
         n40549, n40550, n40551, n40552, n40553, n40554, n40555, n40556,
         n40557, n40558, n40559, n40560, n40561, n40562, n40563, n40564,
         n40565, n40566, n40567, n40568, n40569, n40570, n40571, n40572,
         n40573, n40574, n40575, n40576, n40577, n40578, n40579, n40580,
         n40581, n40582, n40583, n40584, n40585, n40586, n40587, n40588,
         n40589, n40590, n40591, n40592, n40593, n40594, n40595, n40596,
         n40597, n40598, n40599, n40600, n40601, n40602, n40603, n40604,
         n40605, n40606, n40607, n40608, n40609, n40610, n40611, n40612,
         n40613, n40614, n40615, n40616, n40617, n40618, n40619, n40620,
         n40621, n40622, n40623, n40624, n40625, n40626, n40627, n40628,
         n40629, n40630, n40631, n40632, n40633, n40634, n40635, n40636,
         n40637, n40638, n40639, n40640, n40641, n40642, n40643, n40644,
         n40645, n40646, n40647, n40648, n40649, n40650, n40651, n40652,
         n40653, n40654, n40655, n40656, n40657, n40658, n40659, n40660,
         n40661, n40662, n40663, n40664, n40665, n40666, n40667, n40668,
         n40669, n40670, n40671, n40672, n40673, n40674, n40675, n40676,
         n40677, n40678, n40679, n40680, n40681, n40682, n40683, n40684,
         n40685, n40686, n40687, n40688, n40689, n40690, n40691, n40692,
         n40693, n40694, n40695, n40696, n40697, n40698, n40699, n40700,
         n40701, n40702, n40703, n40704, n40705, n40706, n40707, n40708,
         n40709, n40710, n40711, n40712, n40713, n40714, n40715, n40716,
         n40717, n40718, n40719, n40720, n40721, n40722, n40723, n40724,
         n40725, n40726, n40727, n40728, n40729, n40730, n40731, n40732,
         n40733, n40734, n40735, n40736, n40737, n40738, n40739, n40740,
         n40741, n40742, n40743, n40744, n40745, n40746, n40747, n40748,
         n40749, n40750, n40751, n40752, n40753, n40754, n40755, n40756,
         n40757, n40758, n40759, n40760, n40761, n40762, n40763, n40764,
         n40765, n40766, n40767, n40768, n40769, n40770, n40771, n40772,
         n40773, n40774, n40775, n40776, n40777, n40778, n40779, n40780,
         n40781, n40782, n40783, n40784, n40785, n40786, n40787, n40788,
         n40789, n40790, n40791, n40792, n40793, n40794, n40795, n40796,
         n40797, n40798, n40799, n40800, n40801, n40802, n40803, n40804,
         n40805, n40806, n40807, n40808, n40809, n40810, n40811, n40812,
         n40813, n40814, n40815, n40816, n40817, n40818, n40819, n40820,
         n40821, n40822, n40823, n40824, n40825, n40826, n40827, n40828,
         n40829, n40830, n40831, n40832, n40833, n40834, n40835, n40836,
         n40837, n40838, n40839, n40840, n40841, n40842, n40843, n40844,
         n40845, n40846, n40847, n40848, n40849, n40850, n40851, n40852,
         n40853, n40854, n40855, n40856, n40857, n40858, n40859, n40860,
         n40861, n40862, n40863, n40864, n40865, n40866, n40867, n40868,
         n40869, n40870, n40871, n40872, n40873, n40874, n40875, n40876,
         n40877, n40878, n40879, n40880, n40881, n40882, n40883, n40884,
         n40885, n40886, n40887, n40888, n40889, n40890, n40891, n40892,
         n40893, n40894, n40895, n40896, n40897, n40898, n40899, n40900,
         n40901, n40902, n40903, n40904, n40905, n40906, n40907, n40908,
         n40909, n40910, n40911, n40912, n40913, n40914, n40915, n40916,
         n40917, n40918, n40919, n40920, n40921, n40922, n40923, n40924,
         n40925, n40926, n40927, n40928, n40929, n40930, n40931, n40932,
         n40933, n40934, n40935, n40936, n40937, n40938, n40939, n40940,
         n40941, n40942, n40943, n40944, n40945, n40946, n40947, n40948,
         n40949, n40950, n40951, n40952, n40953, n40954, n40955, n40956,
         n40957, n40958, n40959, n40960, n40961, n40962, n40963, n40964,
         n40965, n40966, n40967, n40968, n40969, n40970, n40971, n40972,
         n40973, n40974, n40975, n40976, n40977, n40978, n40979, n40980,
         n40981, n40982, n40983, n40984, n40985, n40986, n40987, n40988,
         n40989, n40990, n40991, n40992, n40993, n40994, n40995, n40996,
         n40997, n40998, n40999, n41000, n41001, n41002, n41003, n41004,
         n41005, n41006, n41007, n41008, n41009, n41010, n41011, n41012,
         n41013, n41014, n41015, n41016, n41017, n41018, n41019, n41020,
         n41021, n41022, n41023, n41024, n41025, n41026, n41027, n41028,
         n41029, n41030, n41031, n41032, n41033, n41034, n41035, n41036,
         n41037, n41038, n41039, n41040, n41041, n41042, n41043, n41044,
         n41045, n41046, n41047, n41048, n41049, n41050, n41051, n41052,
         n41053, n41054, n41055, n41056, n41057, n41058, n41059, n41060,
         n41061, n41062, n41063, n41064, n41065, n41066, n41067, n41068,
         n41069, n41070, n41071, n41072, n41073, n41074, n41075, n41076,
         n41077, n41078, n41079, n41080, n41081, n41082, n41083, n41084,
         n41085, n41086, n41087, n41088, n41089, n41090, n41091, n41092,
         n41093, n41094, n41095, n41096, n41097, n41098, n41099, n41100,
         n41101, n41102, n41103, n41104, n41105, n41106, n41107, n41108,
         n41109, n41110, n41111, n41112, n41113, n41114, n41115, n41116,
         n41117, n41118, n41119, n41120, n41121, n41122, n41123, n41124,
         n41125, n41126, n41127, n41128, n41129, n41130, n41131, n41132,
         n41133, n41134, n41135, n41136, n41137, n41138, n41139, n41140,
         n41141, n41142, n41143, n41144, n41145, n41146, n41147, n41148,
         n41149, n41150, n41151, n41152, n41153, n41154, n41155, n41156,
         n41157, n41158, n41159, n41160, n41161, n41162, n41163, n41164,
         n41165, n41166, n41167, n41168, n41169, n41170, n41171, n41172,
         n41173, n41174, n41175, n41176, n41177, n41178, n41179, n41180,
         n41181, n41182, n41183, n41184, n41185, n41186, n41187, n41188,
         n41189, n41190, n41191, n41192, n41193, n41194, n41195, n41196,
         n41197, n41198, n41199, n41200, n41201, n41202, n41203, n41204,
         n41205, n41206, n41207, n41208, n41209, n41210, n41211, n41212,
         n41213, n41214, n41215, n41216, n41217, n41218, n41219, n41220,
         n41221, n41222, n41223, n41224, n41225, n41226, n41227, n41228,
         n41229, n41230, n41231, n41232, n41233, n41234, n41235, n41236,
         n41237, n41238, n41239, n41240, n41241, n41242, n41243, n41244,
         n41245, n41246, n41247, n41248, n41249, n41250, n41251, n41252,
         n41253, n41254, n41255, n41256, n41257, n41258, n41259, n41260,
         n41261, n41262, n41263, n41264, n41265, n41266, n41267, n41268,
         n41269, n41270, n41271, n41272, n41273, n41274, n41275, n41276,
         n41277, n41278, n41279, n41280, n41281, n41282, n41283, n41284,
         n41285, n41286, n41287, n41288, n41289, n41290, n41291, n41292,
         n41293, n41294, n41295, n41296, n41297, n41298, n41299, n41300,
         n41301, n41302, n41303, n41304, n41305, n41306, n41307, n41308,
         n41309, n41310, n41311, n41312, n41313, n41314, n41315, n41316,
         n41317, n41318, n41319, n41320, n41321, n41322, n41323, n41324,
         n41325, n41326, n41327, n41328, n41329, n41330, n41331, n41332,
         n41333, n41334, n41335, n41336, n41337, n41338, n41339, n41340,
         n41341, n41342, n41343, n41344, n41345, n41346, n41347, n41348,
         n41349, n41350, n41351, n41352, n41353, n41354, n41355, n41356,
         n41357, n41358, n41359, n41360, n41361, n41362, n41363, n41364,
         n41365, n41366, n41367, n41368, n41369, n41370, n41371, n41372,
         n41373, n41374, n41375, n41376, n41377, n41378, n41379, n41380,
         n41381, n41382, n41383, n41384, n41385, n41386, n41387, n41388,
         n41389, n41390, n41391, n41392, n41393, n41394, n41395, n41396,
         n41397, n41398, n41399, n41400, n41401, n41402, n41403, n41404,
         n41405, n41406, n41407, n41408, n41409, n41410, n41411, n41412,
         n41413, n41414, n41415, n41416, n41417, n41418, n41419, n41420,
         n41421, n41422, n41423, n41424, n41425, n41426, n41427, n41428,
         n41429, n41430, n41431, n41432, n41433, n41434, n41435, n41436,
         n41437, n41438, n41439, n41440, n41441, n41442, n41443, n41444,
         n41445, n41446, n41447, n41448, n41449, n41450, n41451, n41452,
         n41453, n41454, n41455, n41456, n41457, n41458, n41459, n41460,
         n41461, n41462, n41463, n41464, n41465, n41466, n41467, n41468,
         n41469, n41470, n41471, n41472, n41473, n41474, n41475, n41476,
         n41477, n41478, n41479, n41480, n41481, n41482, n41483, n41484,
         n41485, n41486, n41487, n41488, n41489, n41490, n41491, n41492,
         n41493, n41494, n41495, n41496, n41497, n41498, n41499, n41500,
         n41501, n41502, n41503, n41504, n41505, n41506, n41507, n41508,
         n41509, n41510, n41511, n41512, n41513, n41514, n41515, n41516,
         n41517, n41518, n41519, n41520, n41521, n41522, n41523, n41524,
         n41525, n41526, n41527, n41528, n41529, n41530, n41531, n41532,
         n41533, n41534, n41535, n41536, n41537, n41538, n41539, n41540,
         n41541, n41542, n41543, n41544, n41545, n41546, n41547, n41548,
         n41549, n41550, n41551, n41552, n41553, n41554, n41555, n41556,
         n41557, n41558, n41559, n41560, n41561, n41562, n41563, n41564,
         n41565, n41566, n41567, n41568, n41569, n41570, n41571, n41572,
         n41573, n41574, n41575, n41576, n41577, n41578, n41579, n41580,
         n41581, n41582, n41583, n41584, n41585, n41586, n41587, n41588,
         n41589, n41590, n41591, n41592, n41593, n41594, n41595, n41596,
         n41597, n41598, n41599, n41600, n41601, n41602, n41603, n41604,
         n41605, n41606, n41607, n41608, n41609, n41610, n41611, n41612,
         n41613, n41614, n41615, n41616, n41617, n41618, n41619, n41620,
         n41621, n41622, n41623, n41624, n41625, n41626, n41627, n41628,
         n41629, n41630, n41631, n41632, n41633, n41634, n41635, n41636,
         n41637, n41638, n41639, n41640, n41641, n41642, n41643, n41644,
         n41645, n41646, n41647, n41648, n41649, n41650, n41651, n41652,
         n41653, n41654, n41655, n41656, n41657, n41658, n41659, n41660,
         n41661, n41662, n41663, n41664, n41665, n41666, n41667, n41668,
         n41669, n41670, n41671, n41672, n41673, n41674, n41675, n41676,
         n41677, n41678, n41679, n41680, n41681, n41682, n41683, n41684,
         n41685, n41686, n41687, n41688, n41689, n41690, n41691, n41692,
         n41693, n41694, n41695, n41696, n41697, n41698, n41699, n41700,
         n41701, n41702, n41703, n41704, n41705, n41706, n41707, n41708,
         n41709, n41710, n41711, n41712, n41713, n41714, n41715, n41716,
         n41717, n41718, n41719, n41720, n41721, n41722, n41723, n41724,
         n41725, n41726, n41727, n41728, n41729, n41730, n41731, n41732,
         n41733, n41734, n41735, n41736, n41737, n41738, n41739, n41740,
         n41741, n41742, n41743, n41744, n41745, n41746, n41747, n41748,
         n41749, n41750, n41751, n41752, n41753, n41754, n41755, n41756,
         n41757, n41758, n41759, n41760, n41761, n41762, n41763, n41764,
         n41765, n41766, n41767, n41768, n41769, n41770, n41771, n41772,
         n41773, n41774, n41775, n41776, n41777, n41778, n41779, n41780,
         n41781, n41782, n41783, n41784, n41785, n41786, n41787, n41788,
         n41789, n41790, n41791, n41792, n41793, n41794, n41795, n41796,
         n41797, n41798, n41799, n41800, n41801, n41802, n41803, n41804,
         n41805, n41806, n41807, n41808, n41809, n41810, n41811, n41812,
         n41813, n41814, n41815, n41816, n41817, n41818, n41819, n41820,
         n41821, n41822, n41823, n41824, n41825, n41826, n41827, n41828,
         n41829, n41830, n41831, n41832, n41833, n41834, n41835, n41836,
         n41837, n41838, n41839, n41840, n41841, n41842, n41843, n41844,
         n41845, n41846, n41847, n41848, n41849, n41850, n41851, n41852,
         n41853, n41854, n41855, n41856, n41857, n41858, n41859, n41860,
         n41861, n41862, n41863, n41864, n41865, n41866, n41867, n41868,
         n41869, n41870, n41871, n41872, n41873, n41874, n41875, n41876,
         n41877, n41878, n41879, n41880, n41881, n41882, n41883, n41884,
         n41885, n41886, n41887, n41888, n41889, n41890, n41891, n41892,
         n41893, n41894, n41895, n41896, n41897, n41898, n41899, n41900,
         n41901, n41902, n41903, n41904, n41905, n41906, n41907, n41908,
         n41909, n41910, n41911, n41912, n41913, n41914, n41915, n41916,
         n41917, n41918, n41919, n41920, n41921, n41922, n41923, n41924,
         n41925, n41926, n41927, n41928, n41929, n41930, n41931, n41932,
         n41933, n41934, n41935, n41936, n41937, n41938, n41939, n41940,
         n41941, n41942, n41943, n41944, n41945, n41946, n41947, n41948,
         n41949, n41950, n41951, n41952, n41953, n41954, n41955, n41956,
         n41957, n41958, n41959, n41960, n41961, n41962, n41963, n41964,
         n41965, n41966, n41967, n41968, n41969, n41970, n41971, n41972,
         n41973, n41974, n41975, n41976, n41977, n41978, n41979, n41980,
         n41981, n41982, n41983, n41984, n41985, n41986, n41987, n41988,
         n41989, n41990, n41991, n41992, n41993, n41994, n41995, n41996,
         n41997, n41998, n41999, n42000, n42001, n42002, n42003, n42004,
         n42005, n42006, n42007, n42008, n42009, n42010, n42011, n42012,
         n42013, n42014, n42015, n42016, n42017, n42018, n42019, n42020,
         n42021, n42022, n42023, n42024, n42025, n42026, n42027, n42028,
         n42029, n42030, n42031, n42032, n42033, n42034, n42035, n42036,
         n42037, n42038, n42039, n42040, n42041, n42042, n42043, n42044,
         n42045, n42046, n42047, n42048, n42049, n42050, n42051, n42052,
         n42053, n42054, n42055, n42056, n42057, n42058, n42059, n42060,
         n42061, n42062, n42063, n42064, n42065, n42066, n42067, n42068,
         n42069, n42070, n42071, n42072, n42073, n42074, n42075, n42076,
         n42077, n42078, n42079, n42080, n42081, n42082, n42083, n42084,
         n42085, n42086, n42087, n42088, n42089, n42090, n42091, n42092,
         n42093, n42094, n42095, n42096, n42097, n42098, n42099, n42100,
         n42101, n42102, n42103, n42104, n42105, n42106, n42107, n42108,
         n42109, n42110, n42111, n42112, n42113, n42114, n42115, n42116,
         n42117, n42118, n42119, n42120, n42121, n42122, n42123, n42124,
         n42125, n42126, n42127, n42128, n42129, n42130, n42131, n42132,
         n42133, n42134, n42135, n42136, n42137, n42138, n42139, n42140,
         n42141, n42142, n42143, n42144, n42145, n42146, n42147, n42148,
         n42149, n42150, n42151, n42152, n42153, n42154, n42155, n42156,
         n42157, n42158, n42159, n42160, n42161, n42162, n42163, n42164,
         n42165, n42166, n42167, n42168, n42169, n42170, n42171, n42172,
         n42173, n42174, n42175, n42176, n42177, n42178, n42179, n42180,
         n42181, n42182, n42183, n42184, n42185, n42186, n42187, n42188,
         n42189, n42190, n42191, n42192, n42193, n42194, n42195, n42196,
         n42197, n42198, n42199, n42200, n42201, n42202, n42203, n42204,
         n42205, n42206, n42207, n42208, n42209, n42210, n42211, n42212,
         n42213, n42214, n42215, n42216, n42217, n42218, n42219, n42220,
         n42221, n42222, n42223, n42224, n42225, n42226, n42227, n42228,
         n42229, n42230, n42231, n42232, n42233, n42234, n42235, n42236,
         n42237, n42238, n42239, n42240, n42241, n42242, n42243, n42244,
         n42245, n42246, n42247, n42248, n42249, n42250, n42251, n42252,
         n42253, n42254, n42255, n42256, n42257, n42258, n42259, n42260,
         n42261, n42262, n42263, n42264, n42265, n42266, n42267, n42268,
         n42269, n42270, n42271, n42272, n42273, n42274, n42275, n42276,
         n42277, n42278, n42279, n42280, n42281, n42282, n42283, n42284,
         n42285, n42286, n42287, n42288, n42289, n42290, n42291, n42292,
         n42293, n42294, n42295, n42296, n42297, n42298, n42299, n42300,
         n42301, n42302, n42303, n42304, n42305, n42306, n42307, n42308,
         n42309, n42310, n42311, n42312, n42313, n42314, n42315, n42316,
         n42317, n42318, n42319, n42320, n42321, n42322, n42323, n42324,
         n42325, n42326, n42327, n42328, n42329, n42330, n42331, n42332,
         n42333, n42334, n42335, n42336, n42337, n42338, n42339, n42340,
         n42341, n42342, n42343, n42344, n42345, n42346, n42347, n42348,
         n42349, n42350, n42351, n42352, n42353, n42354, n42355, n42356,
         n42357, n42358, n42359, n42360, n42361, n42362, n42363, n42364,
         n42365, n42366, n42367, n42368, n42369, n42370, n42371, n42372,
         n42373, n42374, n42375, n42376, n42377, n42378, n42379, n42380,
         n42381, n42382, n42383, n42384, n42385, n42386, n42387, n42388,
         n42389, n42390, n42391, n42392, n42393, n42394, n42395, n42396,
         n42397, n42398, n42399, n42400, n42401, n42402, n42403, n42404,
         n42405, n42406, n42407, n42408, n42409, n42410, n42411, n42412,
         n42413, n42414, n42415, n42416, n42417, n42418, n42419, n42420,
         n42421, n42422, n42423, n42424, n42425, n42426, n42427, n42428,
         n42429, n42430, n42431, n42432, n42433, n42434, n42435, n42436,
         n42437, n42438, n42439, n42440, n42441, n42442, n42443, n42444,
         n42445, n42446, n42447, n42448, n42449, n42450, n42451, n42452,
         n42453, n42454, n42455, n42456, n42457, n42458, n42459, n42460,
         n42461, n42462, n42463, n42464, n42465, n42466, n42467, n42468,
         n42469, n42470, n42471, n42472, n42473, n42474, n42475, n42476,
         n42477, n42478, n42479, n42480, n42481, n42482, n42483, n42484,
         n42485, n42486, n42487, n42488, n42489, n42490, n42491, n42492,
         n42493, n42494, n42495, n42496, n42497, n42498, n42499, n42500,
         n42501, n42502, n42503, n42504, n42505, n42506, n42507, n42508,
         n42509, n42510, n42511, n42512, n42513, n42514, n42515, n42516,
         n42517, n42518, n42519, n42520, n42521, n42522, n42523, n42524,
         n42525, n42526, n42527, n42528, n42529, n42530, n42531, n42532,
         n42533, n42534, n42535, n42536, n42537, n42538, n42539, n42540,
         n42541, n42542, n42543, n42544, n42545, n42546, n42547, n42548,
         n42549, n42550, n42551, n42552, n42553, n42554, n42555, n42556,
         n42557, n42558, n42559, n42560, n42561, n42562, n42563, n42564,
         n42565, n42566, n42567, n42568, n42569, n42570, n42571, n42572,
         n42573, n42574, n42575, n42576, n42577, n42578, n42579, n42580,
         n42581, n42582, n42583, n42584, n42585, n42586, n42587, n42588,
         n42589, n42590, n42591, n42592, n42593, n42594, n42595, n42596,
         n42597, n42598, n42599, n42600, n42601, n42602, n42603, n42604,
         n42605, n42606, n42607, n42608, n42609, n42610, n42611, n42612,
         n42613, n42614, n42615, n42616, n42617, n42618, n42619, n42620,
         n42621, n42622, n42623, n42624, n42625, n42626, n42627, n42628,
         n42629, n42630, n42631, n42632, n42633, n42634, n42635, n42636,
         n42637, n42638, n42639, n42640, n42641, n42642, n42643, n42644,
         n42645, n42646, n42647, n42648, n42649, n42650, n42651, n42652,
         n42653, n42654, n42655, n42656, n42657, n42658, n42659, n42660,
         n42661, n42662, n42663, n42664, n42665, n42666, n42667, n42668,
         n42669, n42670, n42671, n42672, n42673, n42674, n42675, n42676,
         n42677, n42678, n42679, n42680, n42681, n42682, n42683, n42684,
         n42685, n42686, n42687, n42688, n42689, n42690, n42691, n42692,
         n42693, n42694, n42695, n42696, n42697, n42698, n42699, n42700,
         n42701, n42702, n42703, n42704, n42705, n42706, n42707, n42708,
         n42709, n42710, n42711, n42712, n42713, n42714, n42715, n42716,
         n42717, n42718, n42719, n42720, n42721, n42722, n42723, n42724,
         n42725, n42726, n42727, n42728, n42729, n42730, n42731, n42732,
         n42733, n42734, n42735, n42736, n42737, n42738, n42739, n42740,
         n42741, n42742, n42743, n42744, n42745, n42746, n42747, n42748,
         n42749, n42750, n42751, n42752, n42753, n42754, n42755, n42756,
         n42757, n42758, n42759, n42760, n42761, n42762, n42763, n42764,
         n42765, n42766, n42767, n42768, n42769, n42770, n42771, n42772,
         n42773, n42774, n42775, n42776, n42777, n42778, n42779, n42780,
         n42781, n42782, n42783, n42784, n42785, n42786, n42787, n42788,
         n42789, n42790, n42791, n42792, n42793, n42794, n42795, n42796,
         n42797, n42798, n42799, n42800, n42801, n42802, n42803, n42804,
         n42805, n42806, n42807, n42808, n42809, n42810, n42811, n42812,
         n42813, n42814, n42815, n42816, n42817, n42818, n42819, n42820,
         n42821, n42822, n42823, n42824, n42825, n42826, n42827, n42828,
         n42829, n42830, n42831, n42832, n42833, n42834, n42835, n42836,
         n42837, n42838, n42839, n42840, n42841, n42842, n42843, n42844,
         n42845, n42846, n42847, n42848, n42849, n42850, n42851, n42852,
         n42853, n42854, n42855, n42856, n42857, n42858, n42859, n42860,
         n42861, n42862, n42863, n42864, n42865, n42866, n42867, n42868,
         n42869, n42870, n42871, n42872, n42873, n42874, n42875, n42876,
         n42877, n42878, n42879, n42880, n42881, n42882, n42883, n42884,
         n42885, n42886, n42887, n42888, n42889, n42890, n42891, n42892,
         n42893, n42894, n42895, n42896, n42897, n42898, n42899, n42900,
         n42901, n42902, n42903, n42904, n42905, n42906, n42907, n42908,
         n42909, n42910, n42911, n42912, n42913, n42914, n42915, n42916,
         n42917, n42918, n42919, n42920, n42921, n42922, n42923, n42924,
         n42925, n42926, n42927, n42928, n42929, n42930, n42931, n42932,
         n42933, n42934, n42935, n42936, n42937, n42938, n42939, n42940,
         n42941, n42942, n42943, n42944, n42945, n42946, n42947, n42948,
         n42949, n42950, n42951, n42952, n42953, n42954, n42955, n42956,
         n42957, n42958, n42959, n42960, n42961, n42962, n42963, n42964,
         n42965, n42966, n42967, n42968, n42969, n42970, n42971, n42972,
         n42973, n42974, n42975, n42976, n42977, n42978, n42979, n42980,
         n42981, n42982, n42983, n42984, n42985, n42986, n42987, n42988,
         n42989, n42990, n42991, n42992, n42993, n42994, n42995, n42996,
         n42997, n42998, n42999, n43000, n43001, n43002, n43003, n43004,
         n43005, n43006, n43007, n43008, n43009, n43010, n43011, n43012,
         n43013, n43014, n43015, n43016, n43017, n43018, n43019, n43020,
         n43021, n43022, n43023, n43024, n43025, n43026, n43027, n43028,
         n43029, n43030, n43031, n43032, n43033, n43034, n43035, n43036,
         n43037, n43038, n43039, n43040, n43041, n43042, n43043, n43044,
         n43045, n43046, n43047, n43048, n43049, n43050, n43051, n43052,
         n43053, n43054, n43055, n43056, n43057, n43058, n43059, n43060,
         n43061, n43062, n43063, n43064, n43065, n43066, n43067, n43068,
         n43069, n43070, n43071, n43072, n43073, n43074, n43075, n43076,
         n43077, n43078, n43079, n43080, n43081, n43082, n43083, n43084,
         n43085, n43086, n43087, n43088, n43089, n43090, n43091, n43092,
         n43093, n43094, n43095, n43096, n43097, n43098, n43099, n43100,
         n43101, n43102, n43103, n43104, n43105, n43106, n43107, n43108,
         n43109, n43110, n43111, n43112, n43113, n43114, n43115, n43116,
         n43117, n43118, n43119, n43120, n43121, n43122, n43123, n43124,
         n43125, n43126, n43127, n43128, n43129, n43130, n43131, n43132,
         n43133, n43134, n43135, n43136, n43137, n43138, n43139, n43140,
         n43141, n43142, n43143, n43144, n43145, n43146, n43147, n43148,
         n43149, n43150, n43151, n43152, n43153, n43154, n43155, n43156,
         n43157, n43158, n43159, n43160, n43161, n43162, n43163, n43164,
         n43165, n43166, n43167, n43168, n43169, n43170, n43171, n43172,
         n43173, n43174, n43175, n43176, n43177, n43178, n43179, n43180,
         n43181, n43182, n43183, n43184, n43185, n43186, n43187, n43188,
         n43189, n43190, n43191, n43192, n43193, n43194, n43195, n43196,
         n43197, n43198, n43199, n43200, n43201, n43202, n43203, n43204,
         n43205, n43206, n43207, n43208, n43209, n43210, n43211, n43212,
         n43213, n43214, n43215, n43216, n43217, n43218, n43219, n43220,
         n43221, n43222, n43223, n43224, n43225, n43226, n43227, n43228,
         n43229, n43230, n43231, n43232, n43233, n43234, n43235, n43236,
         n43237, n43238, n43239, n43240, n43241, n43242, n43243, n43244,
         n43245, n43246, n43247, n43248, n43249, n43250, n43251, n43252,
         n43253, n43254, n43255, n43256, n43257, n43258, n43259, n43260,
         n43261, n43262, n43263, n43264, n43265, n43266, n43267, n43268,
         n43269, n43270, n43271, n43272, n43273, n43274, n43275, n43276,
         n43277, n43278, n43279, n43280, n43281, n43282, n43283, n43284,
         n43285, n43286, n43287, n43288, n43289, n43290, n43291, n43292,
         n43293, n43294, n43295, n43296, n43297, n43298, n43299, n43300,
         n43301, n43302, n43303, n43304, n43305, n43306, n43307, n43308,
         n43309, n43310, n43311, n43312, n43313, n43314, n43315, n43316,
         n43317, n43318, n43319, n43320, n43321, n43322, n43323, n43324,
         n43325, n43326, n43327, n43328, n43329, n43330, n43331, n43332,
         n43333, n43334, n43335, n43336, n43337, n43338, n43339, n43340,
         n43341, n43342, n43343, n43344, n43345, n43346, n43347, n43348,
         n43349, n43350, n43351, n43352, n43353, n43354, n43355, n43356,
         n43357, n43358, n43359, n43360, n43361, n43362, n43363, n43364,
         n43365, n43366, n43367, n43368, n43369, n43370, n43371, n43372,
         n43373, n43374, n43375, n43376, n43377, n43378, n43379, n43380,
         n43381, n43382, n43383, n43384, n43385, n43386, n43387, n43388,
         n43389, n43390, n43391, n43392, n43393, n43394, n43395, n43396,
         n43397, n43398, n43399, n43400, n43401, n43402, n43403, n43404,
         n43405, n43406, n43407, n43408, n43409, n43410, n43411, n43412,
         n43413, n43414, n43415, n43416, n43417, n43418, n43419, n43420,
         n43421, n43422, n43423, n43424, n43425, n43426, n43427, n43428,
         n43429, n43430, n43431, n43432, n43433, n43434, n43435, n43436,
         n43437, n43438, n43439, n43440, n43441, n43442, n43443, n43444,
         n43445, n43446, n43447, n43448, n43449, n43450, n43451, n43452,
         n43453, n43454, n43455, n43456, n43457, n43458, n43459, n43460,
         n43461, n43462, n43463, n43464, n43465, n43466, n43467, n43468,
         n43469, n43470, n43471, n43472, n43473, n43474, n43475, n43476,
         n43477, n43478, n43479, n43480, n43481, n43482, n43483, n43484,
         n43485, n43486, n43487, n43488, n43489, n43490, n43491, n43492,
         n43493, n43494, n43495, n43496, n43497, n43498, n43499, n43500,
         n43501, n43502, n43503, n43504, n43505, n43506, n43507, n43508,
         n43509, n43510, n43511, n43512, n43513, n43514, n43515, n43516,
         n43517, n43518, n43519, n43520, n43521, n43522, n43523, n43524,
         n43525, n43526, n43527, n43528, n43529, n43530, n43531, n43532,
         n43533, n43534, n43535, n43536, n43537, n43538, n43539, n43540,
         n43541, n43542, n43543, n43544, n43545, n43546, n43547, n43548,
         n43549, n43550, n43551, n43552, n43553, n43554, n43555, n43556,
         n43557, n43558, n43559, n43560, n43561, n43562, n43563, n43564,
         n43565, n43566, n43567, n43568, n43569, n43570, n43571, n43572,
         n43573, n43574, n43575, n43576, n43577, n43578, n43579, n43580,
         n43581, n43582, n43583, n43584, n43585, n43586, n43587, n43588,
         n43589, n43590, n43591, n43592, n43593, n43594, n43595, n43596,
         n43597, n43598, n43599, n43600, n43601, n43602, n43603, n43604,
         n43605, n43606, n43607, n43608, n43609, n43610, n43611, n43612,
         n43613, n43614, n43615, n43616, n43617, n43618, n43619, n43620,
         n43621, n43622, n43623, n43624, n43625, n43626, n43627, n43628,
         n43629, n43630, n43631, n43632, n43633, n43634, n43635, n43636,
         n43637, n43638, n43639, n43640, n43641, n43642, n43643, n43644,
         n43645, n43646, n43647, n43648, n43649, n43650, n43651, n43652,
         n43653, n43654, n43655, n43656, n43657, n43658, n43659, n43660,
         n43661, n43662, n43663, n43664, n43665, n43666, n43667, n43668,
         n43669, n43670, n43671, n43672, n43673, n43674, n43675, n43676,
         n43677, n43678, n43679, n43680, n43681, n43682, n43683, n43684,
         n43685, n43686, n43687, n43688, n43689, n43690, n43691, n43692,
         n43693, n43694, n43695, n43696, n43697, n43698, n43699, n43700,
         n43701, n43702, n43703, n43704, n43705, n43706, n43707, n43708,
         n43709, n43710, n43711, n43712, n43713, n43714, n43715, n43716,
         n43717, n43718, n43719, n43720, n43721, n43722, n43723, n43724,
         n43725, n43726, n43727, n43728, n43729, n43730, n43731, n43732,
         n43733, n43734, n43735, n43736, n43737, n43738, n43739, n43740,
         n43741, n43742, n43743, n43744, n43745, n43746, n43747, n43748,
         n43749, n43750, n43751, n43752, n43753, n43754, n43755, n43756,
         n43757, n43758, n43759, n43760, n43761, n43762, n43763, n43764,
         n43765, n43766, n43767, n43768, n43769, n43770, n43771, n43772,
         n43773, n43774, n43775, n43776, n43777, n43778, n43779, n43780,
         n43781, n43782, n43783, n43784, n43785, n43786, n43787, n43788,
         n43789, n43790, n43791, n43792, n43793, n43794, n43795, n43796,
         n43797, n43798, n43799, n43800, n43801, n43802, n43803, n43804,
         n43805, n43806, n43807, n43808, n43809, n43810, n43811, n43812,
         n43813, n43814, n43815, n43816, n43817, n43818, n43819, n43820,
         n43821, n43822, n43823, n43824, n43825, n43826, n43827, n43828,
         n43829, n43830, n43831, n43832, n43833, n43834, n43835, n43836,
         n43837, n43838, n43839, n43840, n43841, n43842, n43843, n43844,
         n43845, n43846, n43847, n43848, n43849, n43850, n43851, n43852,
         n43853, n43854, n43855, n43856, n43857, n43858, n43859, n43860,
         n43861, n43862, n43863, n43864, n43865, n43866, n43867, n43868,
         n43869, n43870, n43871, n43872, n43873, n43874, n43875, n43876,
         n43877, n43878, n43879, n43880, n43881, n43882, n43883, n43884,
         n43885, n43886, n43887, n43888, n43889, n43890, n43891, n43892,
         n43893, n43894, n43895, n43896, n43897, n43898, n43899, n43900,
         n43901, n43902, n43903, n43904, n43905, n43906, n43907, n43908,
         n43909, n43910, n43911, n43912, n43913, n43914, n43915, n43916,
         n43917, n43918, n43919, n43920, n43921, n43922, n43923, n43924,
         n43925, n43926, n43927, n43928, n43929, n43930, n43931, n43932,
         n43933, n43934, n43935, n43936, n43937, n43938, n43939, n43940,
         n43941, n43942, n43943, n43944, n43945, n43946, n43947, n43948,
         n43949, n43950, n43951, n43952, n43953, n43954, n43955, n43956,
         n43957, n43958, n43959, n43960, n43961, n43962, n43963, n43964,
         n43965, n43966, n43967, n43968, n43969, n43970, n43971, n43972,
         n43973, n43974, n43975, n43976, n43977, n43978, n43979, n43980,
         n43981, n43982, n43983, n43984, n43985, n43986, n43987, n43988,
         n43989, n43990, n43991, n43992, n43993, n43994, n43995, n43996,
         n43997, n43998, n43999, n44000, n44001, n44002, n44003, n44004,
         n44005, n44006, n44007, n44008, n44009, n44010, n44011, n44012,
         n44013, n44014, n44015, n44016, n44017, n44018, n44019, n44020,
         n44021, n44022, n44023, n44024, n44025, n44026, n44027, n44028,
         n44029, n44030, n44031, n44032, n44033, n44034, n44035, n44036,
         n44037, n44038, n44039, n44040, n44041, n44042, n44043, n44044,
         n44045, n44046, n44047, n44048, n44049, n44050, n44051, n44052,
         n44053, n44054, n44055, n44056, n44057, n44058, n44059, n44060,
         n44061, n44062, n44063, n44064, n44065, n44066, n44067, n44068,
         n44069, n44070, n44071, n44072, n44073, n44074, n44075, n44076,
         n44077, n44078, n44079, n44080, n44081, n44082, n44083, n44084,
         n44085, n44086, n44087, n44088, n44089, n44090, n44091, n44092,
         n44093, n44094, n44095, n44096, n44097, n44098, n44099, n44100,
         n44101, n44102, n44103, n44104, n44105, n44106, n44107, n44108,
         n44109, n44110, n44111, n44112, n44113, n44114, n44115, n44116,
         n44117, n44118, n44119, n44120, n44121, n44122, n44123, n44124,
         n44125, n44126, n44127, n44128, n44129, n44130, n44131, n44132,
         n44133, n44134, n44135, n44136, n44137, n44138, n44139, n44140,
         n44141, n44142, n44143, n44144, n44145, n44146, n44147, n44148,
         n44149, n44150, n44151, n44152, n44153, n44154, n44155, n44156,
         n44157, n44158, n44159, n44160, n44161, n44162, n44163, n44164,
         n44165, n44166, n44167, n44168, n44169, n44170, n44171, n44172,
         n44173, n44174, n44175, n44176, n44177, n44178, n44179, n44180,
         n44181, n44182, n44183, n44184, n44185, n44186, n44187, n44188,
         n44189, n44190, n44191, n44192, n44193, n44194, n44195, n44196,
         n44197, n44198, n44199, n44200, n44201, n44202, n44203, n44204,
         n44205, n44206, n44207, n44208, n44209, n44210, n44211, n44212,
         n44213, n44214, n44215, n44216, n44217, n44218, n44219, n44220,
         n44221, n44222, n44223, n44224, n44225, n44226, n44227, n44228,
         n44229, n44230, n44231, n44232, n44233, n44234, n44235, n44236,
         n44237, n44238, n44239, n44240, n44241, n44242, n44243, n44244,
         n44245, n44246, n44247, n44248, n44249, n44250, n44251, n44252,
         n44253, n44254, n44255, n44256, n44257, n44258, n44259, n44260,
         n44261, n44262, n44263, n44264, n44265, n44266, n44267, n44268,
         n44269, n44270, n44271, n44272, n44273, n44274, n44275, n44276,
         n44277, n44278, n44279, n44280, n44281, n44282, n44283, n44284,
         n44285, n44286, n44287, n44288, n44289, n44290, n44291, n44292,
         n44293, n44294, n44295, n44296, n44297, n44298, n44299, n44300,
         n44301, n44302, n44303, n44304, n44305, n44306, n44307, n44308,
         n44309, n44310, n44311, n44312, n44313, n44314, n44315, n44316,
         n44317, n44318, n44319, n44320, n44321, n44322, n44323, n44324,
         n44325, n44326, n44327, n44328, n44329, n44330, n44331, n44332,
         n44333, n44334, n44335, n44336, n44337, n44338, n44339, n44340,
         n44341, n44342, n44343, n44344, n44345, n44346, n44347, n44348,
         n44349, n44350, n44351, n44352, n44353, n44354, n44355, n44356,
         n44357, n44358, n44359, n44360, n44361, n44362, n44363, n44364,
         n44365, n44366, n44367, n44368, n44369, n44370, n44371, n44372,
         n44373, n44374, n44375, n44376, n44377, n44378, n44379, n44380,
         n44381, n44382, n44383, n44384, n44385, n44386, n44387, n44388,
         n44389, n44390, n44391, n44392, n44393, n44394, n44395, n44396,
         n44397, n44398, n44399, n44400, n44401, n44402, n44403, n44404,
         n44405, n44406, n44407, n44408, n44409, n44410, n44411, n44412,
         n44413, n44414, n44415, n44416, n44417, n44418, n44419, n44420,
         n44421, n44422, n44423, n44424, n44425, n44426, n44427, n44428,
         n44429, n44430, n44431, n44432, n44433, n44434, n44435, n44436,
         n44437, n44438, n44439, n44440, n44441, n44442, n44443, n44444,
         n44445, n44446, n44447, n44448, n44449, n44450, n44451, n44452,
         n44453, n44454, n44455, n44456, n44457, n44458, n44459, n44460,
         n44461, n44462, n44463, n44464, n44465, n44466, n44467, n44468,
         n44469, n44470, n44471, n44472, n44473, n44474, n44475, n44476,
         n44477, n44478, n44479, n44480, n44481, n44482, n44483, n44484,
         n44485, n44486, n44487, n44488, n44489, n44490, n44491, n44492,
         n44493, n44494, n44495, n44496, n44497, n44498, n44499, n44500,
         n44501, n44502, n44503, n44504, n44505, n44506, n44507, n44508,
         n44509, n44510, n44511, n44512, n44513, n44514, n44515, n44516,
         n44517, n44518, n44519, n44520, n44521, n44522, n44523, n44524,
         n44525, n44526, n44527, n44528, n44529, n44530, n44531, n44532,
         n44533, n44534, n44535, n44536, n44537, n44538, n44539, n44540,
         n44541, n44542, n44543, n44544, n44545, n44546, n44547, n44548,
         n44549, n44550, n44551, n44552, n44553, n44554, n44555, n44556,
         n44557, n44558, n44559, n44560, n44561, n44562, n44563, n44564,
         n44565, n44566, n44567, n44568, n44569, n44570, n44571, n44572,
         n44573, n44574, n44575, n44576, n44577, n44578, n44579, n44580,
         n44581, n44582, n44583, n44584, n44585, n44586, n44587, n44588,
         n44589, n44590, n44591, n44592, n44593, n44594, n44595, n44596,
         n44597, n44598, n44599, n44600, n44601, n44602, n44603, n44604,
         n44605, n44606, n44607, n44608, n44609, n44610, n44611, n44612,
         n44613, n44614, n44615, n44616, n44617, n44618, n44619, n44620,
         n44621, n44622, n44623, n44624, n44625, n44626, n44627, n44628,
         n44629, n44630, n44631, n44632, n44633, n44634, n44635, n44636,
         n44637, n44638, n44639, n44640, n44641, n44642, n44643, n44644,
         n44645, n44646, n44647, n44648, n44649, n44650, n44651, n44652,
         n44653, n44654, n44655, n44656, n44657, n44658, n44659, n44660,
         n44661, n44662, n44663, n44664, n44665, n44666, n44667, n44668,
         n44669, n44670, n44671, n44672, n44673, n44674, n44675, n44676,
         n44677, n44678, n44679, n44680, n44681, n44682, n44683, n44684,
         n44685, n44686, n44687, n44688, n44689, n44690, n44691, n44692,
         n44693, n44694, n44695, n44696, n44697, n44698, n44699, n44700,
         n44701, n44702, n44703, n44704, n44705, n44706, n44707, n44708,
         n44709, n44710, n44711, n44712, n44713, n44714, n44715, n44716,
         n44717, n44718, n44719, n44720, n44721, n44722, n44723, n44724,
         n44725, n44726, n44727, n44728, n44729, n44730, n44731, n44732,
         n44733, n44734, n44735, n44736, n44737, n44738, n44739, n44740,
         n44741, n44742, n44743, n44744, n44745, n44746, n44747, n44748,
         n44749, n44750, n44751, n44752, n44753, n44754, n44755, n44756,
         n44757, n44758, n44759, n44760, n44761, n44762, n44763, n44764,
         n44765, n44766, n44767, n44768, n44769, n44770, n44771, n44772,
         n44773, n44774, n44775, n44776, n44777, n44778, n44779, n44780,
         n44781, n44782, n44783, n44784, n44785, n44786, n44787, n44788,
         n44789, n44790, n44791, n44792, n44793, n44794, n44795, n44796,
         n44797, n44798, n44799, n44800, n44801, n44802, n44803, n44804,
         n44805, n44806, n44807, n44808, n44809, n44810, n44811, n44812,
         n44813, n44814, n44815, n44816, n44817, n44818, n44819, n44820,
         n44821, n44822, n44823, n44824, n44825, n44826, n44827, n44828,
         n44829, n44830, n44831, n44832, n44833, n44834, n44835, n44836,
         n44837, n44838, n44839, n44840, n44841, n44842, n44843, n44844,
         n44845, n44846, n44847, n44848, n44849, n44850, n44851, n44852,
         n44853, n44854, n44855, n44856, n44857, n44858, n44859, n44860,
         n44861, n44862, n44863, n44864, n44865, n44866, n44867, n44868,
         n44869, n44870, n44871, n44872, n44873, n44874, n44875, n44876,
         n44877, n44878, n44879, n44880, n44881, n44882, n44883, n44884,
         n44885, n44886, n44887, n44888, n44889, n44890, n44891, n44892,
         n44893, n44894, n44895, n44896, n44897, n44898, n44899, n44900,
         n44901, n44902, n44903, n44904, n44905, n44906, n44907, n44908,
         n44909, n44910, n44911, n44912, n44913, n44914, n44915, n44916,
         n44917, n44918, n44919, n44920, n44921, n44922, n44923, n44924,
         n44925, n44926, n44927, n44928, n44929, n44930, n44931, n44932,
         n44933, n44934, n44935, n44936, n44937, n44938, n44939, n44940,
         n44941, n44942, n44943, n44944, n44945, n44946, n44947, n44948,
         n44949, n44950, n44951, n44952, n44953, n44954, n44955, n44956,
         n44957, n44958, n44959, n44960, n44961, n44962, n44963, n44964,
         n44965, n44966, n44967, n44968, n44969, n44970, n44971, n44972,
         n44973, n44974, n44975, n44976, n44977, n44978, n44979, n44980,
         n44981, n44982, n44983, n44984, n44985, n44986, n44987, n44988,
         n44989, n44990, n44991, n44992, n44993, n44994, n44995, n44996,
         n44997, n44998, n44999, n45000, n45001, n45002, n45003, n45004,
         n45005, n45006, n45007, n45008, n45009, n45010, n45011, n45012,
         n45013, n45014, n45015, n45016, n45017, n45018, n45019, n45020,
         n45021, n45022, n45023, n45024, n45025, n45026, n45027, n45028,
         n45029, n45030, n45031, n45032, n45033, n45034, n45035, n45036,
         n45037, n45038, n45039, n45040, n45041, n45042, n45043, n45044,
         n45045, n45046, n45047, n45048, n45049, n45050, n45051, n45052,
         n45053, n45054, n45055, n45056, n45057, n45058, n45059, n45060,
         n45061, n45062, n45063, n45064, n45065, n45066, n45067, n45068,
         n45069, n45070, n45071, n45072, n45073, n45074, n45075, n45076,
         n45077, n45078, n45079, n45080, n45081, n45082, n45083, n45084,
         n45085, n45086, n45087, n45088, n45089, n45090, n45091, n45092,
         n45093, n45094, n45095, n45096, n45097, n45098, n45099, n45100,
         n45101, n45102, n45103, n45104, n45105, n45106, n45107, n45108,
         n45109, n45110, n45111, n45112, n45113, n45114, n45115, n45116,
         n45117, n45118, n45119, n45120, n45121, n45122, n45123, n45124,
         n45125, n45126, n45127, n45128, n45129, n45130, n45131, n45132,
         n45133, n45134, n45135, n45136, n45137, n45138, n45139, n45140,
         n45141, n45142, n45143, n45144, n45145, n45146, n45147, n45148,
         n45149, n45150, n45151, n45152, n45153, n45154, n45155, n45156,
         n45157, n45158, n45159, n45160, n45161, n45162, n45163, n45164,
         n45165, n45166, n45167, n45168, n45169, n45170, n45171, n45172,
         n45173, n45174, n45175, n45176, n45177, n45178, n45179, n45180,
         n45181, n45182, n45183, n45184, n45185, n45186, n45187, n45188,
         n45189, n45190, n45191, n45192, n45193, n45194, n45195, n45196,
         n45197, n45198, n45199, n45200, n45201, n45202, n45203, n45204,
         n45205, n45206, n45207, n45208, n45209, n45210, n45211, n45212,
         n45213, n45214, n45215, n45216, n45217, n45218, n45219, n45220,
         n45221, n45222, n45223, n45224, n45225, n45226, n45227, n45228,
         n45229, n45230, n45231, n45232, n45233, n45234, n45235, n45236,
         n45237, n45238, n45239, n45240, n45241, n45242, n45243, n45244,
         n45245, n45246, n45247, n45248, n45249, n45250, n45251, n45252,
         n45253, n45254, n45255, n45256, n45257, n45258, n45259, n45260,
         n45261, n45262, n45263, n45264, n45265, n45266, n45267, n45268,
         n45269, n45270, n45271, n45272, n45273, n45274, n45275, n45276,
         n45277, n45278, n45279, n45280, n45281, n45282, n45283, n45284,
         n45285, n45286, n45287, n45288, n45289, n45290, n45291, n45292,
         n45293, n45294, n45295, n45296, n45297, n45298, n45299, n45300,
         n45301, n45302, n45303, n45304, n45305, n45306, n45307, n45308,
         n45309, n45310, n45311, n45312, n45313, n45314, n45315, n45316,
         n45317, n45318, n45319, n45320, n45321, n45322, n45323, n45324,
         n45325, n45326, n45327, n45328, n45329, n45330, n45331, n45332,
         n45333, n45334, n45335, n45336, n45337, n45338, n45339, n45340,
         n45341, n45342, n45343, n45344, n45345, n45346, n45347, n45348,
         n45349, n45350, n45351, n45352, n45353, n45354, n45355, n45356,
         n45357, n45358, n45359, n45360, n45361, n45362, n45363, n45364,
         n45365, n45366, n45367, n45368, n45369, n45370, n45371, n45372,
         n45373, n45374, n45375, n45376, n45377, n45378, n45379, n45380,
         n45381, n45382, n45383, n45384, n45385, n45386, n45387, n45388,
         n45389, n45390, n45391, n45392, n45393, n45394, n45395, n45396,
         n45397, n45398, n45399, n45400, n45401, n45402, n45403, n45404,
         n45405, n45406, n45407, n45408, n45409, n45410, n45411, n45412,
         n45413, n45414, n45415, n45416, n45417, n45418, n45419, n45420,
         n45421, n45422, n45423, n45424, n45425, n45426, n45427, n45428,
         n45429, n45430, n45431, n45432, n45433, n45434, n45435, n45436,
         n45437, n45438, n45439, n45440, n45441, n45442, n45443, n45444,
         n45445, n45446, n45447, n45448, n45449, n45450, n45451, n45452,
         n45453, n45454, n45455, n45456, n45457, n45458, n45459, n45460,
         n45461, n45462, n45463, n45464, n45465, n45466, n45467, n45468,
         n45469, n45470, n45471, n45472, n45473, n45474, n45475, n45476,
         n45477, n45478, n45479, n45480, n45481, n45482, n45483, n45484,
         n45485, n45486, n45487, n45488, n45489, n45490, n45491, n45492,
         n45493, n45494, n45495, n45496, n45497, n45498, n45499, n45500,
         n45501, n45502, n45503, n45504, n45505, n45506, n45507, n45508,
         n45509, n45510, n45511, n45512, n45513, n45514, n45515, n45516,
         n45517, n45518, n45519, n45520, n45521, n45522, n45523, n45524,
         n45525, n45526, n45527, n45528, n45529, n45530, n45531, n45532,
         n45533, n45534, n45535, n45536, n45537, n45538, n45539, n45540,
         n45541, n45542, n45543, n45544, n45545, n45546, n45547, n45548,
         n45549, n45550, n45551, n45552, n45553, n45554, n45555, n45556,
         n45557, n45558, n45559, n45560, n45561, n45562, n45563, n45564,
         n45565, n45566, n45567, n45568, n45569, n45570, n45571, n45572,
         n45573, n45574, n45575, n45576, n45577, n45578, n45579, n45580,
         n45581, n45582, n45583, n45584, n45585, n45586, n45587, n45588,
         n45589, n45590, n45591, n45592, n45593, n45594, n45595, n45596,
         n45597, n45598, n45599, n45600, n45601, n45602, n45603, n45604,
         n45605, n45606, n45607, n45608, n45609, n45610, n45611, n45612,
         n45613, n45614, n45615, n45616, n45617, n45618, n45619, n45620,
         n45621, n45622, n45623, n45624, n45625, n45626, n45627, n45628,
         n45629, n45630, n45631, n45632, n45633, n45634, n45635, n45636,
         n45637, n45638, n45639, n45640, n45641, n45642, n45643, n45644,
         n45645, n45646, n45647, n45648, n45649, n45650, n45651, n45652,
         n45653, n45654, n45655, n45656, n45657, n45658, n45659, n45660,
         n45661, n45662, n45663, n45664, n45665, n45666, n45667, n45668,
         n45669, n45670, n45671, n45672, n45673, n45674, n45675, n45676,
         n45677, n45678, n45679, n45680, n45681, n45682, n45683, n45684,
         n45685, n45686, n45687, n45688, n45689, n45690, n45691, n45692,
         n45693, n45694, n45695, n45696, n45697, n45698, n45699, n45700,
         n45701, n45702, n45703, n45704, n45705, n45706, n45707, n45708,
         n45709, n45710, n45711, n45712, n45713, n45714, n45715, n45716,
         n45717, n45718, n45719, n45720, n45721, n45722, n45723, n45724,
         n45725, n45726, n45727, n45728, n45729, n45730, n45731, n45732,
         n45733, n45734, n45735, n45736, n45737, n45738, n45739, n45740,
         n45741, n45742, n45743, n45744, n45745, n45746, n45747, n45748,
         n45749, n45750, n45751, n45752, n45753, n45754, n45755, n45756,
         n45757, n45758, n45759, n45760, n45761, n45762, n45763, n45764,
         n45765, n45766, n45767, n45768, n45769, n45770, n45771, n45772,
         n45773, n45774, n45775, n45776, n45777, n45778, n45779, n45780,
         n45781, n45782, n45783, n45784, n45785, n45786, n45787, n45788,
         n45789, n45790, n45791, n45792, n45793, n45794, n45795, n45796,
         n45797, n45798, n45799, n45800, n45801, n45802, n45803, n45804,
         n45805, n45806, n45807, n45808, n45809, n45810, n45811, n45812,
         n45813, n45814, n45815, n45816, n45817, n45818, n45819, n45820,
         n45821, n45822, n45823, n45824, n45825, n45826, n45827, n45828,
         n45829, n45830, n45831, n45832, n45833, n45834, n45835, n45836,
         n45837, n45838, n45839, n45840, n45841, n45842, n45843, n45844,
         n45845, n45846, n45847, n45848, n45849, n45850, n45851, n45852,
         n45853, n45854, n45855, n45856, n45857, n45858, n45859, n45860,
         n45861, n45862, n45863, n45864, n45865, n45866, n45867, n45868,
         n45869, n45870, n45871, n45872, n45873, n45874, n45875, n45876,
         n45877, n45878, n45879, n45880, n45881, n45882, n45883, n45884,
         n45885, n45886, n45887, n45888, n45889, n45890, n45891, n45892,
         n45893, n45894, n45895, n45896, n45897, n45898, n45899, n45900,
         n45901, n45902, n45903, n45904, n45905, n45906, n45907, n45908,
         n45909, n45910, n45911, n45912, n45913, n45914, n45915, n45916,
         n45917, n45918, n45919, n45920, n45921, n45922, n45923, n45924,
         n45925, n45926, n45927, n45928, n45929, n45930, n45931, n45932,
         n45933, n45934, n45935, n45936, n45937, n45938, n45939, n45940,
         n45941, n45942, n45943, n45944, n45945, n45946, n45947, n45948,
         n45949, n45950, n45951, n45952, n45953, n45954, n45955, n45956,
         n45957, n45958, n45959, n45960, n45961, n45962, n45963, n45964,
         n45965, n45966, n45967, n45968, n45969, n45970, n45971, n45972,
         n45973, n45974, n45975, n45976, n45977, n45978, n45979, n45980,
         n45981, n45982, n45983, n45984, n45985, n45986, n45987, n45988,
         n45989, n45990, n45991, n45992, n45993, n45994, n45995, n45996,
         n45997, n45998, n45999, n46000, n46001, n46002, n46003, n46004,
         n46005, n46006, n46007, n46008, n46009, n46010, n46011, n46012,
         n46013, n46014, n46015, n46016, n46017, n46018, n46019, n46020,
         n46021, n46022, n46023, n46024, n46025, n46026, n46027, n46028,
         n46029, n46030, n46031, n46032, n46033, n46034, n46035, n46036,
         n46037, n46038, n46039, n46040, n46041, n46042, n46043, n46044,
         n46045, n46046, n46047, n46048, n46049, n46050, n46051, n46052,
         n46053, n46054, n46055, n46056, n46057, n46058, n46059, n46060,
         n46061, n46062, n46063, n46064, n46065, n46066, n46067, n46068,
         n46069, n46070, n46071, n46072, n46073, n46074, n46075, n46076,
         n46077, n46078, n46079, n46080, n46081, n46082, n46083, n46084,
         n46085, n46086, n46087, n46088, n46089, n46090, n46091, n46092,
         n46093, n46094, n46095, n46096, n46097, n46098, n46099, n46100,
         n46101, n46102, n46103, n46104, n46105, n46106, n46107, n46108,
         n46109, n46110, n46111, n46112, n46113, n46114, n46115, n46116,
         n46117, n46118, n46119, n46120, n46121, n46122, n46123, n46124,
         n46125, n46126, n46127, n46128, n46129, n46130, n46131, n46132,
         n46133, n46134, n46135, n46136, n46137, n46138, n46139, n46140,
         n46141, n46142, n46143, n46144, n46145, n46146, n46147, n46148,
         n46149, n46150, n46151, n46152, n46153, n46154, n46155, n46156,
         n46157, n46158, n46159, n46160, n46161, n46162, n46163, n46164,
         n46165, n46166, n46167, n46168, n46169, n46170, n46171, n46172,
         n46173, n46174, n46175, n46176, n46177, n46178, n46179, n46180,
         n46181, n46182, n46183, n46184, n46185, n46186, n46187, n46188,
         n46189, n46190, n46191, n46192, n46193, n46194, n46195, n46196,
         n46197, n46198, n46199, n46200, n46201, n46202, n46203, n46204,
         n46205, n46206, n46207, n46208, n46209, n46210, n46211, n46212,
         n46213, n46214, n46215, n46216, n46217, n46218, n46219, n46220,
         n46221, n46222, n46223, n46224, n46225, n46226, n46227, n46228,
         n46229, n46230, n46231, n46232, n46233, n46234, n46235, n46236,
         n46237, n46238, n46239, n46240, n46241, n46242, n46243, n46244,
         n46245, n46246, n46247, n46248, n46249, n46250, n46251, n46252,
         n46253, n46254, n46255, n46256, n46257, n46258, n46259, n46260,
         n46261, n46262, n46263, n46264, n46265, n46266, n46267, n46268,
         n46269, n46270, n46271, n46272, n46273, n46274, n46275, n46276,
         n46277, n46278, n46279, n46280, n46281, n46282, n46283, n46284,
         n46285, n46286, n46287, n46288, n46289, n46290, n46291, n46292,
         n46293, n46294, n46295, n46296, n46297, n46298, n46299, n46300,
         n46301, n46302, n46303, n46304, n46305, n46306, n46307, n46308,
         n46309, n46310, n46311, n46312, n46313, n46314, n46315, n46316,
         n46317, n46318, n46319, n46320, n46321, n46322, n46323, n46324,
         n46325, n46326, n46327, n46328, n46329, n46330, n46331, n46332,
         n46333, n46334, n46335, n46336, n46337, n46338, n46339, n46340,
         n46341, n46342, n46343, n46344, n46345, n46346, n46347, n46348,
         n46349, n46350, n46351, n46352, n46353, n46354, n46355, n46356,
         n46357, n46358, n46359, n46360, n46361, n46362, n46363, n46364,
         n46365, n46366, n46367, n46368, n46369, n46370, n46371, n46372,
         n46373, n46374, n46375, n46376, n46377, n46378, n46379, n46380,
         n46381, n46382, n46383, n46384, n46385, n46386, n46387, n46388,
         n46389, n46390, n46391, n46392, n46393, n46394, n46395, n46396,
         n46397, n46398, n46399, n46400, n46401, n46402, n46403, n46404,
         n46405, n46406, n46407, n46408, n46409, n46410, n46411, n46412,
         n46413, n46414, n46415, n46416, n46417, n46418, n46419, n46420,
         n46421, n46422, n46423, n46424, n46425, n46426, n46427, n46428,
         n46429, n46430, n46431, n46432, n46433, n46434, n46435, n46436,
         n46437, n46438, n46439, n46440, n46441, n46442, n46443, n46444,
         n46445, n46446, n46447, n46448, n46449, n46450, n46451, n46452,
         n46453, n46454, n46455, n46456, n46457, n46458, n46459, n46460,
         n46461, n46462, n46463, n46464, n46465, n46466, n46467, n46468,
         n46469, n46470, n46471, n46472, n46473, n46474, n46475, n46476,
         n46477, n46478, n46479, n46480, n46481, n46482, n46483, n46484,
         n46485, n46486, n46487, n46488, n46489, n46490, n46491, n46492,
         n46493, n46494, n46495, n46496, n46497, n46498, n46499, n46500,
         n46501, n46502, n46503, n46504, n46505, n46506, n46507, n46508,
         n46509, n46510, n46511, n46512, n46513, n46514, n46515, n46516,
         n46517, n46518, n46519, n46520, n46521, n46522, n46523, n46524,
         n46525, n46526, n46527, n46528, n46529, n46530, n46531, n46532,
         n46533, n46534, n46535, n46536, n46537, n46538, n46539, n46540,
         n46541, n46542, n46543, n46544, n46545, n46546, n46547, n46548,
         n46549, n46550, n46551, n46552, n46553, n46554, n46555, n46556,
         n46557, n46558, n46559, n46560, n46561, n46562, n46563, n46564,
         n46565, n46566, n46567, n46568, n46569, n46570, n46571, n46572,
         n46573, n46574, n46575, n46576, n46577, n46578, n46579, n46580,
         n46581, n46582, n46583, n46584, n46585, n46586, n46587, n46588,
         n46589, n46590, n46591, n46592, n46593, n46594, n46595, n46596,
         n46597, n46598, n46599, n46600, n46601, n46602, n46603, n46604,
         n46605, n46606, n46607, n46608, n46609, n46610, n46611, n46612,
         n46613, n46614, n46615, n46616, n46617, n46618, n46619, n46620,
         n46621, n46622, n46623, n46624, n46625, n46626, n46627, n46628,
         n46629, n46630, n46631, n46632, n46633, n46634, n46635, n46636,
         n46637, n46638, n46639, n46640, n46641, n46642, n46643, n46644,
         n46645, n46646, n46647, n46648, n46649, n46650, n46651, n46652,
         n46653, n46654, n46655, n46656, n46657, n46658, n46659, n46660,
         n46661, n46662, n46663, n46664, n46665, n46666, n46667, n46668,
         n46669, n46670, n46671, n46672, n46673, n46674, n46675, n46676,
         n46677, n46678, n46679, n46680, n46681, n46682, n46683, n46684,
         n46685, n46686, n46687, n46688, n46689, n46690, n46691, n46692,
         n46693, n46694, n46695, n46696, n46697, n46698, n46699, n46700,
         n46701, n46702, n46703, n46704, n46705, n46706, n46707, n46708,
         n46709, n46710, n46711, n46712, n46713, n46714, n46715, n46716,
         n46717, n46718, n46719, n46720, n46721, n46722, n46723, n46724,
         n46725, n46726, n46727, n46728, n46729, n46730, n46731, n46732,
         n46733, n46734, n46735, n46736, n46737, n46738, n46739, n46740,
         n46741, n46742, n46743, n46744, n46745, n46746, n46747, n46748,
         n46749, n46750, n46751, n46752, n46753, n46754, n46755, n46756,
         n46757, n46758, n46759, n46760, n46761, n46762, n46763, n46764,
         n46765, n46766, n46767, n46768, n46769, n46770, n46771, n46772,
         n46773, n46774, n46775, n46776, n46777, n46778, n46779, n46780,
         n46781, n46782, n46783, n46784, n46785, n46786, n46787, n46788,
         n46789, n46790, n46791, n46792, n46793, n46794, n46795, n46796,
         n46797, n46798, n46799, n46800, n46801, n46802, n46803, n46804,
         n46805, n46806, n46807, n46808, n46809, n46810, n46811, n46812,
         n46813, n46814, n46815, n46816, n46817, n46818, n46819, n46820,
         n46821, n46822, n46823, n46824, n46825, n46826, n46827, n46828,
         n46829, n46830, n46831, n46832, n46833, n46834, n46835, n46836,
         n46837, n46838, n46839, n46840, n46841, n46842, n46843, n46844,
         n46845, n46846, n46847, n46848, n46849, n46850, n46851, n46852,
         n46853, n46854, n46855, n46856, n46857, n46858, n46859, n46860,
         n46861, n46862, n46863, n46864, n46865, n46866, n46867, n46868,
         n46869, n46870, n46871, n46872, n46873, n46874, n46875, n46876,
         n46877, n46878, n46879, n46880, n46881, n46882, n46883, n46884,
         n46885, n46886, n46887, n46888, n46889, n46890, n46891, n46892,
         n46893, n46894, n46895, n46896, n46897, n46898, n46899, n46900,
         n46901, n46902, n46903, n46904, n46905, n46906, n46907, n46908,
         n46909, n46910, n46911, n46912, n46913, n46914, n46915, n46916,
         n46917, n46918, n46919, n46920, n46921, n46922, n46923, n46924,
         n46925, n46926, n46927, n46928, n46929, n46930, n46931, n46932,
         n46933, n46934, n46935, n46936, n46937, n46938, n46939, n46940,
         n46941, n46942, n46943, n46944, n46945, n46946, n46947, n46948,
         n46949, n46950, n46951, n46952, n46953, n46954, n46955, n46956,
         n46957, n46958, n46959, n46960, n46961, n46962, n46963, n46964,
         n46965, n46966, n46967, n46968, n46969, n46970, n46971, n46972,
         n46973, n46974, n46975, n46976, n46977, n46978, n46979, n46980,
         n46981, n46982, n46983, n46984, n46985, n46986, n46987, n46988,
         n46989, n46990, n46991, n46992, n46993, n46994, n46995, n46996,
         n46997, n46998, n46999, n47000, n47001, n47002, n47003, n47004,
         n47005, n47006, n47007, n47008, n47009, n47010, n47011, n47012,
         n47013, n47014, n47015, n47016, n47017, n47018, n47019, n47020,
         n47021, n47022, n47023, n47024, n47025, n47026, n47027, n47028,
         n47029, n47030, n47031, n47032, n47033, n47034, n47035, n47036,
         n47037, n47038, n47039, n47040, n47041, n47042, n47043, n47044,
         n47045, n47046, n47047, n47048, n47049, n47050, n47051, n47052,
         n47053, n47054, n47055, n47056, n47057, n47058, n47059, n47060,
         n47061, n47062, n47063, n47064, n47065, n47066, n47067, n47068,
         n47069, n47070, n47071, n47072, n47073, n47074, n47075, n47076,
         n47077, n47078, n47079, n47080, n47081, n47082, n47083, n47084,
         n47085, n47086, n47087, n47088, n47089, n47090, n47091, n47092,
         n47093, n47094, n47095, n47096, n47097, n47098, n47099, n47100,
         n47101, n47102, n47103, n47104, n47105, n47106, n47107, n47108,
         n47109, n47110, n47111, n47112, n47113, n47114, n47115, n47116,
         n47117, n47118, n47119, n47120, n47121, n47122, n47123, n47124,
         n47125, n47126, n47127, n47128, n47129, n47130, n47131, n47132,
         n47133, n47134, n47135, n47136, n47137, n47138, n47139, n47140,
         n47141, n47142, n47143, n47144, n47145, n47146, n47147, n47148,
         n47149, n47150, n47151, n47152, n47153, n47154, n47155, n47156,
         n47157, n47158, n47159, n47160, n47161, n47162, n47163, n47164,
         n47165, n47166, n47167, n47168, n47169, n47170, n47171, n47172,
         n47173, n47174, n47175, n47176, n47177, n47178, n47179, n47180,
         n47181, n47182, n47183, n47184, n47185, n47186, n47187, n47188,
         n47189, n47190, n47191, n47192, n47193, n47194, n47195, n47196,
         n47197, n47198, n47199, n47200, n47201, n47202, n47203, n47204,
         n47205, n47206, n47207, n47208, n47209, n47210, n47211, n47212,
         n47213, n47214, n47215, n47216, n47217, n47218, n47219, n47220,
         n47221, n47222, n47223, n47224, n47225, n47226, n47227, n47228,
         n47229, n47230, n47231, n47232, n47233, n47234, n47235, n47236,
         n47237, n47238, n47239, n47240, n47241, n47242, n47243, n47244,
         n47245, n47246, n47247, n47248, n47249, n47250, n47251, n47252,
         n47253, n47254, n47255, n47256, n47257, n47258, n47259, n47260,
         n47261, n47262, n47263, n47264, n47265, n47266, n47267, n47268,
         n47269, n47270, n47271, n47272, n47273, n47274, n47275, n47276,
         n47277, n47278, n47279, n47280, n47281, n47282, n47283, n47284,
         n47285, n47286, n47287, n47288, n47289, n47290, n47291, n47292,
         n47293, n47294, n47295, n47296, n47297, n47298, n47299, n47300,
         n47301, n47302, n47303, n47304, n47305, n47306, n47307, n47308,
         n47309, n47310, n47311, n47312, n47313, n47314, n47315, n47316,
         n47317, n47318, n47319, n47320, n47321, n47322, n47323, n47324,
         n47325, n47326, n47327, n47328, n47329, n47330, n47331, n47332,
         n47333, n47334, n47335, n47336, n47337, n47338, n47339, n47340,
         n47341, n47342, n47343, n47344, n47345, n47346, n47347, n47348,
         n47349, n47350, n47351, n47352, n47353, n47354, n47355, n47356,
         n47357, n47358, n47359, n47360, n47361, n47362, n47363, n47364,
         n47365, n47366, n47367, n47368, n47369, n47370, n47371, n47372,
         n47373, n47374, n47375, n47376, n47377, n47378, n47379, n47380,
         n47381, n47382, n47383, n47384, n47385, n47386, n47387, n47388,
         n47389, n47390, n47391, n47392, n47393, n47394, n47395, n47396,
         n47397, n47398, n47399, n47400, n47401, n47402, n47403, n47404,
         n47405, n47406, n47407, n47408, n47409, n47410, n47411, n47412,
         n47413, n47414, n47415, n47416, n47417, n47418, n47419, n47420,
         n47421, n47422, n47423, n47424, n47425, n47426, n47427, n47428,
         n47429, n47430, n47431, n47432, n47433, n47434, n47435, n47436,
         n47437, n47438, n47439, n47440, n47441, n47442, n47443, n47444,
         n47445, n47446, n47447, n47448, n47449, n47450, n47451, n47452,
         n47453, n47454, n47455, n47456, n47457, n47458, n47459, n47460,
         n47461, n47462, n47463, n47464, n47465, n47466, n47467, n47468,
         n47469, n47470, n47471, n47472, n47473, n47474, n47475, n47476,
         n47477, n47478, n47479, n47480, n47481, n47482, n47483, n47484,
         n47485, n47486, n47487, n47488, n47489, n47490, n47491, n47492,
         n47493, n47494, n47495, n47496, n47497, n47498, n47499, n47500,
         n47501, n47502, n47503, n47504, n47505, n47506, n47507, n47508,
         n47509, n47510, n47511, n47512, n47513, n47514, n47515, n47516,
         n47517, n47518, n47519, n47520, n47521, n47522, n47523, n47524,
         n47525, n47526, n47527, n47528, n47529, n47530, n47531, n47532,
         n47533, n47534, n47535, n47536, n47537, n47538, n47539, n47540,
         n47541, n47542, n47543, n47544, n47545, n47546, n47547, n47548,
         n47549, n47550, n47551, n47552, n47553, n47554, n47555, n47556,
         n47557, n47558, n47559, n47560, n47561, n47562, n47563, n47564,
         n47565, n47566, n47567, n47568, n47569, n47570, n47571, n47572,
         n47573, n47574, n47575, n47576, n47577, n47578, n47579, n47580,
         n47581, n47582, n47583, n47584, n47585, n47586, n47587, n47588,
         n47589, n47590, n47591, n47592, n47593, n47594, n47595, n47596,
         n47597, n47598, n47599, n47600, n47601, n47602, n47603, n47604,
         n47605, n47606, n47607, n47608, n47609, n47610, n47611, n47612,
         n47613, n47614, n47615, n47616, n47617, n47618, n47619, n47620,
         n47621, n47622, n47623, n47624, n47625, n47626, n47627, n47628,
         n47629, n47630, n47631, n47632, n47633, n47634, n47635, n47636,
         n47637, n47638, n47639, n47640, n47641, n47642, n47643, n47644,
         n47645, n47646, n47647, n47648, n47649, n47650, n47651, n47652,
         n47653, n47654, n47655, n47656, n47657, n47658, n47659, n47660,
         n47661, n47662, n47663, n47664, n47665, n47666, n47667, n47668,
         n47669, n47670, n47671, n47672, n47673, n47674, n47675, n47676,
         n47677, n47678, n47679, n47680, n47681, n47682, n47683, n47684,
         n47685, n47686, n47687, n47688, n47689, n47690, n47691, n47692,
         n47693, n47694, n47695, n47696, n47697, n47698, n47699, n47700,
         n47701, n47702, n47703, n47704, n47705, n47706, n47707, n47708,
         n47709, n47710, n47711, n47712, n47713, n47714, n47715, n47716,
         n47717, n47718, n47719, n47720, n47721, n47722, n47723, n47724,
         n47725, n47726, n47727, n47728, n47729, n47730, n47731, n47732,
         n47733, n47734, n47735, n47736, n47737, n47738, n47739, n47740,
         n47741, n47742, n47743, n47744, n47745, n47746, n47747, n47748,
         n47749, n47750, n47751, n47752, n47753, n47754, n47755, n47756,
         n47757, n47758, n47759, n47760, n47761, n47762, n47763, n47764,
         n47765, n47766, n47767, n47768, n47769, n47770, n47771, n47772,
         n47773, n47774, n47775, n47776, n47777, n47778, n47779, n47780,
         n47781, n47782, n47783, n47784, n47785, n47786, n47787, n47788,
         n47789, n47790, n47791, n47792, n47793, n47794, n47795, n47796,
         n47797, n47798, n47799, n47800, n47801, n47802, n47803, n47804,
         n47805, n47806, n47807, n47808, n47809, n47810, n47811, n47812,
         n47813, n47814, n47815, n47816, n47817, n47818, n47819, n47820,
         n47821, n47822, n47823, n47824, n47825, n47826, n47827, n47828,
         n47829, n47830, n47831, n47832, n47833, n47834, n47835, n47836,
         n47837, n47838, n47839, n47840, n47841, n47842, n47843, n47844,
         n47845, n47846, n47847, n47848, n47849, n47850, n47851, n47852,
         n47853, n47854, n47855, n47856, n47857, n47858, n47859, n47860,
         n47861, n47862, n47863, n47864, n47865, n47866, n47867, n47868,
         n47869, n47870, n47871, n47872, n47873, n47874, n47875, n47876,
         n47877, n47878, n47879, n47880, n47881, n47882, n47883, n47884,
         n47885, n47886, n47887, n47888, n47889, n47890, n47891, n47892,
         n47893, n47894, n47895, n47896, n47897, n47898, n47899, n47900,
         n47901, n47902, n47903, n47904, n47905, n47906, n47907, n47908,
         n47909, n47910, n47911, n47912, n47913, n47914, n47915, n47916,
         n47917, n47918, n47919, n47920, n47921, n47922, n47923, n47924,
         n47925, n47926, n47927, n47928, n47929, n47930, n47931, n47932,
         n47933, n47934, n47935, n47936, n47937, n47938, n47939, n47940,
         n47941, n47942, n47943, n47944, n47945, n47946, n47947, n47948,
         n47949, n47950, n47951, n47952, n47953, n47954, n47955, n47956,
         n47957, n47958, n47959, n47960, n47961, n47962, n47963, n47964,
         n47965, n47966, n47967, n47968, n47969, n47970, n47971, n47972,
         n47973, n47974, n47975, n47976, n47977, n47978, n47979, n47980,
         n47981, n47982, n47983, n47984, n47985, n47986, n47987, n47988,
         n47989, n47990, n47991, n47992, n47993, n47994, n47995, n47996,
         n47997, n47998, n47999, n48000, n48001, n48002, n48003, n48004,
         n48005, n48006, n48007, n48008, n48009, n48010, n48011, n48012,
         n48013, n48014, n48015, n48016, n48017, n48018, n48019, n48020,
         n48021, n48022, n48023, n48024, n48025, n48026, n48027, n48028,
         n48029, n48030, n48031, n48032, n48033, n48034, n48035, n48036,
         n48037, n48038, n48039, n48040, n48041, n48042, n48043, n48044,
         n48045, n48046, n48047, n48048, n48049, n48050, n48051, n48052,
         n48053, n48054, n48055, n48056, n48057, n48058, n48059, n48060,
         n48061, n48062, n48063, n48064, n48065, n48066, n48067, n48068,
         n48069, n48070, n48071, n48072, n48073, n48074, n48075, n48076,
         n48077, n48078, n48079, n48080, n48081, n48082, n48083, n48084,
         n48085, n48086, n48087, n48088, n48089, n48090, n48091, n48092,
         n48093, n48094, n48095, n48096, n48097, n48098, n48099, n48100,
         n48101, n48102, n48103, n48104, n48105, n48106, n48107, n48108,
         n48109, n48110, n48111, n48112, n48113, n48114, n48115, n48116,
         n48117, n48118, n48119, n48120, n48121, n48122, n48123, n48124,
         n48125, n48126, n48127, n48128, n48129, n48130, n48131, n48132,
         n48133, n48134, n48135, n48136, n48137, n48138, n48139, n48140,
         n48141, n48142, n48143, n48144, n48145, n48146, n48147, n48148,
         n48149, n48150, n48151, n48152, n48153, n48154, n48155, n48156,
         n48157, n48158, n48159, n48160, n48161, n48162, n48163, n48164,
         n48165, n48166, n48167, n48168, n48169, n48170, n48171, n48172,
         n48173, n48174, n48175, n48176, n48177, n48178, n48179, n48180,
         n48181, n48182, n48183, n48184, n48185, n48186, n48187, n48188,
         n48189, n48190, n48191, n48192, n48193, n48194, n48195, n48196,
         n48197, n48198, n48199, n48200, n48201, n48202, n48203, n48204,
         n48205, n48206, n48207, n48208, n48209, n48210, n48211, n48212,
         n48213, n48214, n48215, n48216, n48217, n48218, n48219, n48220,
         n48221, n48222, n48223, n48224, n48225, n48226, n48227, n48228,
         n48229, n48230, n48231, n48232, n48233, n48234, n48235, n48236,
         n48237, n48238, n48239, n48240, n48241, n48242, n48243, n48244,
         n48245, n48246, n48247, n48248, n48249, n48250, n48251, n48252,
         n48253, n48254, n48255, n48256, n48257, n48258, n48259, n48260,
         n48261, n48262, n48263, n48264, n48265, n48266, n48267, n48268,
         n48269, n48270, n48271, n48272, n48273, n48274, n48275, n48276,
         n48277, n48278, n48279, n48280, n48281, n48282, n48283, n48284,
         n48285, n48286, n48287, n48288, n48289, n48290, n48291, n48292,
         n48293, n48294, n48295, n48296, n48297, n48298, n48299, n48300,
         n48301, n48302, n48303, n48304, n48305, n48306, n48307, n48308,
         n48309, n48310, n48311, n48312, n48313, n48314, n48315, n48316,
         n48317, n48318, n48319, n48320, n48321, n48322, n48323, n48324,
         n48325, n48326, n48327, n48328, n48329, n48330, n48331, n48332,
         n48333, n48334, n48335, n48336, n48337, n48338, n48339, n48340,
         n48341, n48342, n48343, n48344, n48345, n48346, n48347, n48348,
         n48349, n48350, n48351, n48352, n48353, n48354, n48355, n48356,
         n48357, n48358, n48359, n48360, n48361, n48362, n48363, n48364,
         n48365, n48366, n48367, n48368, n48369, n48370, n48371, n48372,
         n48373, n48374, n48375, n48376, n48377, n48378, n48379, n48380,
         n48381, n48382, n48383, n48384, n48385, n48386, n48387, n48388,
         n48389, n48390, n48391, n48392, n48393, n48394, n48395, n48396,
         n48397, n48398, n48399, n48400, n48401, n48402, n48403, n48404,
         n48405, n48406, n48407, n48408, n48409, n48410, n48411, n48412,
         n48413, n48414, n48415, n48416, n48417, n48418, n48419, n48420,
         n48421, n48422, n48423, n48424, n48425, n48426, n48427, n48428,
         n48429, n48430, n48431, n48432, n48433, n48434, n48435, n48436,
         n48437, n48438, n48439, n48440, n48441, n48442, n48443, n48444,
         n48445, n48446, n48447, n48448, n48449, n48450, n48451, n48452,
         n48453, n48454, n48455, n48456, n48457, n48458, n48459, n48460,
         n48461, n48462, n48463, n48464, n48465, n48466, n48467, n48468,
         n48469, n48470, n48471, n48472, n48473, n48474, n48475, n48476,
         n48477, n48478, n48479, n48480, n48481, n48482, n48483, n48484,
         n48485, n48486, n48487, n48488, n48489, n48490, n48491, n48492,
         n48493, n48494, n48495, n48496, n48497, n48498, n48499, n48500,
         n48501, n48502, n48503, n48504, n48505, n48506, n48507, n48508,
         n48509, n48510, n48511, n48512, n48513, n48514, n48515, n48516,
         n48517, n48518, n48519, n48520, n48521, n48522, n48523, n48524,
         n48525, n48526, n48527, n48528, n48529, n48530, n48531, n48532,
         n48533, n48534, n48535, n48536, n48537, n48538, n48539, n48540,
         n48541, n48542, n48543, n48544, n48545, n48546, n48547, n48548,
         n48549, n48550, n48551, n48552, n48553, n48554, n48555, n48556,
         n48557, n48558, n48559, n48560, n48561, n48562, n48563, n48564,
         n48565, n48566, n48567, n48568, n48569, n48570, n48571, n48572,
         n48573, n48574, n48575, n48576, n48577, n48578, n48579, n48580,
         n48581, n48582, n48583, n48584, n48585, n48586, n48587, n48588,
         n48589, n48590, n48591, n48592, n48593, n48594, n48595, n48596,
         n48597, n48598, n48599, n48600, n48601, n48602, n48603, n48604,
         n48605, n48606, n48607, n48608, n48609, n48610, n48611, n48612,
         n48613, n48614, n48615, n48616, n48617, n48618, n48619, n48620,
         n48621, n48622, n48623, n48624, n48625, n48626, n48627, n48628,
         n48629, n48630, n48631, n48632, n48633, n48634, n48635, n48636,
         n48637, n48638, n48639, n48640, n48641, n48642, n48643, n48644,
         n48645, n48646, n48647, n48648, n48649, n48650, n48651, n48652,
         n48653, n48654, n48655, n48656, n48657, n48658, n48659, n48660,
         n48661, n48662, n48663, n48664, n48665, n48666, n48667, n48668,
         n48669, n48670, n48671, n48672, n48673, n48674, n48675, n48676,
         n48677, n48678, n48679, n48680, n48681, n48682, n48683, n48684,
         n48685, n48686, n48687, n48688, n48689, n48690, n48691, n48692,
         n48693, n48694, n48695, n48696, n48697, n48698, n48699, n48700,
         n48701, n48702, n48703, n48704, n48705, n48706, n48707, n48708,
         n48709, n48710, n48711, n48712, n48713, n48714, n48715, n48716,
         n48717, n48718, n48719, n48720, n48721, n48722, n48723, n48724,
         n48725, n48726, n48727, n48728, n48729, n48730, n48731, n48732,
         n48733, n48734, n48735, n48736, n48737, n48738, n48739, n48740,
         n48741, n48742, n48743, n48744, n48745, n48746, n48747, n48748,
         n48749, n48750, n48751, n48752, n48753, n48754, n48755, n48756,
         n48757, n48758, n48759, n48760, n48761, n48762, n48763, n48764,
         n48765, n48766, n48767, n48768, n48769, n48770, n48771, n48772,
         n48773, n48774, n48775, n48776, n48777, n48778, n48779, n48780,
         n48781, n48782, n48783, n48784, n48785, n48786, n48787, n48788,
         n48789, n48790, n48791, n48792, n48793, n48794, n48795, n48796,
         n48797, n48798, n48799, n48800, n48801, n48802, n48803, n48804,
         n48805, n48806, n48807, n48808, n48809, n48810, n48811, n48812,
         n48813, n48814, n48815, n48816, n48817, n48818, n48819, n48820,
         n48821, n48822, n48823, n48824, n48825, n48826, n48827, n48828,
         n48829, n48830, n48831, n48832, n48833, n48834, n48835, n48836,
         n48837, n48838, n48839, n48840, n48841, n48842, n48843, n48844,
         n48845, n48846, n48847, n48848, n48849, n48850, n48851, n48852,
         n48853, n48854, n48855, n48856, n48857, n48858, n48859, n48860,
         n48861, n48862, n48863, n48864, n48865, n48866, n48867, n48868,
         n48869, n48870, n48871, n48872, n48873, n48874, n48875, n48876,
         n48877, n48878, n48879, n48880, n48881, n48882, n48883, n48884,
         n48885, n48886, n48887, n48888, n48889, n48890, n48891, n48892,
         n48893, n48894, n48895, n48896, n48897, n48898, n48899, n48900,
         n48901, n48902, n48903, n48904, n48905, n48906, n48907, n48908,
         n48909, n48910, n48911, n48912, n48913, n48914, n48915, n48916,
         n48917, n48918, n48919, n48920, n48921, n48922, n48923, n48924,
         n48925, n48926, n48927, n48928, n48929, n48930, n48931, n48932,
         n48933, n48934, n48935, n48936, n48937, n48938, n48939, n48940,
         n48941, n48942, n48943, n48944, n48945, n48946, n48947, n48948,
         n48949, n48950, n48951, n48952, n48953, n48954, n48955, n48956,
         n48957, n48958, n48959, n48960, n48961, n48962, n48963, n48964,
         n48965, n48966, n48967, n48968, n48969, n48970, n48971, n48972,
         n48973, n48974, n48975, n48976, n48977, n48978, n48979, n48980,
         n48981, n48982, n48983, n48984, n48985, n48986, n48987, n48988,
         n48989, n48990, n48991, n48992, n48993, n48994, n48995, n48996,
         n48997, n48998, n48999, n49000, n49001, n49002, n49003, n49004,
         n49005, n49006, n49007, n49008, n49009, n49010, n49011, n49012,
         n49013, n49014, n49015, n49016, n49017, n49018, n49019, n49020,
         n49021, n49022, n49023, n49024, n49025, n49026, n49027, n49028,
         n49029, n49030, n49031, n49032, n49033, n49034, n49035, n49036,
         n49037, n49038, n49039, n49040, n49041, n49042, n49043, n49044,
         n49045, n49046, n49047, n49048, n49049, n49050, n49051, n49052,
         n49053, n49054, n49055, n49056, n49057, n49058, n49059, n49060,
         n49061, n49062, n49063, n49064, n49065, n49066, n49067, n49068,
         n49069, n49070, n49071, n49072, n49073, n49074, n49075, n49076,
         n49077, n49078, n49079, n49080, n49081, n49082, n49083, n49084,
         n49085, n49086, n49087, n49088, n49089, n49090, n49091, n49092,
         n49093, n49094, n49095, n49096, n49097, n49098, n49099, n49100,
         n49101, n49102, n49103, n49104, n49105, n49106, n49107, n49108,
         n49109, n49110, n49111, n49112, n49113, n49114, n49115, n49116,
         n49117, n49118, n49119, n49120, n49121, n49122, n49123, n49124,
         n49125, n49126, n49127, n49128, n49129, n49130, n49131, n49132,
         n49133, n49134, n49135, n49136, n49137, n49138, n49139, n49140,
         n49141, n49142, n49143, n49144, n49145, n49146, n49147, n49148,
         n49149, n49150, n49151, n49152, n49153, n49154, n49155, n49156,
         n49157, n49158, n49159, n49160, n49161, n49162, n49163, n49164,
         n49165, n49166, n49167, n49168, n49169, n49170, n49171, n49172,
         n49173, n49174, n49175, n49176, n49177, n49178, n49179, n49180,
         n49181, n49182, n49183, n49184, n49185, n49186, n49187, n49188,
         n49189, n49190, n49191, n49192, n49193, n49194, n49195, n49196,
         n49197, n49198, n49199, n49200, n49201, n49202, n49203, n49204,
         n49205, n49206, n49207, n49208, n49209, n49210, n49211, n49212,
         n49213, n49214, n49215, n49216, n49217, n49218, n49219, n49220,
         n49221, n49222, n49223, n49224, n49225, n49226, n49227, n49228,
         n49229, n49230, n49231, n49232, n49233, n49234, n49235, n49236,
         n49237, n49238, n49239, n49240, n49241, n49242, n49243, n49244,
         n49245, n49246, n49247, n49248, n49249, n49250, n49251, n49252,
         n49253, n49254, n49255, n49256, n49257, n49258, n49259, n49260,
         n49261, n49262, n49263, n49264, n49265, n49266, n49267, n49268,
         n49269, n49270, n49271, n49272, n49273, n49274, n49275, n49276,
         n49277, n49278, n49279, n49280, n49281, n49282, n49283, n49284,
         n49285, n49286, n49287, n49288, n49289, n49290, n49291, n49292,
         n49293, n49294, n49295, n49296, n49297, n49298, n49299, n49300,
         n49301, n49302, n49303, n49304, n49305, n49306, n49307, n49308,
         n49309, n49310, n49311, n49312, n49313, n49314, n49315, n49316,
         n49317, n49318, n49319, n49320, n49321, n49322, n49323, n49324,
         n49325, n49326, n49327, n49328, n49329, n49330, n49331, n49332,
         n49333, n49334, n49335, n49336, n49337, n49338, n49339, n49340,
         n49341, n49342, n49343, n49344, n49345, n49346, n49347, n49348,
         n49349, n49350, n49351, n49352, n49353, n49354, n49355, n49356,
         n49357, n49358, n49359, n49360, n49361, n49362, n49363, n49364,
         n49365, n49366, n49367, n49368, n49369, n49370, n49371, n49372,
         n49373, n49374, n49375, n49376, n49377, n49378, n49379, n49380,
         n49381, n49382, n49383, n49384, n49385, n49386, n49387, n49388,
         n49389, n49390, n49391, n49392, n49393, n49394, n49395, n49396,
         n49397, n49398, n49399, n49400, n49401, n49402, n49403, n49404,
         n49405, n49406, n49407, n49408, n49409, n49410, n49411, n49412,
         n49413, n49414, n49415, n49416, n49417, n49418, n49419, n49420,
         n49421, n49422, n49423, n49424, n49425, n49426, n49427, n49428,
         n49429, n49430, n49431, n49432, n49433, n49434, n49435, n49436,
         n49437, n49438, n49439, n49440, n49441, n49442, n49443, n49444,
         n49445, n49446, n49447, n49448, n49449, n49450, n49451, n49452,
         n49453, n49454, n49455, n49456, n49457, n49458, n49459, n49460,
         n49461, n49462, n49463, n49464, n49465, n49466, n49467, n49468,
         n49469, n49470, n49471, n49472, n49473, n49474, n49475, n49476,
         n49477, n49478, n49479, n49480, n49481, n49482, n49483, n49484,
         n49485, n49486, n49487, n49488, n49489, n49490, n49491, n49492,
         n49493, n49494, n49495, n49496, n49497, n49498, n49499, n49500,
         n49501, n49502, n49503, n49504, n49505, n49506, n49507, n49508,
         n49509, n49510, n49511, n49512, n49513, n49514, n49515, n49516,
         n49517, n49518, n49519, n49520, n49521, n49522, n49523, n49524,
         n49525, n49526, n49527, n49528, n49529, n49530, n49531, n49532,
         n49533, n49534, n49535, n49536, n49537, n49538, n49539, n49540,
         n49541, n49542, n49543, n49544, n49545, n49546, n49547, n49548,
         n49549, n49550, n49551, n49552, n49553, n49554, n49555, n49556,
         n49557, n49558, n49559, n49560, n49561, n49562, n49563, n49564,
         n49565, n49566, n49567, n49568, n49569, n49570, n49571, n49572,
         n49573, n49574, n49575, n49576, n49577, n49578, n49579, n49580,
         n49581, n49582, n49583, n49584, n49585, n49586, n49587, n49588,
         n49589, n49590, n49591, n49592, n49593, n49594, n49595, n49596,
         n49597, n49598, n49599, n49600, n49601, n49602, n49603, n49604,
         n49605, n49606, n49607, n49608, n49609, n49610, n49611, n49612,
         n49613, n49614, n49615, n49616, n49617, n49618, n49619, n49620,
         n49621, n49622, n49623, n49624, n49625, n49626, n49627, n49628,
         n49629, n49630, n49631, n49632, n49633, n49634, n49635, n49636,
         n49637, n49638, n49639, n49640, n49641, n49642, n49643, n49644,
         n49645, n49646, n49647, n49648, n49649, n49650, n49651, n49652,
         n49653, n49654, n49655, n49656, n49657, n49658, n49659, n49660,
         n49661, n49662, n49663, n49664, n49665, n49666, n49667, n49668,
         n49669, n49670, n49671, n49672, n49673, n49674, n49675, n49676,
         n49677, n49678, n49679, n49680, n49681, n49682, n49683, n49684,
         n49685, n49686, n49687, n49688, n49689, n49690, n49691, n49692,
         n49693, n49694, n49695, n49696, n49697, n49698, n49699, n49700,
         n49701, n49702, n49703, n49704, n49705, n49706, n49707, n49708,
         n49709, n49710, n49711, n49712, n49713, n49714, n49715, n49716,
         n49717, n49718, n49719, n49720, n49721, n49722, n49723, n49724,
         n49725, n49726, n49727, n49728, n49729, n49730, n49731, n49732,
         n49733, n49734, n49735, n49736, n49737, n49738, n49739, n49740,
         n49741, n49742, n49743, n49744, n49745, n49746, n49747, n49748,
         n49749, n49750, n49751, n49752, n49753, n49754, n49755, n49756,
         n49757, n49758, n49759, n49760, n49761, n49762, n49763, n49764,
         n49765, n49766, n49767, n49768, n49769, n49770, n49771, n49772,
         n49773, n49774, n49775, n49776, n49777, n49778, n49779, n49780,
         n49781, n49782, n49783, n49784, n49785, n49786, n49787, n49788,
         n49789, n49790, n49791, n49792, n49793, n49794, n49795, n49796,
         n49797, n49798, n49799, n49800, n49801, n49802, n49803, n49804,
         n49805, n49806, n49807, n49808, n49809, n49810, n49811, n49812,
         n49813, n49814, n49815, n49816, n49817, n49818, n49819, n49820,
         n49821, n49822, n49823, n49824, n49825, n49826, n49827, n49828,
         n49829, n49830, n49831, n49832, n49833, n49834, n49835, n49836,
         n49837, n49838, n49839, n49840, n49841, n49842, n49843, n49844,
         n49845, n49846, n49847, n49848, n49849, n49850, n49851, n49852,
         n49853, n49854, n49855, n49856, n49857, n49858, n49859, n49860,
         n49861, n49862, n49863, n49864, n49865, n49866, n49867, n49868,
         n49869, n49870, n49871, n49872, n49873, n49874, n49875, n49876,
         n49877, n49878, n49879, n49880, n49881, n49882, n49883, n49884,
         n49885, n49886, n49887, n49888, n49889, n49890, n49891, n49892,
         n49893, n49894, n49895, n49896, n49897, n49898, n49899, n49900,
         n49901, n49902, n49903, n49904, n49905, n49906, n49907, n49908,
         n49909, n49910, n49911, n49912, n49913, n49914, n49915, n49916,
         n49917, n49918, n49919, n49920, n49921, n49922, n49923, n49924,
         n49925, n49926, n49927, n49928, n49929, n49930, n49931, n49932,
         n49933, n49934, n49935, n49936, n49937, n49938, n49939, n49940,
         n49941, n49942, n49943, n49944, n49945, n49946, n49947, n49948,
         n49949, n49950, n49951, n49952, n49953, n49954, n49955, n49956,
         n49957, n49958, n49959, n49960, n49961, n49962, n49963, n49964,
         n49965, n49966, n49967, n49968, n49969, n49970, n49971, n49972,
         n49973, n49974, n49975, n49976, n49977, n49978, n49979, n49980,
         n49981, n49982, n49983, n49984, n49985, n49986, n49987, n49988,
         n49989, n49990, n49991, n49992, n49993, n49994, n49995, n49996,
         n49997, n49998, n49999, n50000, n50001, n50002, n50003, n50004,
         n50005, n50006, n50007, n50008, n50009, n50010, n50011, n50012,
         n50013, n50014, n50015, n50016, n50017, n50018, n50019, n50020,
         n50021, n50022, n50023, n50024, n50025, n50026, n50027, n50028,
         n50029, n50030, n50031, n50032, n50033, n50034, n50035, n50036,
         n50037, n50038, n50039, n50040, n50041, n50042, n50043, n50044,
         n50045, n50046, n50047, n50048, n50049, n50050, n50051, n50052,
         n50053, n50054, n50055, n50056, n50057, n50058, n50059, n50060,
         n50061, n50062, n50063, n50064, n50065, n50066, n50067, n50068,
         n50069, n50070, n50071, n50072, n50073, n50074, n50075, n50076,
         n50077, n50078, n50079, n50080, n50081, n50082, n50083, n50084,
         n50085, n50086, n50087, n50088, n50089, n50090, n50091, n50092,
         n50093, n50094, n50095, n50096, n50097, n50098, n50099, n50100,
         n50101, n50102, n50103, n50104, n50105, n50106, n50107, n50108,
         n50109, n50110, n50111, n50112, n50113, n50114, n50115, n50116,
         n50117, n50118, n50119, n50120, n50121, n50122, n50123, n50124,
         n50125, n50126, n50127, n50128, n50129, n50130, n50131, n50132,
         n50133, n50134, n50135, n50136, n50137, n50138, n50139, n50140,
         n50141, n50142, n50143, n50144, n50145, n50146, n50147, n50148,
         n50149, n50150, n50151, n50152, n50153, n50154, n50155, n50156,
         n50157, n50158, n50159, n50160, n50161, n50162, n50163, n50164,
         n50165, n50166, n50167, n50168, n50169, n50170, n50171, n50172,
         n50173, n50174, n50175, n50176, n50177, n50178, n50179, n50180,
         n50181, n50182, n50183, n50184, n50185, n50186, n50187, n50188,
         n50189, n50190, n50191, n50192, n50193, n50194, n50195, n50196,
         n50197, n50198, n50199, n50200, n50201, n50202, n50203, n50204,
         n50205, n50206, n50207, n50208, n50209, n50210, n50211, n50212,
         n50213, n50214, n50215, n50216, n50217, n50218, n50219, n50220,
         n50221, n50222, n50223, n50224, n50225, n50226, n50227, n50228,
         n50229, n50230, n50231, n50232, n50233, n50234, n50235, n50236,
         n50237, n50238, n50239, n50240, n50241, n50242, n50243, n50244,
         n50245, n50246, n50247, n50248, n50249, n50250, n50251, n50252,
         n50253, n50254, n50255, n50256, n50257, n50258, n50259, n50260,
         n50261, n50262, n50263, n50264, n50265, n50266, n50267, n50268,
         n50269, n50270, n50271, n50272, n50273, n50274, n50275, n50276,
         n50277, n50278, n50279, n50280, n50281, n50282, n50283, n50284,
         n50285, n50286, n50287, n50288, n50289, n50290, n50291, n50292,
         n50293, n50294, n50295, n50296, n50297, n50298, n50299, n50300,
         n50301, n50302, n50303, n50304, n50305, n50306, n50307, n50308,
         n50309, n50310, n50311, n50312, n50313, n50314, n50315, n50316,
         n50317, n50318, n50319, n50320, n50321, n50322, n50323, n50324,
         n50325, n50326, n50327, n50328, n50329, n50330, n50331, n50332,
         n50333, n50334, n50335, n50336, n50337, n50338, n50339, n50340,
         n50341, n50342, n50343, n50344, n50345, n50346, n50347, n50348,
         n50349, n50350, n50351, n50352, n50353, n50354, n50355, n50356,
         n50357, n50358, n50359, n50360, n50361, n50362, n50363, n50364,
         n50365, n50366, n50367, n50368, n50369, n50370, n50371, n50372,
         n50373, n50374, n50375, n50376, n50377, n50378, n50379, n50380,
         n50381, n50382, n50383, n50384, n50385, n50386, n50387, n50388,
         n50389, n50390, n50391, n50392, n50393, n50394, n50395, n50396,
         n50397, n50398, n50399, n50400, n50401, n50402, n50403, n50404,
         n50405, n50406, n50407, n50408, n50409, n50410, n50411, n50412,
         n50413, n50414, n50415, n50416, n50417, n50418, n50419, n50420,
         n50421, n50422, n50423, n50424, n50425, n50426, n50427, n50428,
         n50429, n50430, n50431, n50432, n50433, n50434, n50435, n50436,
         n50437, n50438, n50439, n50440, n50441, n50442, n50443, n50444,
         n50445, n50446, n50447, n50448, n50449, n50450, n50451, n50452,
         n50453, n50454, n50455, n50456, n50457, n50458, n50459, n50460,
         n50461, n50462, n50463, n50464, n50465, n50466, n50467, n50468,
         n50469, n50470, n50471, n50472, n50473, n50474, n50475, n50476,
         n50477, n50478, n50479, n50480, n50481, n50482, n50483, n50484,
         n50485, n50486, n50487, n50488, n50489, n50490, n50491, n50492,
         n50493, n50494, n50495, n50496, n50497, n50498, n50499, n50500,
         n50501, n50502, n50503, n50504, n50505, n50506, n50507, n50508,
         n50509, n50510, n50511, n50512, n50513, n50514, n50515, n50516,
         n50517, n50518, n50519, n50520, n50521, n50522, n50523, n50524,
         n50525, n50526, n50527, n50528, n50529, n50530, n50531, n50532,
         n50533, n50534, n50535, n50536, n50537, n50538, n50539, n50540,
         n50541, n50542, n50543, n50544, n50545, n50546, n50547, n50548,
         n50549, n50550, n50551, n50552, n50553, n50554, n50555, n50556,
         n50557, n50558, n50559, n50560, n50561, n50562, n50563, n50564,
         n50565, n50566, n50567, n50568, n50569, n50570, n50571, n50572,
         n50573, n50574, n50575, n50576, n50577, n50578, n50579, n50580,
         n50581, n50582, n50583, n50584, n50585, n50586, n50587, n50588,
         n50589, n50590, n50591, n50592, n50593, n50594, n50595, n50596,
         n50597, n50598, n50599, n50600, n50601, n50602, n50603, n50604,
         n50605, n50606, n50607, n50608, n50609, n50610, n50611, n50612,
         n50613, n50614, n50615, n50616, n50617, n50618, n50619, n50620,
         n50621, n50622, n50623, n50624, n50625, n50626, n50627, n50628,
         n50629, n50630, n50631, n50632, n50633, n50634, n50635, n50636,
         n50637, n50638, n50639, n50640, n50641, n50642, n50643, n50644,
         n50645, n50646, n50647, n50648, n50649, n50650, n50651, n50652,
         n50653, n50654, n50655, n50656, n50657, n50658, n50659, n50660,
         n50661, n50662, n50663, n50664, n50665, n50666, n50667, n50668,
         n50669, n50670, n50671, n50672, n50673, n50674, n50675, n50676,
         n50677, n50678, n50679, n50680, n50681, n50682, n50683, n50684,
         n50685, n50686, n50687, n50688, n50689, n50690, n50691, n50692,
         n50693, n50694, n50695, n50696, n50697, n50698, n50699, n50700,
         n50701, n50702, n50703, n50704, n50705, n50706, n50707, n50708,
         n50709, n50710, n50711, n50712, n50713, n50714, n50715, n50716,
         n50717, n50718, n50719, n50720, n50721, n50722, n50723, n50724,
         n50725, n50726, n50727, n50728, n50729, n50730, n50731, n50732,
         n50733, n50734, n50735, n50736, n50737, n50738, n50739, n50740,
         n50741, n50742, n50743, n50744, n50745, n50746, n50747, n50748,
         n50749, n50750, n50751, n50752, n50753, n50754, n50755, n50756,
         n50757, n50758, n50759, n50760, n50761, n50762, n50763, n50764,
         n50765, n50766, n50767, n50768, n50769, n50770, n50771, n50772,
         n50773, n50774, n50775, n50776, n50777, n50778, n50779, n50780,
         n50781, n50782, n50783, n50784, n50785, n50786, n50787, n50788,
         n50789, n50790, n50791, n50792, n50793, n50794, n50795, n50796,
         n50797, n50798, n50799, n50800, n50801, n50802, n50803, n50804,
         n50805, n50806, n50807, n50808, n50809, n50810, n50811, n50812,
         n50813, n50814, n50815, n50816, n50817, n50818, n50819, n50820,
         n50821, n50822, n50823, n50824, n50825, n50826, n50827, n50828,
         n50829, n50830, n50831, n50832, n50833, n50834, n50835, n50836,
         n50837, n50838, n50839, n50840, n50841, n50842, n50843, n50844,
         n50845, n50846, n50847, n50848, n50849, n50850, n50851, n50852,
         n50853, n50854, n50855, n50856, n50857, n50858, n50859, n50860,
         n50861, n50862, n50863, n50864, n50865, n50866, n50867, n50868,
         n50869, n50870, n50871, n50872, n50873, n50874, n50875, n50876,
         n50877, n50878, n50879, n50880, n50881, n50882, n50883, n50884,
         n50885, n50886, n50887, n50888, n50889, n50890, n50891, n50892,
         n50893, n50894, n50895, n50896, n50897, n50898, n50899, n50900,
         n50901, n50902, n50903, n50904, n50905, n50906, n50907, n50908,
         n50909, n50910, n50911, n50912, n50913, n50914, n50915, n50916,
         n50917, n50918, n50919, n50920, n50921, n50922, n50923, n50924,
         n50925, n50926, n50927, n50928, n50929, n50930, n50931, n50932,
         n50933, n50934, n50935, n50936, n50937, n50938, n50939, n50940,
         n50941, n50942, n50943, n50944, n50945, n50946, n50947, n50948,
         n50949, n50950, n50951, n50952, n50953, n50954, n50955, n50956,
         n50957, n50958, n50959, n50960, n50961, n50962, n50963, n50964,
         n50965, n50966, n50967, n50968, n50969, n50970, n50971, n50972,
         n50973, n50974, n50975, n50976, n50977, n50978, n50979, n50980,
         n50981, n50982, n50983, n50984, n50985, n50986, n50987, n50988,
         n50989, n50990, n50991, n50992, n50993, n50994, n50995, n50996,
         n50997, n50998, n50999, n51000, n51001, n51002, n51003, n51004,
         n51005, n51006, n51007, n51008, n51009, n51010, n51011, n51012,
         n51013, n51014, n51015, n51016, n51017, n51018, n51019, n51020,
         n51021, n51022, n51023, n51024, n51025, n51026, n51027, n51028,
         n51029, n51030, n51031, n51032, n51033, n51034, n51035, n51036,
         n51037, n51038, n51039, n51040, n51041, n51042, n51043, n51044,
         n51045, n51046, n51047, n51048, n51049, n51050, n51051, n51052,
         n51053, n51054, n51055, n51056, n51057, n51058, n51059, n51060,
         n51061, n51062, n51063, n51064, n51065, n51066, n51067, n51068,
         n51069, n51070, n51071, n51072, n51073, n51074, n51075, n51076,
         n51077, n51078, n51079, n51080, n51081, n51082, n51083, n51084,
         n51085, n51086, n51087, n51088, n51089, n51090, n51091, n51092,
         n51093, n51094, n51095, n51096, n51097, n51098, n51099, n51100,
         n51101, n51102, n51103, n51104, n51105, n51106, n51107, n51108,
         n51109, n51110, n51111, n51112, n51113, n51114, n51115, n51116,
         n51117, n51118, n51119, n51120, n51121, n51122, n51123, n51124,
         n51125, n51126, n51127, n51128, n51129, n51130, n51131, n51132,
         n51133, n51134, n51135, n51136, n51137, n51138, n51139, n51140,
         n51141, n51142, n51143, n51144, n51145, n51146, n51147, n51148,
         n51149, n51150, n51151, n51152, n51153, n51154, n51155, n51156,
         n51157, n51158, n51159, n51160, n51161, n51162, n51163, n51164,
         n51165, n51166, n51167, n51168, n51169, n51170, n51171, n51172,
         n51173, n51174, n51175, n51176, n51177, n51178, n51179, n51180,
         n51181, n51182, n51183, n51184, n51185, n51186, n51187, n51188,
         n51189, n51190, n51191, n51192, n51193, n51194, n51195, n51196,
         n51197, n51198, n51199, n51200, n51201, n51202, n51203, n51204,
         n51205, n51206, n51207, n51208, n51209, n51210, n51211, n51212,
         n51213, n51214, n51215, n51216, n51217, n51218, n51219, n51220,
         n51221, n51222, n51223, n51224, n51225, n51226, n51227, n51228,
         n51229, n51230, n51231, n51232, n51233, n51234, n51235, n51236,
         n51237, n51238, n51239, n51240, n51241, n51242, n51243, n51244,
         n51245, n51246, n51247, n51248, n51249, n51250, n51251, n51252,
         n51253, n51254, n51255, n51256, n51257, n51258, n51259, n51260,
         n51261, n51262, n51263, n51264, n51265, n51266, n51267, n51268,
         n51269, n51270, n51271, n51272, n51273, n51274, n51275, n51276,
         n51277, n51278, n51279, n51280, n51281, n51282, n51283, n51284,
         n51285, n51286, n51287, n51288, n51289, n51290, n51291, n51292,
         n51293, n51294, n51295, n51296, n51297, n51298, n51299, n51300,
         n51301, n51302, n51303, n51304, n51305, n51306, n51307, n51308,
         n51309, n51310, n51311, n51312, n51313, n51314, n51315, n51316,
         n51317, n51318, n51319, n51320, n51321, n51322, n51323, n51324,
         n51325, n51326, n51327, n51328, n51329, n51330, n51331, n51332,
         n51333, n51334, n51335, n51336, n51337, n51338, n51339, n51340,
         n51341, n51342, n51343, n51344, n51345, n51346, n51347, n51348,
         n51349, n51350, n51351, n51352, n51353, n51354, n51355, n51356,
         n51357, n51358, n51359, n51360, n51361, n51362, n51363, n51364,
         n51365, n51366, n51367, n51368, n51369, n51370, n51371, n51372,
         n51373, n51374, n51375, n51376, n51377, n51378, n51379, n51380,
         n51381, n51382, n51383, n51384, n51385, n51386, n51387, n51388,
         n51389, n51390, n51391, n51392, n51393, n51394, n51395, n51396,
         n51397, n51398, n51399, n51400, n51401, n51402, n51403, n51404,
         n51405, n51406, n51407, n51408, n51409, n51410, n51411, n51412,
         n51413, n51414, n51415, n51416, n51417, n51418, n51419, n51420,
         n51421, n51422, n51423, n51424, n51425, n51426, n51427, n51428,
         n51429, n51430, n51431, n51432, n51433, n51434, n51435, n51436,
         n51437, n51438, n51439, n51440, n51441, n51442, n51443, n51444,
         n51445, n51446, n51447, n51448, n51449, n51450, n51451, n51452,
         n51453, n51454, n51455, n51456, n51457, n51458, n51459, n51460,
         n51461, n51462, n51463, n51464, n51465, n51466, n51467, n51468,
         n51469, n51470, n51471, n51472, n51473, n51474, n51475, n51476,
         n51477, n51478, n51479, n51480, n51481, n51482, n51483, n51484,
         n51485, n51486, n51487, n51488, n51489, n51490, n51491, n51492,
         n51493, n51494, n51495, n51496, n51497, n51498, n51499, n51500,
         n51501, n51502, n51503, n51504, n51505, n51506, n51507, n51508,
         n51509, n51510, n51511, n51512, n51513, n51514, n51515, n51516,
         n51517, n51518, n51519, n51520, n51521, n51522, n51523, n51524,
         n51525, n51526, n51527, n51528, n51529, n51530, n51531, n51532,
         n51533, n51534, n51535, n51536, n51537, n51538, n51539, n51540,
         n51541, n51542, n51543, n51544, n51545, n51546, n51547, n51548,
         n51549, n51550, n51551, n51552, n51553, n51554, n51555, n51556,
         n51557, n51558, n51559, n51560, n51561, n51562, n51563, n51564,
         n51565, n51566, n51567, n51568, n51569, n51570, n51571, n51572,
         n51573, n51574, n51575, n51576, n51577, n51578, n51579, n51580,
         n51581, n51582, n51583, n51584, n51585, n51586, n51587, n51588,
         n51589, n51590, n51591, n51592, n51593, n51594, n51595, n51596,
         n51597, n51598, n51599, n51600, n51601, n51602, n51603, n51604,
         n51605, n51606, n51607, n51608, n51609, n51610, n51611, n51612,
         n51613, n51614, n51615, n51616, n51617, n51618, n51619, n51620,
         n51621, n51622, n51623, n51624, n51625, n51626, n51627, n51628,
         n51629, n51630, n51631, n51632, n51633, n51634, n51635, n51636,
         n51637, n51638, n51639, n51640, n51641, n51642, n51643, n51644,
         n51645, n51646, n51647, n51648, n51649, n51650, n51651, n51652,
         n51653, n51654, n51655, n51656, n51657, n51658, n51659, n51660,
         n51661, n51662, n51663, n51664, n51665, n51666, n51667, n51668,
         n51669, n51670, n51671, n51672, n51673, n51674, n51675, n51676,
         n51677, n51678, n51679, n51680, n51681, n51682, n51683, n51684,
         n51685, n51686, n51687, n51688, n51689, n51690, n51691, n51692,
         n51693, n51694, n51695, n51696, n51697, n51698, n51699, n51700,
         n51701, n51702, n51703, n51704, n51705, n51706, n51707, n51708,
         n51709, n51710, n51711, n51712, n51713, n51714, n51715, n51716,
         n51717, n51718, n51719, n51720, n51721, n51722, n51723, n51724,
         n51725, n51726, n51727, n51728, n51729, n51730, n51731, n51732,
         n51733, n51734, n51735, n51736, n51737, n51738, n51739, n51740,
         n51741, n51742, n51743, n51744, n51745, n51746, n51747, n51748,
         n51749, n51750, n51751, n51752, n51753, n51754, n51755, n51756,
         n51757, n51758, n51759, n51760, n51761, n51762, n51763, n51764,
         n51765, n51766, n51767, n51768, n51769, n51770, n51771, n51772,
         n51773, n51774, n51775, n51776, n51777, n51778, n51779, n51780,
         n51781, n51782, n51783, n51784, n51785, n51786, n51787, n51788,
         n51789, n51790, n51791, n51792, n51793, n51794, n51795, n51796,
         n51797, n51798, n51799, n51800, n51801, n51802, n51803, n51804,
         n51805, n51806, n51807, n51808, n51809, n51810, n51811, n51812,
         n51813, n51814, n51815, n51816, n51817, n51818, n51819, n51820,
         n51821, n51822, n51823, n51824, n51825, n51826, n51827, n51828,
         n51829, n51830, n51831, n51832, n51833, n51834, n51835, n51836,
         n51837, n51838, n51839, n51840, n51841, n51842, n51843, n51844,
         n51845, n51846, n51847, n51848, n51849, n51850, n51851, n51852,
         n51853, n51854, n51855, n51856, n51857, n51858, n51859, n51860,
         n51861, n51862, n51863, n51864, n51865, n51866, n51867, n51868,
         n51869, n51870, n51871, n51872, n51873, n51874, n51875, n51876,
         n51877, n51878, n51879, n51880, n51881, n51882, n51883, n51884,
         n51885, n51886, n51887, n51888, n51889, n51890, n51891, n51892,
         n51893, n51894, n51895, n51896, n51897, n51898, n51899, n51900,
         n51901, n51902, n51903, n51904, n51905, n51906, n51907, n51908,
         n51909, n51910, n51911, n51912, n51913, n51914, n51915, n51916,
         n51917, n51918, n51919, n51920, n51921, n51922, n51923, n51924,
         n51925, n51926, n51927, n51928, n51929, n51930, n51931, n51932,
         n51933, n51934, n51935, n51936, n51937, n51938, n51939, n51940,
         n51941, n51942, n51943, n51944, n51945, n51946, n51947, n51948,
         n51949, n51950, n51951, n51952, n51953, n51954, n51955, n51956,
         n51957, n51958, n51959, n51960, n51961, n51962, n51963, n51964,
         n51965, n51966, n51967, n51968, n51969, n51970, n51971, n51972,
         n51973, n51974, n51975, n51976, n51977, n51978, n51979, n51980,
         n51981, n51982, n51983, n51984, n51985, n51986, n51987, n51988,
         n51989, n51990, n51991, n51992, n51993, n51994, n51995, n51996,
         n51997, n51998, n51999, n52000, n52001, n52002, n52003, n52004,
         n52005, n52006, n52007, n52008, n52009, n52010, n52011, n52012,
         n52013, n52014, n52015, n52016, n52017, n52018, n52019, n52020,
         n52021, n52022, n52023, n52024, n52025, n52026, n52027, n52028,
         n52029, n52030, n52031, n52032, n52033, n52034, n52035, n52036,
         n52037, n52038, n52039, n52040, n52041, n52042, n52043, n52044,
         n52045, n52046, n52047, n52048, n52049, n52050, n52051, n52052,
         n52053, n52054, n52055, n52056, n52057, n52058, n52059, n52060,
         n52061, n52062, n52063, n52064, n52065, n52066, n52067, n52068,
         n52069, n52070, n52071, n52072, n52073, n52074, n52075, n52076,
         n52077, n52078, n52079, n52080, n52081, n52082, n52083, n52084,
         n52085, n52086, n52087, n52088, n52089, n52090, n52091, n52092,
         n52093, n52094, n52095, n52096, n52097, n52098, n52099, n52100,
         n52101, n52102, n52103, n52104, n52105, n52106, n52107, n52108,
         n52109, n52110, n52111, n52112, n52113, n52114, n52115, n52116,
         n52117, n52118, n52119, n52120, n52121, n52122, n52123, n52124,
         n52125, n52126, n52127, n52128, n52129, n52130, n52131, n52132,
         n52133, n52134, n52135, n52136, n52137, n52138, n52139, n52140,
         n52141, n52142, n52143, n52144, n52145, n52146, n52147, n52148,
         n52149, n52150, n52151, n52152, n52153, n52154, n52155, n52156,
         n52157, n52158, n52159, n52160, n52161, n52162, n52163, n52164,
         n52165, n52166, n52167, n52168, n52169, n52170, n52171, n52172,
         n52173, n52174, n52175, n52176, n52177, n52178, n52179, n52180,
         n52181, n52182, n52183, n52184, n52185, n52186, n52187, n52188,
         n52189, n52190, n52191, n52192, n52193, n52194, n52195, n52196,
         n52197, n52198, n52199, n52200, n52201, n52202, n52203, n52204,
         n52205, n52206, n52207, n52208, n52209, n52210, n52211, n52212,
         n52213, n52214, n52215, n52216, n52217, n52218, n52219, n52220,
         n52221, n52222, n52223, n52224, n52225, n52226, n52227, n52228,
         n52229, n52230, n52231, n52232, n52233, n52234, n52235, n52236,
         n52237, n52238, n52239, n52240, n52241, n52242, n52243, n52244,
         n52245, n52246, n52247, n52248, n52249, n52250, n52251, n52252,
         n52253, n52254, n52255, n52256, n52257, n52258, n52259, n52260,
         n52261, n52262, n52263, n52264, n52265, n52266, n52267, n52268,
         n52269, n52270, n52271, n52272, n52273, n52274, n52275, n52276,
         n52277, n52278, n52279, n52280, n52281, n52282, n52283, n52284,
         n52285, n52286, n52287, n52288, n52289, n52290, n52291, n52292,
         n52293, n52294, n52295, n52296, n52297, n52298, n52299, n52300,
         n52301, n52302, n52303, n52304, n52305, n52306, n52307, n52308,
         n52309, n52310, n52311, n52312, n52313, n52314, n52315, n52316,
         n52317, n52318, n52319, n52320, n52321, n52322, n52323, n52324,
         n52325, n52326, n52327, n52328, n52329, n52330, n52331, n52332,
         n52333, n52334, n52335, n52336, n52337, n52338, n52339, n52340,
         n52341, n52342, n52343, n52344, n52345, n52346, n52347, n52348,
         n52349, n52350, n52351, n52352, n52353, n52354, n52355, n52356,
         n52357, n52358, n52359, n52360, n52361, n52362, n52363, n52364,
         n52365, n52366, n52367, n52368, n52369, n52370, n52371, n52372,
         n52373, n52374, n52375, n52376, n52377, n52378, n52379, n52380,
         n52381, n52382, n52383, n52384, n52385, n52386, n52387, n52388,
         n52389, n52390, n52391, n52392, n52393, n52394, n52395, n52396,
         n52397, n52398, n52399, n52400, n52401, n52402, n52403, n52404,
         n52405, n52406, n52407, n52408, n52409, n52410, n52411, n52412,
         n52413, n52414, n52415, n52416, n52417, n52418, n52419, n52420,
         n52421, n52422, n52423, n52424, n52425, n52426, n52427, n52428,
         n52429, n52430, n52431, n52432, n52433, n52434, n52435, n52436,
         n52437, n52438, n52439, n52440, n52441, n52442, n52443, n52444,
         n52445, n52446, n52447, n52448, n52449, n52450, n52451, n52452,
         n52453, n52454, n52455, n52456, n52457, n52458, n52459, n52460,
         n52461, n52462, n52463, n52464, n52465, n52466, n52467, n52468,
         n52469, n52470, n52471, n52472, n52473, n52474, n52475, n52476,
         n52477, n52478, n52479, n52480, n52481, n52482, n52483, n52484,
         n52485, n52486, n52487, n52488, n52489, n52490, n52491, n52492,
         n52493, n52494, n52495, n52496, n52497, n52498, n52499, n52500,
         n52501, n52502, n52503, n52504, n52505, n52506, n52507, n52508,
         n52509, n52510, n52511, n52512, n52513, n52514, n52515, n52516,
         n52517, n52518, n52519, n52520, n52521, n52522, n52523, n52524,
         n52525, n52526, n52527, n52528, n52529, n52530, n52531, n52532,
         n52533, n52534, n52535, n52536, n52537, n52538, n52539, n52540,
         n52541, n52542, n52543, n52544, n52545, n52546, n52547, n52548,
         n52549, n52550, n52551, n52552, n52553, n52554, n52555, n52556,
         n52557, n52558, n52559, n52560, n52561, n52562, n52563, n52564,
         n52565, n52566, n52567, n52568, n52569, n52570, n52571, n52572,
         n52573, n52574, n52575, n52576, n52577, n52578, n52579, n52580,
         n52581, n52582, n52583, n52584, n52585, n52586, n52587, n52588,
         n52589, n52590, n52591, n52592, n52593, n52594, n52595, n52596,
         n52597, n52598, n52599, n52600, n52601, n52602, n52603, n52604,
         n52605, n52606, n52607, n52608, n52609, n52610, n52611, n52612,
         n52613, n52614, n52615, n52616, n52617, n52618, n52619, n52620,
         n52621, n52622, n52623, n52624, n52625, n52626, n52627, n52628,
         n52629, n52630, n52631, n52632, n52633, n52634, n52635, n52636,
         n52637, n52638, n52639, n52640, n52641, n52642, n52643, n52644,
         n52645, n52646, n52647, n52648, n52649, n52650, n52651, n52652,
         n52653, n52654, n52655, n52656, n52657, n52658, n52659, n52660,
         n52661, n52662, n52663, n52664, n52665, n52666, n52667, n52668,
         n52669, n52670, n52671, n52672, n52673, n52674, n52675, n52676,
         n52677, n52678, n52679, n52680, n52681, n52682, n52683, n52684,
         n52685, n52686, n52687, n52688, n52689, n52690, n52691, n52692,
         n52693, n52694, n52695, n52696, n52697, n52698, n52699, n52700,
         n52701, n52702, n52703, n52704, n52705, n52706, n52707, n52708,
         n52709, n52710, n52711, n52712, n52713, n52714, n52715, n52716,
         n52717, n52718, n52719, n52720, n52721, n52722, n52723, n52724,
         n52725, n52726, n52727, n52728, n52729, n52730, n52731, n52732,
         n52733, n52734, n52735, n52736, n52737, n52738, n52739, n52740,
         n52741, n52742, n52743, n52744, n52745, n52746, n52747, n52748,
         n52749, n52750, n52751, n52752, n52753, n52754, n52755, n52756,
         n52757, n52758, n52759, n52760, n52761, n52762, n52763, n52764,
         n52765, n52766, n52767, n52768, n52769, n52770, n52771, n52772,
         n52773, n52774, n52775, n52776, n52777, n52778, n52779, n52780,
         n52781, n52782, n52783, n52784, n52785, n52786, n52787, n52788,
         n52789, n52790, n52791, n52792, n52793, n52794, n52795, n52796,
         n52797, n52798, n52799, n52800, n52801, n52802, n52803, n52804,
         n52805, n52806, n52807, n52808, n52809, n52810, n52811, n52812,
         n52813, n52814, n52815, n52816, n52817, n52818, n52819, n52820,
         n52821, n52822, n52823, n52824, n52825, n52826, n52827, n52828,
         n52829, n52830, n52831, n52832, n52833, n52834, n52835, n52836,
         n52837, n52838, n52839, n52840, n52841, n52842, n52843, n52844,
         n52845, n52846, n52847, n52848, n52849, n52850, n52851, n52852,
         n52853, n52854, n52855, n52856, n52857, n52858, n52859, n52860,
         n52861, n52862, n52863, n52864, n52865, n52866, n52867, n52868,
         n52869, n52870, n52871, n52872, n52873, n52874, n52875, n52876,
         n52877, n52878, n52879, n52880, n52881, n52882, n52883, n52884,
         n52885, n52886, n52887, n52888, n52889, n52890, n52891, n52892,
         n52893, n52894, n52895, n52896, n52897, n52898, n52899, n52900,
         n52901, n52902, n52903, n52904, n52905, n52906, n52907, n52908,
         n52909, n52910, n52911, n52912, n52913, n52914, n52915, n52916,
         n52917, n52918, n52919, n52920, n52921, n52922, n52923, n52924,
         n52925, n52926, n52927, n52928, n52929, n52930, n52931, n52932,
         n52933, n52934, n52935, n52936, n52937, n52938, n52939, n52940,
         n52941, n52942, n52943, n52944, n52945, n52946, n52947, n52948,
         n52949, n52950, n52951, n52952, n52953, n52954, n52955, n52956,
         n52957, n52958, n52959, n52960, n52961, n52962, n52963, n52964,
         n52965, n52966, n52967, n52968, n52969, n52970, n52971, n52972,
         n52973, n52974, n52975, n52976, n52977, n52978, n52979, n52980,
         n52981, n52982, n52983, n52984, n52985, n52986, n52987, n52988,
         n52989, n52990, n52991, n52992, n52993, n52994, n52995, n52996,
         n52997, n52998, n52999, n53000, n53001, n53002, n53003, n53004,
         n53005, n53006, n53007, n53008, n53009, n53010, n53011, n53012,
         n53013, n53014, n53015, n53016, n53017, n53018, n53019, n53020,
         n53021, n53022, n53023, n53024, n53025, n53026, n53027, n53028,
         n53029, n53030, n53031, n53032, n53033, n53034, n53035, n53036,
         n53037, n53038, n53039, n53040, n53041, n53042, n53043, n53044,
         n53045, n53046, n53047, n53048, n53049, n53050, n53051, n53052,
         n53053, n53054, n53055, n53056, n53057, n53058, n53059, n53060,
         n53061, n53062, n53063, n53064, n53065, n53066, n53067, n53068,
         n53069, n53070, n53071, n53072, n53073, n53074, n53075, n53076,
         n53077, n53078, n53079, n53080, n53081, n53082, n53083, n53084,
         n53085, n53086, n53087, n53088, n53089, n53090, n53091, n53092,
         n53093, n53094, n53095, n53096, n53097, n53098, n53099, n53100,
         n53101, n53102, n53103, n53104, n53105, n53106, n53107, n53108,
         n53109, n53110, n53111, n53112, n53113, n53114, n53115, n53116,
         n53117, n53118, n53119, n53120, n53121, n53122, n53123, n53124,
         n53125, n53126, n53127, n53128, n53129, n53130, n53131, n53132,
         n53133, n53134, n53135, n53136, n53137, n53138, n53139, n53140,
         n53141, n53142, n53143, n53144, n53145, n53146, n53147, n53148,
         n53149, n53150, n53151, n53152, n53153, n53154, n53155, n53156,
         n53157, n53158, n53159, n53160, n53161, n53162, n53163, n53164,
         n53165, n53166, n53167, n53168, n53169, n53170, n53171, n53172,
         n53173, n53174, n53175, n53176, n53177, n53178, n53179, n53180,
         n53181, n53182, n53183, n53184, n53185, n53186, n53187, n53188,
         n53189, n53190, n53191, n53192, n53193, n53194, n53195, n53196,
         n53197, n53198, n53199, n53200, n53201, n53202, n53203, n53204,
         n53205, n53206, n53207, n53208, n53209, n53210, n53211, n53212,
         n53213, n53214, n53215, n53216, n53217, n53218, n53219, n53220,
         n53221, n53222, n53223, n53224, n53225, n53226, n53227, n53228,
         n53229, n53230, n53231, n53232, n53233, n53234, n53235, n53236,
         n53237, n53238, n53239, n53240, n53241, n53242, n53243, n53244,
         n53245, n53246, n53247, n53248, n53249, n53250, n53251, n53252,
         n53253, n53254, n53255, n53256, n53257, n53258, n53259, n53260,
         n53261, n53262, n53263, n53264, n53265, n53266, n53267, n53268,
         n53269, n53270, n53271, n53272, n53273, n53274, n53275, n53276,
         n53277, n53278, n53279, n53280, n53281, n53282, n53283, n53284,
         n53285, n53286, n53287, n53288, n53289, n53290, n53291, n53292,
         n53293, n53294, n53295, n53296, n53297, n53298, n53299, n53300,
         n53301, n53302, n53303, n53304, n53305, n53306, n53307, n53308,
         n53309, n53310, n53311, n53312, n53313, n53314, n53315, n53316,
         n53317, n53318, n53319, n53320, n53321, n53322, n53323, n53324,
         n53325, n53326, n53327, n53328, n53329, n53330, n53331, n53332,
         n53333, n53334, n53335, n53336, n53337, n53338, n53339, n53340,
         n53341, n53342, n53343, n53344, n53345, n53346, n53347, n53348,
         n53349, n53350, n53351, n53352, n53353, n53354, n53355, n53356,
         n53357, n53358, n53359, n53360, n53361, n53362, n53363, n53364,
         n53365, n53366, n53367, n53368, n53369, n53370, n53371, n53372,
         n53373, n53374, n53375, n53376, n53377, n53378, n53379, n53380,
         n53381, n53382, n53383, n53384, n53385, n53386, n53387, n53388,
         n53389, n53390, n53391, n53392, n53393, n53394, n53395, n53396,
         n53397, n53398, n53399, n53400, n53401, n53402, n53403, n53404,
         n53405, n53406, n53407, n53408, n53409, n53410, n53411, n53412,
         n53413, n53414, n53415, n53416, n53417, n53418, n53419, n53420,
         n53421, n53422, n53423, n53424, n53425, n53426, n53427, n53428,
         n53429, n53430, n53431, n53432, n53433, n53434, n53435, n53436,
         n53437, n53438, n53439, n53440, n53441, n53442, n53443, n53444,
         n53445, n53446, n53447, n53448, n53449, n53450, n53451, n53452,
         n53453, n53454, n53455, n53456, n53457, n53458, n53459, n53460,
         n53461, n53462, n53463, n53464, n53465, n53466, n53467, n53468,
         n53469, n53470, n53471, n53472, n53473, n53474, n53475, n53476,
         n53477, n53478, n53479, n53480, n53481, n53482, n53483, n53484,
         n53485, n53486, n53487, n53488, n53489, n53490, n53491, n53492,
         n53493, n53494, n53495, n53496, n53497, n53498, n53499, n53500,
         n53501, n53502, n53503, n53504, n53505, n53506, n53507, n53508,
         n53509, n53510, n53511, n53512, n53513, n53514, n53515, n53516,
         n53517, n53518, n53519, n53520, n53521, n53522, n53523, n53524,
         n53525, n53526, n53527, n53528, n53529, n53530, n53531, n53532,
         n53533, n53534, n53535, n53536, n53537, n53538, n53539, n53540,
         n53541, n53542, n53543, n53544, n53545, n53546, n53547, n53548,
         n53549, n53550, n53551, n53552, n53553, n53554, n53555, n53556,
         n53557, n53558, n53559, n53560, n53561, n53562, n53563, n53564,
         n53565, n53566, n53567, n53568, n53569, n53570, n53571, n53572,
         n53573, n53574, n53575, n53576, n53577, n53578, n53579, n53580,
         n53581, n53582, n53583, n53584, n53585, n53586, n53587, n53588,
         n53589, n53590, n53591, n53592, n53593, n53594, n53595, n53596,
         n53597, n53598, n53599, n53600, n53601, n53602, n53603, n53604,
         n53605, n53606, n53607, n53608, n53609, n53610, n53611, n53612,
         n53613, n53614, n53615, n53616, n53617, n53618, n53619, n53620,
         n53621, n53622, n53623, n53624, n53625, n53626, n53627, n53628,
         n53629, n53630, n53631, n53632, n53633, n53634, n53635, n53636,
         n53637, n53638, n53639, n53640, n53641, n53642, n53643, n53644,
         n53645, n53646, n53647, n53648, n53649, n53650, n53651, n53652,
         n53653, n53654, n53655, n53656, n53657, n53658, n53659, n53660,
         n53661, n53662, n53663, n53664, n53665, n53666, n53667, n53668,
         n53669, n53670, n53671, n53672, n53673, n53674, n53675, n53676,
         n53677, n53678, n53679, n53680, n53681, n53682, n53683, n53684,
         n53685, n53686, n53687, n53688, n53689, n53690, n53691, n53692,
         n53693, n53694, n53695, n53696, n53697, n53698, n53699, n53700,
         n53701, n53702, n53703, n53704, n53705, n53706, n53707, n53708,
         n53709, n53710, n53711, n53712, n53713, n53714, n53715, n53716,
         n53717, n53718, n53719, n53720, n53721, n53722, n53723, n53724,
         n53725, n53726, n53727, n53728, n53729, n53730, n53731, n53732,
         n53733, n53734, n53735, n53736, n53737, n53738, n53739, n53740,
         n53741, n53742, n53743, n53744, n53745, n53746, n53747, n53748,
         n53749, n53750, n53751, n53752, n53753, n53754, n53755, n53756,
         n53757, n53758, n53759, n53760, n53761, n53762, n53763, n53764,
         n53765, n53766, n53767, n53768, n53769, n53770, n53771, n53772,
         n53773, n53774, n53775, n53776, n53777, n53778, n53779, n53780,
         n53781, n53782, n53783, n53784, n53785, n53786, n53787, n53788,
         n53789, n53790, n53791, n53792, n53793, n53794, n53795, n53796,
         n53797, n53798, n53799, n53800, n53801, n53802, n53803, n53804,
         n53805, n53806, n53807, n53808, n53809, n53810, n53811, n53812,
         n53813, n53814, n53815, n53816, n53817, n53818, n53819, n53820,
         n53821, n53822, n53823, n53824, n53825, n53826, n53827, n53828,
         n53829, n53830, n53831, n53832, n53833, n53834, n53835, n53836,
         n53837, n53838, n53839, n53840, n53841, n53842, n53843, n53844,
         n53845, n53846, n53847, n53848, n53849, n53850, n53851, n53852,
         n53853, n53854, n53855, n53856, n53857, n53858, n53859, n53860,
         n53861, n53862, n53863, n53864, n53865, n53866, n53867, n53868,
         n53869, n53870, n53871, n53872, n53873, n53874, n53875, n53876,
         n53877, n53878, n53879, n53880, n53881, n53882, n53883, n53884,
         n53885, n53886, n53887, n53888, n53889, n53890, n53891, n53892,
         n53893, n53894, n53895, n53896, n53897, n53898, n53899, n53900,
         n53901, n53902, n53903, n53904, n53905, n53906, n53907, n53908,
         n53909, n53910, n53911, n53912, n53913, n53914, n53915, n53916,
         n53917, n53918, n53919, n53920, n53921, n53922, n53923, n53924,
         n53925, n53926, n53927, n53928, n53929, n53930, n53931, n53932,
         n53933, n53934, n53935, n53936, n53937, n53938, n53939, n53940,
         n53941, n53942, n53943, n53944, n53945, n53946, n53947, n53948,
         n53949, n53950, n53951, n53952, n53953, n53954, n53955, n53956,
         n53957, n53958, n53959, n53960, n53961, n53962, n53963, n53964,
         n53965, n53966, n53967, n53968, n53969, n53970, n53971, n53972,
         n53973, n53974, n53975, n53976, n53977, n53978, n53979, n53980,
         n53981, n53982, n53983, n53984, n53985, n53986, n53987, n53988,
         n53989, n53990, n53991, n53992, n53993, n53994, n53995, n53996,
         n53997, n53998, n53999, n54000, n54001, n54002, n54003, n54004,
         n54005, n54006, n54007, n54008, n54009, n54010, n54011, n54012,
         n54013, n54014, n54015, n54016, n54017, n54018, n54019, n54020,
         n54021, n54022, n54023, n54024, n54025, n54026, n54027, n54028,
         n54029, n54030, n54031, n54032, n54033, n54034, n54035, n54036,
         n54037, n54038, n54039, n54040, n54041, n54042, n54043, n54044,
         n54045, n54046, n54047, n54048, n54049, n54050, n54051, n54052,
         n54053, n54054, n54055, n54056, n54057, n54058, n54059, n54060,
         n54061, n54062, n54063, n54064, n54065, n54066, n54067, n54068,
         n54069, n54070, n54071, n54072, n54073, n54074, n54075, n54076,
         n54077, n54078, n54079, n54080, n54081, n54082, n54083, n54084,
         n54085, n54086, n54087, n54088, n54089, n54090, n54091, n54092,
         n54093, n54094, n54095, n54096, n54097, n54098, n54099, n54100,
         n54101, n54102, n54103, n54104, n54105, n54106, n54107, n54108,
         n54109, n54110, n54111, n54112, n54113, n54114, n54115, n54116,
         n54117, n54118, n54119, n54120, n54121, n54122, n54123, n54124,
         n54125, n54126, n54127, n54128, n54129, n54130, n54131, n54132,
         n54133, n54134, n54135, n54136, n54137, n54138, n54139, n54140,
         n54141, n54142, n54143, n54144, n54145, n54146, n54147, n54148,
         n54149, n54150, n54151, n54152, n54153, n54154, n54155, n54156,
         n54157, n54158, n54159, n54160, n54161, n54162, n54163, n54164,
         n54165, n54166, n54167, n54168, n54169, n54170, n54171, n54172,
         n54173, n54174, n54175, n54176, n54177, n54178, n54179, n54180,
         n54181, n54182, n54183, n54184, n54185, n54186, n54187, n54188,
         n54189, n54190, n54191, n54192, n54193, n54194, n54195, n54196,
         n54197, n54198, n54199, n54200, n54201, n54202, n54203, n54204,
         n54205, n54206, n54207, n54208, n54209, n54210, n54211, n54212,
         n54213, n54214, n54215, n54216, n54217, n54218, n54219, n54220,
         n54221, n54222, n54223, n54224, n54225, n54226, n54227, n54228,
         n54229, n54230, n54231, n54232, n54233, n54234, n54235, n54236,
         n54237, n54238, n54239, n54240, n54241, n54242, n54243, n54244,
         n54245, n54246, n54247, n54248, n54249, n54250, n54251, n54252,
         n54253, n54254, n54255, n54256, n54257, n54258, n54259, n54260,
         n54261, n54262, n54263, n54264, n54265, n54266, n54267, n54268,
         n54269, n54270, n54271, n54272, n54273, n54274, n54275, n54276,
         n54277, n54278, n54279, n54280, n54281, n54282, n54283, n54284,
         n54285, n54286, n54287, n54288, n54289, n54290, n54291, n54292,
         n54293, n54294, n54295, n54296, n54297, n54298, n54299, n54300,
         n54301, n54302, n54303, n54304, n54305, n54306, n54307, n54308,
         n54309, n54310, n54311, n54312, n54313, n54314, n54315, n54316,
         n54317, n54318, n54319, n54320, n54321, n54322, n54323, n54324,
         n54325, n54326, n54327, n54328, n54329, n54330, n54331, n54332,
         n54333, n54334, n54335, n54336, n54337, n54338, n54339, n54340,
         n54341, n54342, n54343, n54344, n54345, n54346, n54347, n54348,
         n54349, n54350, n54351, n54352, n54353, n54354, n54355, n54356,
         n54357, n54358, n54359, n54360, n54361, n54362, n54363, n54364,
         n54365, n54366, n54367, n54368, n54369, n54370, n54371, n54372,
         n54373, n54374, n54375, n54376, n54377, n54378, n54379, n54380,
         n54381, n54382, n54383, n54384, n54385, n54386, n54387, n54388,
         n54389, n54390, n54391, n54392, n54393, n54394, n54395, n54396,
         n54397, n54398, n54399, n54400, n54401, n54402, n54403, n54404,
         n54405, n54406, n54407, n54408, n54409, n54410, n54411, n54412,
         n54413, n54414, n54415, n54416, n54417, n54418, n54419, n54420,
         n54421, n54422, n54423, n54424, n54425, n54426, n54427, n54428,
         n54429, n54430, n54431, n54432, n54433, n54434, n54435, n54436,
         n54437, n54438, n54439, n54440, n54441, n54442, n54443, n54444,
         n54445, n54446, n54447, n54448, n54449, n54450, n54451, n54452,
         n54453, n54454, n54455, n54456, n54457, n54458, n54459, n54460,
         n54461, n54462, n54463, n54464, n54465, n54466, n54467, n54468,
         n54469, n54470, n54471, n54472, n54473, n54474, n54475, n54476,
         n54477, n54478, n54479, n54480, n54481, n54482, n54483, n54484,
         n54485, n54486, n54487, n54488, n54489, n54490, n54491, n54492,
         n54493, n54494, n54495, n54496, n54497, n54498, n54499, n54500,
         n54501, n54502, n54503, n54504, n54505, n54506, n54507, n54508,
         n54509, n54510, n54511, n54512, n54513, n54514, n54515, n54516,
         n54517, n54518, n54519, n54520, n54521, n54522, n54523, n54524,
         n54525, n54526, n54527, n54528, n54529, n54530, n54531, n54532,
         n54533, n54534, n54535, n54536, n54537, n54538, n54539, n54540,
         n54541, n54542, n54543, n54544, n54545, n54546, n54547, n54548,
         n54549, n54550, n54551, n54552, n54553, n54554, n54555, n54556,
         n54557, n54558, n54559, n54560, n54561, n54562, n54563, n54564,
         n54565, n54566, n54567, n54568, n54569, n54570, n54571, n54572,
         n54573, n54574, n54575, n54576, n54577, n54578, n54579, n54580,
         n54581, n54582, n54583, n54584, n54585, n54586, n54587, n54588,
         n54589, n54590, n54591, n54592, n54593, n54594, n54595, n54596,
         n54597, n54598, n54599, n54600, n54601, n54602, n54603, n54604,
         n54605, n54606, n54607, n54608, n54609, n54610, n54611, n54612,
         n54613, n54614, n54615, n54616, n54617, n54618, n54619, n54620,
         n54621, n54622, n54623, n54624, n54625, n54626, n54627, n54628,
         n54629, n54630, n54631, n54632, n54633, n54634, n54635, n54636,
         n54637, n54638, n54639, n54640, n54641, n54642, n54643, n54644,
         n54645, n54646, n54647, n54648, n54649, n54650, n54651, n54652,
         n54653, n54654, n54655, n54656, n54657, n54658, n54659, n54660,
         n54661, n54662, n54663, n54664, n54665, n54666, n54667, n54668,
         n54669, n54670, n54671, n54672, n54673, n54674, n54675, n54676,
         n54677, n54678, n54679, n54680, n54681, n54682, n54683, n54684,
         n54685, n54686, n54687, n54688, n54689, n54690, n54691, n54692,
         n54693, n54694, n54695, n54696, n54697, n54698, n54699, n54700,
         n54701, n54702, n54703, n54704, n54705, n54706, n54707, n54708,
         n54709, n54710, n54711, n54712, n54713, n54714, n54715, n54716,
         n54717, n54718, n54719, n54720, n54721, n54722, n54723, n54724,
         n54725, n54726, n54727, n54728, n54729, n54730, n54731, n54732,
         n54733, n54734, n54735, n54736, n54737, n54738, n54739, n54740,
         n54741, n54742, n54743, n54744, n54745, n54746, n54747, n54748,
         n54749, n54750, n54751, n54752, n54753, n54754, n54755, n54756,
         n54757, n54758, n54759, n54760, n54761, n54762, n54763, n54764,
         n54765, n54766, n54767, n54768, n54769, n54770, n54771, n54772,
         n54773, n54774, n54775, n54776, n54777, n54778, n54779, n54780,
         n54781, n54782, n54783, n54784, n54785, n54786, n54787, n54788,
         n54789, n54790, n54791, n54792, n54793, n54794, n54795, n54796,
         n54797, n54798, n54799, n54800, n54801, n54802, n54803, n54804,
         n54805, n54806, n54807, n54808, n54809, n54810, n54811, n54812,
         n54813, n54814, n54815, n54816, n54817, n54818, n54819, n54820,
         n54821, n54822, n54823, n54824, n54825, n54826, n54827, n54828,
         n54829, n54830, n54831, n54832, n54833, n54834, n54835, n54836,
         n54837, n54838, n54839, n54840, n54841, n54842, n54843, n54844,
         n54845, n54846, n54847, n54848, n54849, n54850, n54851, n54852,
         n54853, n54854, n54855, n54856, n54857, n54858, n54859, n54860,
         n54861, n54862, n54863, n54864, n54865, n54866, n54867, n54868,
         n54869, n54870, n54871, n54872, n54873, n54874, n54875, n54876,
         n54877, n54878, n54879, n54880, n54881, n54882, n54883, n54884,
         n54885, n54886, n54887, n54888, n54889, n54890, n54891, n54892,
         n54893, n54894, n54895, n54896, n54897, n54898, n54899, n54900,
         n54901, n54902, n54903, n54904, n54905, n54906, n54907, n54908,
         n54909, n54910, n54911, n54912, n54913, n54914, n54915, n54916,
         n54917, n54918, n54919, n54920, n54921, n54922, n54923, n54924,
         n54925, n54926, n54927, n54928, n54929, n54930, n54931, n54932,
         n54933, n54934, n54935, n54936, n54937, n54938, n54939, n54940,
         n54941, n54942, n54943, n54944, n54945, n54946, n54947, n54948,
         n54949, n54950, n54951, n54952, n54953, n54954, n54955, n54956,
         n54957, n54958, n54959, n54960, n54961, n54962, n54963, n54964,
         n54965, n54966, n54967, n54968, n54969, n54970, n54971, n54972,
         n54973, n54974, n54975, n54976, n54977, n54978, n54979, n54980,
         n54981, n54982, n54983, n54984, n54985, n54986, n54987, n54988,
         n54989, n54990, n54991, n54992, n54993, n54994, n54995, n54996,
         n54997, n54998, n54999, n55000, n55001, n55002, n55003, n55004,
         n55005, n55006, n55007, n55008, n55009, n55010, n55011, n55012,
         n55013, n55014, n55015, n55016, n55017, n55018, n55019, n55020,
         n55021, n55022, n55023, n55024, n55025, n55026, n55027, n55028,
         n55029, n55030, n55031, n55032, n55033, n55034, n55035, n55036,
         n55037, n55038, n55039, n55040, n55041, n55042, n55043, n55044,
         n55045, n55046, n55047, n55048, n55049, n55050, n55051, n55052,
         n55053, n55054, n55055, n55056, n55057, n55058, n55059, n55060,
         n55061, n55062, n55063, n55064, n55065, n55066, n55067, n55068,
         n55069, n55070, n55071, n55072, n55073, n55074, n55075, n55076,
         n55077, n55078, n55079, n55080, n55081, n55082, n55083, n55084,
         n55085, n55086, n55087, n55088, n55089, n55090, n55091, n55092,
         n55093, n55094, n55095, n55096, n55097, n55098, n55099, n55100,
         n55101, n55102, n55103, n55104, n55105, n55106, n55107, n55108,
         n55109, n55110, n55111, n55112, n55113, n55114, n55115, n55116,
         n55117, n55118, n55119, n55120, n55121, n55122, n55123, n55124,
         n55125, n55126, n55127, n55128, n55129, n55130, n55131, n55132,
         n55133, n55134, n55135, n55136, n55137, n55138, n55139, n55140,
         n55141, n55142, n55143, n55144, n55145, n55146, n55147, n55148,
         n55149, n55150, n55151, n55152, n55153, n55154, n55155, n55156,
         n55157, n55158, n55159, n55160, n55161, n55162, n55163, n55164,
         n55165, n55166, n55167, n55168, n55169, n55170, n55171, n55172,
         n55173, n55174, n55175, n55176, n55177, n55178, n55179, n55180,
         n55181, n55182, n55183, n55184, n55185, n55186, n55187, n55188,
         n55189, n55190, n55191, n55192, n55193, n55194, n55195, n55196,
         n55197, n55198, n55199, n55200, n55201, n55202, n55203, n55204,
         n55205, n55206, n55207, n55208, n55209, n55210, n55211, n55212,
         n55213, n55214, n55215, n55216, n55217, n55218, n55219, n55220,
         n55221, n55222, n55223, n55224, n55225, n55226, n55227, n55228,
         n55229, n55230, n55231, n55232, n55233, n55234, n55235, n55236,
         n55237, n55238, n55239, n55240, n55241, n55242, n55243, n55244,
         n55245, n55246, n55247, n55248, n55249, n55250, n55251, n55252,
         n55253, n55254, n55255, n55256, n55257, n55258, n55259, n55260,
         n55261, n55262, n55263, n55264, n55265, n55266, n55267, n55268,
         n55269, n55270, n55271, n55272, n55273, n55274, n55275, n55276,
         n55277, n55278, n55279, n55280, n55281, n55282, n55283, n55284,
         n55285, n55286, n55287, n55288, n55289, n55290, n55291, n55292,
         n55293, n55294, n55295, n55296, n55297, n55298, n55299, n55300,
         n55301, n55302, n55303, n55304, n55305, n55306, n55307, n55308,
         n55309, n55310, n55311, n55312, n55313, n55314, n55315, n55316,
         n55317, n55318, n55319, n55320, n55321, n55322, n55323, n55324,
         n55325, n55326, n55327, n55328, n55329, n55330, n55331, n55332,
         n55333, n55334, n55335, n55336, n55337, n55338, n55339, n55340,
         n55341, n55342, n55343, n55344, n55345, n55346, n55347, n55348,
         n55349, n55350, n55351, n55352, n55353, n55354, n55355, n55356,
         n55357, n55358, n55359, n55360, n55361, n55362, n55363, n55364,
         n55365, n55366, n55367, n55368, n55369, n55370, n55371, n55372,
         n55373, n55374, n55375, n55376, n55377, n55378, n55379, n55380,
         n55381, n55382, n55383, n55384, n55385, n55386, n55387, n55388,
         n55389, n55390, n55391, n55392, n55393, n55394, n55395, n55396,
         n55397, n55398, n55399, n55400, n55401, n55402, n55403, n55404,
         n55405, n55406, n55407, n55408, n55409, n55410, n55411, n55412,
         n55413, n55414, n55415, n55416, n55417, n55418, n55419, n55420,
         n55421, n55422, n55423, n55424, n55425, n55426, n55427, n55428,
         n55429, n55430, n55431, n55432, n55433, n55434, n55435, n55436,
         n55437, n55438, n55439, n55440, n55441, n55442, n55443, n55444,
         n55445, n55446, n55447, n55448, n55449, n55450, n55451, n55452,
         n55453, n55454, n55455, n55456, n55457, n55458, n55459, n55460,
         n55461, n55462, n55463, n55464, n55465, n55466, n55467, n55468,
         n55469, n55470, n55471, n55472, n55473, n55474, n55475, n55476,
         n55477, n55478, n55479, n55480, n55481, n55482, n55483, n55484,
         n55485, n55486, n55487, n55488, n55489, n55490, n55491, n55492,
         n55493, n55494, n55495, n55496, n55497, n55498, n55499, n55500,
         n55501, n55502, n55503, n55504, n55505, n55506, n55507, n55508,
         n55509, n55510, n55511, n55512, n55513, n55514, n55515, n55516,
         n55517, n55518, n55519, n55520, n55521, n55522, n55523, n55524,
         n55525, n55526, n55527, n55528, n55529, n55530, n55531, n55532,
         n55533, n55534, n55535, n55536, n55537, n55538, n55539, n55540,
         n55541, n55542, n55543, n55544, n55545, n55546, n55547, n55548,
         n55549, n55550, n55551, n55552, n55553, n55554, n55555, n55556,
         n55557, n55558, n55559, n55560, n55561, n55562, n55563, n55564,
         n55565, n55566, n55567, n55568, n55569, n55570, n55571, n55572,
         n55573, n55574, n55575, n55576, n55577, n55578, n55579, n55580,
         n55581, n55582, n55583, n55584, n55585, n55586, n55587, n55588,
         n55589, n55590, n55591, n55592, n55593, n55594, n55595, n55596,
         n55597, n55598, n55599, n55600, n55601, n55602, n55603, n55604,
         n55605, n55606, n55607, n55608, n55609, n55610, n55611, n55612,
         n55613, n55614, n55615, n55616, n55617, n55618, n55619, n55620,
         n55621, n55622, n55623, n55624, n55625, n55626, n55627, n55628,
         n55629, n55630, n55631, n55632, n55633, n55634, n55635, n55636,
         n55637, n55638, n55639, n55640, n55641, n55642, n55643, n55644,
         n55645, n55646, n55647, n55648, n55649, n55650, n55651, n55652,
         n55653, n55654, n55655, n55656, n55657, n55658, n55659, n55660,
         n55661, n55662, n55663, n55664, n55665, n55666, n55667, n55668,
         n55669, n55670, n55671, n55672, n55673, n55674, n55675, n55676,
         n55677, n55678, n55679, n55680, n55681, n55682, n55683, n55684,
         n55685, n55686, n55687, n55688, n55689, n55690, n55691, n55692,
         n55693, n55694, n55695, n55696, n55697, n55698, n55699, n55700,
         n55701, n55702, n55703, n55704, n55705, n55706, n55707, n55708,
         n55709, n55710, n55711, n55712, n55713, n55714, n55715, n55716,
         n55717, n55718, n55719, n55720, n55721, n55722, n55723, n55724,
         n55725, n55726, n55727, n55728, n55729, n55730, n55731, n55732,
         n55733, n55734, n55735, n55736, n55737, n55738, n55739, n55740,
         n55741, n55742, n55743, n55744, n55745, n55746, n55747, n55748,
         n55749, n55750, n55751, n55752, n55753, n55754, n55755, n55756,
         n55757, n55758, n55759, n55760, n55761, n55762, n55763, n55764,
         n55765, n55766, n55767, n55768, n55769, n55770, n55771, n55772,
         n55773, n55774, n55775, n55776, n55777, n55778, n55779, n55780,
         n55781, n55782, n55783, n55784, n55785, n55786, n55787, n55788,
         n55789, n55790, n55791, n55792, n55793, n55794, n55795, n55796,
         n55797, n55798, n55799, n55800, n55801, n55802, n55803, n55804,
         n55805, n55806, n55807, n55808, n55809, n55810, n55811, n55812,
         n55813, n55814, n55815, n55816, n55817, n55818, n55819, n55820,
         n55821, n55822, n55823, n55824, n55825, n55826, n55827, n55828,
         n55829, n55830, n55831, n55832, n55833, n55834, n55835, n55836,
         n55837, n55838, n55839, n55840, n55841, n55842, n55843, n55844,
         n55845, n55846, n55847, n55848, n55849, n55850, n55851, n55852,
         n55853, n55854, n55855, n55856, n55857, n55858, n55859, n55860,
         n55861, n55862, n55863, n55864, n55865, n55866, n55867, n55868,
         n55869, n55870, n55871, n55872, n55873, n55874, n55875, n55876,
         n55877, n55878, n55879, n55880, n55881, n55882, n55883, n55884,
         n55885, n55886, n55887, n55888, n55889, n55890, n55891, n55892,
         n55893, n55894, n55895, n55896, n55897, n55898, n55899, n55900,
         n55901, n55902, n55903, n55904, n55905, n55906, n55907, n55908,
         n55909, n55910, n55911, n55912, n55913, n55914, n55915, n55916,
         n55917, n55918, n55919, n55920, n55921, n55922, n55923, n55924,
         n55925, n55926, n55927, n55928, n55929, n55930, n55931, n55932,
         n55933, n55934, n55935, n55936, n55937, n55938, n55939, n55940,
         n55941, n55942, n55943, n55944, n55945, n55946, n55947, n55948,
         n55949, n55950, n55951, n55952, n55953, n55954, n55955, n55956,
         n55957, n55958, n55959, n55960, n55961, n55962, n55963, n55964,
         n55965, n55966, n55967, n55968, n55969, n55970, n55971, n55972,
         n55973, n55974, n55975, n55976, n55977, n55978, n55979, n55980,
         n55981, n55982, n55983, n55984, n55985, n55986, n55987, n55988,
         n55989, n55990, n55991, n55992, n55993, n55994, n55995, n55996,
         n55997, n55998, n55999, n56000, n56001, n56002, n56003, n56004,
         n56005, n56006, n56007, n56008, n56009, n56010, n56011, n56012,
         n56013, n56014, n56015, n56016, n56017, n56018, n56019, n56020,
         n56021, n56022, n56023, n56024, n56025, n56026, n56027, n56028,
         n56029, n56030, n56031, n56032, n56033, n56034, n56035, n56036,
         n56037, n56038, n56039, n56040, n56041, n56042, n56043, n56044,
         n56045, n56046, n56047, n56048, n56049, n56050, n56051, n56052,
         n56053, n56054, n56055, n56056, n56057, n56058, n56059, n56060,
         n56061, n56062, n56063, n56064, n56065, n56066, n56067, n56068,
         n56069, n56070, n56071, n56072, n56073, n56074, n56075, n56076,
         n56077, n56078, n56079, n56080, n56081, n56082, n56083, n56084,
         n56085, n56086, n56087, n56088, n56089, n56090, n56091, n56092,
         n56093, n56094, n56095, n56096, n56097, n56098, n56099, n56100,
         n56101, n56102, n56103, n56104, n56105, n56106, n56107, n56108,
         n56109, n56110, n56111, n56112, n56113, n56114, n56115, n56116,
         n56117, n56118, n56119, n56120, n56121, n56122, n56123, n56124,
         n56125, n56126, n56127, n56128, n56129, n56130, n56131, n56132,
         n56133, n56134, n56135, n56136, n56137, n56138, n56139, n56140,
         n56141, n56142, n56143, n56144, n56145, n56146, n56147, n56148,
         n56149, n56150, n56151, n56152, n56153, n56154, n56155, n56156,
         n56157, n56158, n56159, n56160, n56161, n56162, n56163, n56164,
         n56165, n56166, n56167, n56168, n56169, n56170, n56171, n56172,
         n56173, n56174, n56175, n56176, n56177, n56178, n56179, n56180,
         n56181, n56182, n56183, n56184, n56185, n56186, n56187, n56188,
         n56189, n56190, n56191, n56192, n56193, n56194, n56195, n56196,
         n56197, n56198, n56199, n56200, n56201, n56202, n56203, n56204,
         n56205, n56206, n56207, n56208, n56209, n56210, n56211, n56212,
         n56213, n56214, n56215, n56216, n56217, n56218, n56219, n56220,
         n56221, n56222, n56223, n56224, n56225, n56226, n56227, n56228,
         n56229, n56230, n56231, n56232, n56233, n56234, n56235, n56236,
         n56237, n56238, n56239, n56240, n56241, n56242, n56243, n56244,
         n56245, n56246, n56247, n56248, n56249, n56250, n56251, n56252,
         n56253, n56254, n56255, n56256, n56257, n56258, n56259, n56260,
         n56261, n56262, n56263, n56264, n56265, n56266, n56267, n56268,
         n56269, n56270, n56271, n56272, n56273, n56274, n56275, n56276,
         n56277, n56278, n56279, n56280, n56281, n56282, n56283, n56284,
         n56285, n56286, n56287, n56288, n56289, n56290, n56291, n56292,
         n56293, n56294, n56295, n56296, n56297, n56298, n56299, n56300,
         n56301, n56302, n56303, n56304, n56305, n56306, n56307, n56308,
         n56309, n56310, n56311, n56312, n56313, n56314, n56315, n56316,
         n56317, n56318, n56319, n56320, n56321, n56322, n56323, n56324,
         n56325, n56326, n56327, n56328, n56329, n56330, n56331, n56332,
         n56333, n56334, n56335, n56336, n56337, n56338, n56339, n56340,
         n56341, n56342, n56343, n56344, n56345, n56346, n56347, n56348,
         n56349, n56350, n56351, n56352, n56353, n56354, n56355, n56356,
         n56357, n56358, n56359, n56360, n56361, n56362, n56363, n56364,
         n56365, n56366, n56367, n56368, n56369, n56370, n56371, n56372,
         n56373, n56374, n56375, n56376, n56377, n56378, n56379, n56380,
         n56381, n56382, n56383, n56384, n56385, n56386, n56387, n56388,
         n56389, n56390, n56391, n56392, n56393, n56394, n56395, n56396,
         n56397, n56398, n56399, n56400, n56401, n56402, n56403, n56404,
         n56405, n56406, n56407, n56408, n56409, n56410, n56411, n56412,
         n56413, n56414, n56415, n56416, n56417, n56418, n56419, n56420,
         n56421, n56422, n56423, n56424, n56425, n56426, n56427, n56428,
         n56429, n56430, n56431, n56432, n56433, n56434, n56435, n56436,
         n56437, n56438, n56439, n56440, n56441, n56442, n56443, n56444,
         n56445, n56446, n56447, n56448, n56449, n56450, n56451, n56452,
         n56453, n56454, n56455, n56456, n56457, n56458, n56459, n56460,
         n56461, n56462, n56463, n56464, n56465, n56466, n56467, n56468,
         n56469, n56470, n56471, n56472, n56473, n56474, n56475, n56476,
         n56477, n56478, n56479, n56480, n56481, n56482, n56483, n56484,
         n56485, n56486, n56487, n56488, n56489, n56490, n56491, n56492,
         n56493, n56494, n56495, n56496, n56497, n56498, n56499, n56500,
         n56501, n56502, n56503, n56504, n56505, n56506, n56507, n56508,
         n56509, n56510, n56511, n56512, n56513, n56514, n56515, n56516,
         n56517, n56518, n56519, n56520, n56521, n56522, n56523, n56524,
         n56525, n56526, n56527, n56528, n56529, n56530, n56531, n56532,
         n56533, n56534, n56535, n56536, n56537, n56538, n56539, n56540,
         n56541, n56542, n56543, n56544, n56545, n56546, n56547, n56548,
         n56549, n56550, n56551, n56552, n56553, n56554, n56555, n56556,
         n56557, n56558, n56559, n56560, n56561, n56562, n56563, n56564,
         n56565, n56566, n56567, n56568, n56569, n56570, n56571, n56572,
         n56573, n56574, n56575, n56576, n56577, n56578, n56579, n56580,
         n56581, n56582, n56583, n56584, n56585, n56586, n56587, n56588,
         n56589, n56590, n56591, n56592, n56593, n56594, n56595, n56596,
         n56597, n56598, n56599, n56600, n56601, n56602, n56603, n56604,
         n56605, n56606, n56607, n56608, n56609, n56610, n56611, n56612,
         n56613, n56614, n56615, n56616, n56617, n56618, n56619, n56620,
         n56621, n56622, n56623, n56624, n56625, n56626, n56627, n56628,
         n56629, n56630, n56631, n56632, n56633, n56634, n56635, n56636,
         n56637, n56638, n56639, n56640, n56641, n56642, n56643, n56644,
         n56645, n56646, n56647, n56648, n56649, n56650, n56651, n56652,
         n56653, n56654, n56655, n56656, n56657, n56658, n56659, n56660,
         n56661, n56662, n56663, n56664, n56665, n56666, n56667, n56668,
         n56669, n56670, n56671, n56672, n56673, n56674, n56675, n56676,
         n56677, n56678, n56679, n56680, n56681, n56682, n56683, n56684,
         n56685, n56686, n56687, n56688, n56689, n56690, n56691, n56692,
         n56693, n56694, n56695, n56696, n56697, n56698, n56699, n56700,
         n56701, n56702, n56703, n56704, n56705, n56706, n56707, n56708,
         n56709, n56710, n56711, n56712, n56713, n56714, n56715, n56716,
         n56717, n56718, n56719, n56720, n56721, n56722, n56723, n56724,
         n56725, n56726, n56727, n56728, n56729, n56730, n56731, n56732,
         n56733, n56734, n56735, n56736, n56737, n56738, n56739, n56740,
         n56741, n56742, n56743, n56744, n56745, n56746, n56747, n56748,
         n56749, n56750, n56751, n56752, n56753, n56754, n56755, n56756,
         n56757, n56758, n56759, n56760, n56761, n56762, n56763, n56764,
         n56765, n56766, n56767, n56768, n56769, n56770, n56771, n56772,
         n56773, n56774, n56775, n56776, n56777, n56778, n56779, n56780,
         n56781, n56782, n56783, n56784, n56785, n56786, n56787, n56788,
         n56789, n56790, n56791, n56792, n56793, n56794, n56795, n56796,
         n56797, n56798, n56799, n56800, n56801, n56802, n56803, n56804,
         n56805, n56806, n56807, n56808, n56809, n56810, n56811, n56812,
         n56813, n56814, n56815, n56816, n56817, n56818, n56819, n56820,
         n56821, n56822, n56823, n56824, n56825, n56826, n56827, n56828,
         n56829, n56830, n56831, n56832, n56833, n56834, n56835, n56836,
         n56837, n56838, n56839, n56840, n56841, n56842, n56843, n56844,
         n56845, n56846, n56847, n56848, n56849, n56850, n56851, n56852,
         n56853, n56854, n56855, n56856, n56857, n56858, n56859, n56860,
         n56861, n56862, n56863, n56864, n56865, n56866, n56867, n56868,
         n56869, n56870, n56871, n56872, n56873, n56874, n56875, n56876,
         n56877, n56878, n56879, n56880, n56881, n56882, n56883, n56884,
         n56885, n56886, n56887, n56888, n56889, n56890, n56891, n56892,
         n56893, n56894, n56895, n56896, n56897, n56898, n56899, n56900,
         n56901, n56902, n56903, n56904, n56905, n56906, n56907, n56908,
         n56909, n56910, n56911, n56912, n56913, n56914, n56915, n56916,
         n56917, n56918, n56919, n56920, n56921, n56922, n56923, n56924,
         n56925, n56926, n56927, n56928, n56929, n56930, n56931, n56932,
         n56933, n56934, n56935, n56936, n56937, n56938, n56939, n56940,
         n56941, n56942, n56943, n56944, n56945, n56946, n56947, n56948,
         n56949, n56950, n56951, n56952, n56953, n56954, n56955, n56956,
         n56957, n56958, n56959, n56960, n56961, n56962, n56963, n56964,
         n56965, n56966, n56967, n56968, n56969, n56970, n56971, n56972,
         n56973, n56974, n56975, n56976, n56977, n56978, n56979, n56980,
         n56981, n56982, n56983, n56984, n56985, n56986, n56987, n56988,
         n56989, n56990, n56991, n56992, n56993, n56994, n56995, n56996,
         n56997, n56998, n56999, n57000, n57001, n57002, n57003, n57004,
         n57005, n57006, n57007, n57008, n57009, n57010, n57011, n57012,
         n57013, n57014, n57015, n57016, n57017, n57018, n57019, n57020,
         n57021, n57022, n57023, n57024, n57025, n57026, n57027, n57028,
         n57029, n57030, n57031, n57032, n57033, n57034, n57035, n57036,
         n57037, n57038, n57039, n57040, n57041, n57042, n57043, n57044,
         n57045, n57046, n57047, n57048, n57049, n57050, n57051, n57052,
         n57053, n57054, n57055, n57056, n57057, n57058, n57059, n57060,
         n57061, n57062, n57063, n57064, n57065, n57066, n57067, n57068,
         n57069, n57070, n57071, n57072, n57073, n57074, n57075, n57076,
         n57077, n57078, n57079, n57080, n57081, n57082, n57083, n57084,
         n57085, n57086, n57087, n57088, n57089, n57090, n57091, n57092,
         n57093, n57094, n57095, n57096, n57097, n57098, n57099, n57100,
         n57101, n57102, n57103, n57104, n57105, n57106, n57107, n57108,
         n57109, n57110, n57111, n57112, n57113, n57114, n57115, n57116,
         n57117, n57118, n57119, n57120, n57121, n57122, n57123, n57124,
         n57125, n57126, n57127, n57128, n57129, n57130, n57131, n57132,
         n57133, n57134, n57135, n57136, n57137, n57138, n57139, n57140,
         n57141, n57142, n57143, n57144, n57145, n57146, n57147, n57148,
         n57149, n57150, n57151, n57152, n57153, n57154, n57155, n57156,
         n57157, n57158, n57159, n57160, n57161, n57162, n57163, n57164,
         n57165, n57166, n57167, n57168, n57169, n57170, n57171, n57172,
         n57173, n57174, n57175, n57176, n57177, n57178, n57179, n57180,
         n57181, n57182, n57183, n57184, n57185, n57186, n57187, n57188,
         n57189, n57190, n57191, n57192, n57193, n57194, n57195, n57196,
         n57197, n57198, n57199, n57200, n57201, n57202, n57203, n57204,
         n57205, n57206, n57207, n57208, n57209, n57210, n57211, n57212,
         n57213, n57214, n57215, n57216, n57217, n57218, n57219, n57220,
         n57221, n57222, n57223, n57224, n57225, n57226, n57227, n57228,
         n57229, n57230, n57231, n57232, n57233, n57234, n57235, n57236,
         n57237, n57238, n57239, n57240, n57241, n57242, n57243, n57244,
         n57245, n57246, n57247, n57248, n57249, n57250, n57251, n57252,
         n57253, n57254, n57255, n57256, n57257, n57258, n57259, n57260,
         n57261, n57262, n57263, n57264, n57265, n57266, n57267, n57268,
         n57269, n57270, n57271, n57272, n57273, n57274, n57275, n57276,
         n57277, n57278, n57279, n57280, n57281, n57282, n57283, n57284,
         n57285, n57286, n57287, n57288, n57289, n57290, n57291, n57292,
         n57293, n57294, n57295, n57296, n57297, n57298, n57299, n57300,
         n57301, n57302, n57303, n57304, n57305, n57306, n57307, n57308,
         n57309, n57310, n57311, n57312, n57313, n57314, n57315, n57316,
         n57317, n57318, n57319, n57320, n57321, n57322, n57323, n57324,
         n57325, n57326, n57327, n57328, n57329, n57330, n57331, n57332,
         n57333, n57334, n57335, n57336, n57337, n57338, n57339, n57340,
         n57341, n57342, n57343, n57344, n57345, n57346, n57347, n57348,
         n57349, n57350, n57351, n57352, n57353, n57354, n57355, n57356,
         n57357, n57358, n57359, n57360, n57361, n57362, n57363, n57364,
         n57365, n57366, n57367, n57368, n57369, n57370, n57371, n57372,
         n57373, n57374, n57375, n57376, n57377, n57378, n57379, n57380,
         n57381, n57382, n57383, n57384, n57385, n57386, n57387, n57388,
         n57389, n57390, n57391, n57392, n57393, n57394, n57395, n57396,
         n57397, n57398, n57399, n57400, n57401, n57402, n57403, n57404,
         n57405, n57406, n57407, n57408, n57409, n57410, n57411, n57412,
         n57413, n57414, n57415, n57416, n57417, n57418, n57419, n57420,
         n57421, n57422, n57423, n57424, n57425, n57426, n57427, n57428,
         n57429, n57430, n57431, n57432, n57433, n57434, n57435, n57436,
         n57437, n57438, n57439, n57440, n57441, n57442, n57443, n57444,
         n57445, n57446, n57447, n57448, n57449, n57450, n57451, n57452,
         n57453, n57454, n57455, n57456, n57457, n57458, n57459, n57460,
         n57461, n57462, n57463, n57464, n57465, n57466, n57467, n57468,
         n57469, n57470, n57471, n57472, n57473, n57474, n57475, n57476,
         n57477, n57478, n57479, n57480, n57481, n57482, n57483, n57484,
         n57485, n57486, n57487, n57488, n57489, n57490, n57491, n57492,
         n57493, n57494, n57495, n57496, n57497, n57498, n57499, n57500,
         n57501, n57502, n57503, n57504, n57505, n57506, n57507, n57508,
         n57509, n57510, n57511, n57512, n57513, n57514, n57515, n57516,
         n57517, n57518, n57519, n57520, n57521, n57522, n57523, n57524,
         n57525, n57526, n57527, n57528, n57529, n57530, n57531, n57532,
         n57533, n57534, n57535, n57536, n57537, n57538, n57539, n57540,
         n57541, n57542, n57543, n57544, n57545, n57546, n57547, n57548,
         n57549, n57550, n57551, n57552, n57553, n57554, n57555, n57556,
         n57557, n57558, n57559, n57560, n57561, n57562, n57563, n57564,
         n57565, n57566, n57567, n57568, n57569, n57570, n57571, n57572,
         n57573, n57574, n57575, n57576, n57577, n57578, n57579, n57580,
         n57581, n57582, n57583, n57584, n57585, n57586, n57587, n57588,
         n57589, n57590, n57591, n57592, n57593, n57594, n57595, n57596,
         n57597, n57598, n57599, n57600, n57601, n57602, n57603, n57604,
         n57605, n57606, n57607, n57608, n57609, n57610, n57611, n57612,
         n57613, n57614, n57615, n57616, n57617, n57618, n57619, n57620,
         n57621, n57622, n57623, n57624, n57625, n57626, n57627, n57628,
         n57629, n57630, n57631, n57632, n57633, n57634, n57635, n57636,
         n57637, n57638, n57639, n57640, n57641, n57642, n57643, n57644,
         n57645, n57646, n57647, n57648, n57649, n57650, n57651, n57652,
         n57653, n57654, n57655, n57656, n57657, n57658, n57659, n57660,
         n57661, n57662, n57663, n57664, n57665, n57666, n57667, n57668,
         n57669, n57670, n57671, n57672, n57673, n57674, n57675, n57676,
         n57677, n57678, n57679, n57680, n57681, n57682, n57683, n57684,
         n57685, n57686, n57687, n57688, n57689, n57690, n57691, n57692,
         n57693, n57694, n57695, n57696, n57697, n57698, n57699, n57700,
         n57701, n57702, n57703, n57704, n57705, n57706, n57707, n57708,
         n57709, n57710, n57711, n57712, n57713, n57714, n57715, n57716,
         n57717, n57718, n57719, n57720, n57721, n57722, n57723, n57724,
         n57725, n57726, n57727, n57728, n57729, n57730, n57731, n57732,
         n57733, n57734, n57735, n57736, n57737, n57738, n57739, n57740,
         n57741, n57742, n57743, n57744, n57745, n57746, n57747, n57748,
         n57749, n57750, n57751, n57752, n57753, n57754, n57755, n57756,
         n57757, n57758, n57759, n57760, n57761, n57762, n57763, n57764,
         n57765, n57766, n57767, n57768, n57769, n57770, n57771, n57772,
         n57773, n57774, n57775, n57776, n57777, n57778, n57779, n57780,
         n57781, n57782, n57783, n57784, n57785, n57786, n57787, n57788,
         n57789, n57790, n57791, n57792, n57793, n57794, n57795, n57796,
         n57797, n57798, n57799, n57800, n57801, n57802, n57803, n57804,
         n57805, n57806, n57807, n57808, n57809, n57810, n57811, n57812,
         n57813, n57814, n57815, n57816, n57817, n57818, n57819, n57820,
         n57821, n57822, n57823, n57824, n57825, n57826, n57827, n57828,
         n57829, n57830, n57831, n57832, n57833, n57834, n57835, n57836,
         n57837, n57838, n57839, n57840, n57841, n57842, n57843, n57844,
         n57845, n57846, n57847, n57848, n57849, n57850, n57851, n57852,
         n57853, n57854, n57855, n57856, n57857, n57858, n57859, n57860,
         n57861, n57862, n57863, n57864, n57865, n57866, n57867, n57868,
         n57869, n57870, n57871, n57872, n57873, n57874, n57875, n57876,
         n57877, n57878, n57879, n57880, n57881, n57882, n57883, n57884,
         n57885, n57886, n57887, n57888, n57889, n57890, n57891, n57892,
         n57893, n57894, n57895, n57896, n57897, n57898, n57899, n57900,
         n57901, n57902, n57903, n57904, n57905, n57906, n57907, n57908,
         n57909, n57910, n57911, n57912, n57913, n57914, n57915, n57916,
         n57917, n57918, n57919, n57920, n57921, n57922, n57923, n57924,
         n57925, n57926, n57927, n57928, n57929, n57930, n57931, n57932,
         n57933, n57934, n57935, n57936, n57937, n57938, n57939, n57940,
         n57941, n57942, n57943, n57944, n57945, n57946, n57947, n57948,
         n57949, n57950, n57951, n57952, n57953, n57954, n57955, n57956,
         n57957, n57958, n57959, n57960, n57961, n57962, n57963, n57964,
         n57965, n57966, n57967, n57968, n57969, n57970, n57971, n57972,
         n57973, n57974, n57975, n57976, n57977, n57978, n57979, n57980,
         n57981, n57982, n57983, n57984, n57985, n57986, n57987, n57988,
         n57989, n57990, n57991, n57992, n57993, n57994, n57995, n57996,
         n57997, n57998, n57999, n58000, n58001, n58002, n58003, n58004,
         n58005, n58006, n58007, n58008, n58009, n58010, n58011, n58012,
         n58013, n58014, n58015, n58016, n58017, n58018, n58019, n58020,
         n58021, n58022, n58023, n58024, n58025, n58026, n58027, n58028,
         n58029, n58030, n58031, n58032, n58033, n58034, n58035, n58036,
         n58037, n58038, n58039, n58040, n58041, n58042, n58043, n58044,
         n58045, n58046, n58047, n58048, n58049, n58050, n58051, n58052,
         n58053, n58054, n58055, n58056, n58057, n58058, n58059, n58060,
         n58061, n58062, n58063, n58064, n58065, n58066, n58067, n58068,
         n58069, n58070, n58071, n58072, n58073, n58074, n58075, n58076,
         n58077, n58078, n58079, n58080, n58081, n58082, n58083, n58084,
         n58085, n58086, n58087, n58088, n58089, n58090, n58091, n58092,
         n58093, n58094, n58095, n58096, n58097, n58098, n58099, n58100,
         n58101, n58102, n58103, n58104, n58105, n58106, n58107, n58108,
         n58109, n58110, n58111, n58112, n58113, n58114, n58115, n58116,
         n58117, n58118, n58119, n58120, n58121, n58122, n58123, n58124,
         n58125, n58126, n58127, n58128, n58129, n58130, n58131, n58132,
         n58133, n58134, n58135, n58136, n58137, n58138, n58139, n58140,
         n58141, n58142, n58143, n58144, n58145, n58146, n58147, n58148,
         n58149, n58150, n58151, n58152, n58153, n58154, n58155, n58156,
         n58157, n58158, n58159, n58160, n58161, n58162, n58163, n58164,
         n58165, n58166, n58167, n58168, n58169, n58170, n58171, n58172,
         n58173, n58174, n58175, n58176, n58177, n58178, n58179, n58180,
         n58181, n58182, n58183, n58184, n58185, n58186, n58187, n58188,
         n58189, n58190, n58191, n58192, n58193, n58194, n58195, n58196,
         n58197, n58198, n58199, n58200, n58201, n58202, n58203, n58204,
         n58205, n58206, n58207, n58208, n58209, n58210, n58211, n58212,
         n58213, n58214, n58215, n58216, n58217, n58218, n58219, n58220,
         n58221, n58222, n58223, n58224, n58225, n58226, n58227, n58228,
         n58229, n58230, n58231, n58232, n58233, n58234, n58235, n58236,
         n58237, n58238, n58239, n58240, n58241, n58242, n58243, n58244,
         n58245, n58246, n58247, n58248, n58249, n58250, n58251, n58252,
         n58253, n58254, n58255, n58256, n58257, n58258, n58259, n58260,
         n58261, n58262, n58263, n58264, n58265, n58266, n58267, n58268,
         n58269, n58270, n58271, n58272, n58273, n58274, n58275, n58276,
         n58277, n58278, n58279, n58280, n58281, n58282, n58283, n58284,
         n58285, n58286, n58287, n58288, n58289, n58290, n58291, n58292,
         n58293, n58294, n58295, n58296, n58297, n58298, n58299, n58300,
         n58301, n58302, n58303, n58304, n58305, n58306, n58307, n58308,
         n58309, n58310, n58311, n58312, n58313, n58314, n58315, n58316,
         n58317, n58318, n58319, n58320, n58321, n58322, n58323, n58324,
         n58325, n58326, n58327, n58328, n58329, n58330, n58331, n58332,
         n58333, n58334, n58335, n58336, n58337, n58338, n58339, n58340,
         n58341, n58342, n58343, n58344, n58345, n58346, n58347, n58348,
         n58349, n58350, n58351, n58352, n58353, n58354, n58355, n58356,
         n58357, n58358, n58359, n58360, n58361, n58362, n58363, n58364,
         n58365, n58366, n58367, n58368, n58369, n58370, n58371, n58372,
         n58373, n58374, n58375, n58376, n58377, n58378, n58379, n58380,
         n58381, n58382, n58383, n58384, n58385, n58386, n58387, n58388,
         n58389, n58390, n58391, n58392, n58393, n58394, n58395, n58396,
         n58397, n58398, n58399, n58400, n58401, n58402, n58403, n58404,
         n58405, n58406, n58407, n58408, n58409, n58410, n58411, n58412,
         n58413, n58414, n58415, n58416, n58417, n58418, n58419, n58420,
         n58421, n58422, n58423, n58424, n58425, n58426, n58427, n58428,
         n58429, n58430, n58431, n58432, n58433, n58434, n58435, n58436,
         n58437, n58438, n58439, n58440, n58441, n58442, n58443, n58444,
         n58445, n58446, n58447, n58448, n58449, n58450, n58451, n58452,
         n58453, n58454, n58455, n58456, n58457, n58458, n58459, n58460,
         n58461, n58462, n58463, n58464, n58465, n58466, n58467, n58468,
         n58469, n58470, n58471, n58472, n58473, n58474, n58475, n58476,
         n58477, n58478, n58479, n58480, n58481, n58482, n58483, n58484,
         n58485, n58486, n58487, n58488, n58489, n58490, n58491, n58492,
         n58493, n58494, n58495, n58496, n58497, n58498, n58499, n58500,
         n58501, n58502, n58503, n58504, n58505, n58506, n58507, n58508,
         n58509, n58510, n58511, n58512, n58513, n58514, n58515, n58516,
         n58517, n58518, n58519, n58520, n58521, n58522, n58523, n58524,
         n58525, n58526, n58527, n58528, n58529, n58530, n58531, n58532,
         n58533, n58534, n58535, n58536, n58537, n58538, n58539, n58540,
         n58541, n58542, n58543, n58544, n58545, n58546, n58547, n58548,
         n58549, n58550, n58551, n58552, n58553, n58554, n58555, n58556,
         n58557, n58558, n58559, n58560, n58561, n58562, n58563, n58564,
         n58565, n58566, n58567, n58568, n58569, n58570, n58571, n58572,
         n58573, n58574, n58575, n58576, n58577, n58578, n58579, n58580,
         n58581, n58582, n58583, n58584, n58585, n58586, n58587, n58588,
         n58589, n58590, n58591, n58592, n58593, n58594, n58595, n58596,
         n58597, n58598, n58599, n58600, n58601, n58602, n58603, n58604,
         n58605, n58606, n58607, n58608, n58609, n58610, n58611, n58612,
         n58613, n58614, n58615, n58616, n58617, n58618, n58619, n58620,
         n58621, n58622, n58623, n58624, n58625, n58626, n58627, n58628,
         n58629, n58630, n58631, n58632, n58633, n58634, n58635, n58636,
         n58637, n58638, n58639, n58640, n58641, n58642, n58643, n58644,
         n58645, n58646, n58647, n58648, n58649, n58650, n58651, n58652,
         n58653, n58654, n58655, n58656, n58657, n58658, n58659, n58660,
         n58661, n58662, n58663, n58664, n58665, n58666, n58667, n58668,
         n58669, n58670, n58671, n58672, n58673, n58674, n58675, n58676,
         n58677, n58678, n58679, n58680, n58681, n58682, n58683, n58684,
         n58685, n58686, n58687, n58688, n58689, n58690, n58691, n58692,
         n58693, n58694, n58695, n58696, n58697, n58698, n58699, n58700,
         n58701, n58702, n58703, n58704, n58705, n58706, n58707, n58708,
         n58709, n58710, n58711, n58712, n58713, n58714, n58715, n58716,
         n58717, n58718, n58719, n58720, n58721, n58722, n58723, n58724,
         n58725, n58726, n58727, n58728, n58729, n58730, n58731, n58732,
         n58733, n58734, n58735, n58736, n58737, n58738, n58739, n58740,
         n58741, n58742, n58743, n58744, n58745, n58746, n58747, n58748,
         n58749, n58750, n58751, n58752, n58753, n58754, n58755, n58756,
         n58757, n58758, n58759, n58760, n58761, n58762, n58763, n58764,
         n58765, n58766, n58767, n58768, n58769, n58770, n58771, n58772,
         n58773, n58774, n58775, n58776, n58777, n58778, n58779, n58780,
         n58781, n58782, n58783, n58784, n58785, n58786, n58787, n58788,
         n58789, n58790, n58791, n58792, n58793, n58794, n58795, n58796,
         n58797, n58798, n58799, n58800, n58801, n58802, n58803, n58804,
         n58805, n58806, n58807, n58808, n58809, n58810, n58811, n58812,
         n58813, n58814, n58815, n58816, n58817, n58818, n58819, n58820,
         n58821, n58822, n58823, n58824, n58825, n58826, n58827, n58828,
         n58829, n58830, n58831, n58832, n58833, n58834, n58835, n58836,
         n58837, n58838, n58839, n58840, n58841, n58842, n58843, n58844,
         n58845, n58846, n58847, n58848, n58849, n58850, n58851, n58852,
         n58853, n58854, n58855, n58856, n58857, n58858, n58859, n58860,
         n58861, n58862, n58863, n58864, n58865, n58866, n58867, n58868,
         n58869, n58870, n58871, n58872, n58873, n58874, n58875, n58876,
         n58877, n58878, n58879, n58880, n58881, n58882, n58883, n58884,
         n58885, n58886, n58887, n58888, n58889, n58890, n58891, n58892,
         n58893, n58894, n58895, n58896, n58897, n58898, n58899, n58900,
         n58901, n58902, n58903, n58904, n58905, n58906, n58907, n58908,
         n58909, n58910, n58911, n58912, n58913, n58914, n58915, n58916,
         n58917, n58918, n58919, n58920, n58921, n58922, n58923, n58924,
         n58925, n58926, n58927, n58928, n58929, n58930, n58931, n58932,
         n58933, n58934, n58935, n58936, n58937, n58938, n58939, n58940,
         n58941, n58942, n58943, n58944, n58945, n58946, n58947, n58948,
         n58949, n58950, n58951, n58952, n58953, n58954, n58955, n58956,
         n58957, n58958, n58959, n58960, n58961, n58962, n58963, n58964,
         n58965, n58966, n58967, n58968, n58969, n58970, n58971, n58972,
         n58973, n58974, n58975, n58976, n58977, n58978, n58979, n58980,
         n58981, n58982, n58983, n58984, n58985, n58986, n58987, n58988,
         n58989, n58990, n58991, n58992, n58993, n58994, n58995, n58996,
         n58997, n58998, n58999, n59000, n59001, n59002, n59003, n59004,
         n59005, n59006, n59007, n59008, n59009, n59010, n59011, n59012,
         n59013, n59014, n59015, n59016, n59017, n59018, n59019, n59020,
         n59021, n59022, n59023, n59024, n59025, n59026, n59027, n59028,
         n59029, n59030, n59031, n59032, n59033, n59034, n59035, n59036,
         n59037, n59038, n59039, n59040, n59041, n59042, n59043, n59044,
         n59045, n59046, n59047, n59048, n59049, n59050, n59051, n59052,
         n59053, n59054, n59055, n59056, n59057, n59058, n59059, n59060,
         n59061, n59062, n59063, n59064, n59065, n59066, n59067, n59068,
         n59069, n59070, n59071, n59072, n59073, n59074, n59075, n59076,
         n59077, n59078, n59079, n59080, n59081, n59082, n59083, n59084,
         n59085, n59086, n59087, n59088, n59089, n59090, n59091, n59092,
         n59093, n59094, n59095, n59096, n59097, n59098, n59099, n59100,
         n59101, n59102, n59103, n59104, n59105, n59106, n59107, n59108,
         n59109, n59110, n59111, n59112, n59113, n59114, n59115, n59116,
         n59117, n59118, n59119, n59120, n59121, n59122, n59123, n59124,
         n59125, n59126, n59127, n59128, n59129, n59130, n59131, n59132,
         n59133, n59134, n59135, n59136, n59137, n59138, n59139, n59140,
         n59141, n59142, n59143, n59144, n59145, n59146, n59147, n59148,
         n59149, n59150, n59151, n59152, n59153, n59154, n59155, n59156,
         n59157, n59158, n59159, n59160, n59161, n59162, n59163, n59164,
         n59165, n59166, n59167, n59168, n59169, n59170, n59171, n59172,
         n59173, n59174, n59175, n59176, n59177, n59178, n59179, n59180,
         n59181, n59182, n59183, n59184, n59185, n59186, n59187, n59188,
         n59189, n59190, n59191, n59192, n59193, n59194, n59195, n59196,
         n59197, n59198, n59199, n59200, n59201, n59202, n59203, n59204,
         n59205, n59206, n59207, n59208, n59209, n59210, n59211, n59212,
         n59213, n59214, n59215, n59216, n59217, n59218, n59219, n59220,
         n59221, n59222, n59223, n59224, n59225, n59226, n59227, n59228,
         n59229, n59230, n59231, n59232, n59233, n59234, n59235, n59236,
         n59237, n59238, n59239, n59240, n59241, n59242, n59243, n59244,
         n59245, n59246, n59247, n59248, n59249, n59250, n59251, n59252,
         n59253, n59254, n59255, n59256, n59257, n59258, n59259, n59260,
         n59261, n59262, n59263, n59264, n59265, n59266, n59267, n59268,
         n59269, n59270, n59271, n59272, n59273, n59274, n59275, n59276,
         n59277, n59278, n59279, n59280, n59281, n59282, n59283, n59284,
         n59285, n59286, n59287, n59288, n59289, n59290, n59291, n59292,
         n59293, n59294, n59295, n59296, n59297, n59298, n59299, n59300,
         n59301, n59302, n59303, n59304, n59305, n59306, n59307, n59308,
         n59309, n59310, n59311, n59312, n59313, n59314, n59315, n59316,
         n59317, n59318, n59319, n59320, n59321, n59322, n59323, n59324,
         n59325, n59326, n59327, n59328, n59329, n59330, n59331, n59332,
         n59333, n59334, n59335, n59336, n59337, n59338, n59339, n59340,
         n59341, n59342, n59343, n59344, n59345, n59346, n59347, n59348,
         n59349, n59350, n59351, n59352, n59353, n59354, n59355, n59356,
         n59357, n59358, n59359, n59360, n59361, n59362, n59363, n59364,
         n59365, n59366, n59367, n59368, n59369, n59370, n59371, n59372,
         n59373, n59374, n59375, n59376, n59377, n59378, n59379, n59380,
         n59381, n59382, n59383, n59384, n59385, n59386, n59387, n59388,
         n59389, n59390, n59391, n59392, n59393, n59394, n59395, n59396,
         n59397, n59398, n59399, n59400, n59401, n59402, n59403, n59404,
         n59405, n59406, n59407, n59408, n59409, n59410, n59411, n59412,
         n59413, n59414, n59415, n59416, n59417, n59418, n59419, n59420,
         n59421, n59422, n59423, n59424, n59425, n59426, n59427, n59428,
         n59429, n59430, n59431, n59432, n59433, n59434, n59435, n59436,
         n59437, n59438, n59439, n59440, n59441, n59442, n59443, n59444,
         n59445, n59446, n59447, n59448, n59449, n59450, n59451, n59452,
         n59453, n59454, n59455, n59456, n59457, n59458, n59459, n59460,
         n59461, n59462, n59463, n59464, n59465, n59466, n59467, n59468,
         n59469, n59470, n59471, n59472, n59473, n59474, n59475, n59476,
         n59477, n59478, n59479, n59480, n59481, n59482, n59483, n59484,
         n59485, n59486, n59487, n59488, n59489, n59490, n59491, n59492,
         n59493, n59494, n59495, n59496, n59497, n59498, n59499, n59500,
         n59501, n59502, n59503, n59504, n59505, n59506, n59507, n59508,
         n59509, n59510, n59511, n59512, n59513, n59514, n59515, n59516,
         n59517, n59518, n59519, n59520, n59521, n59522, n59523, n59524,
         n59525, n59526, n59527, n59528, n59529, n59530, n59531, n59532,
         n59533, n59534, n59535, n59536, n59537, n59538, n59539, n59540,
         n59541, n59542, n59543, n59544, n59545, n59546, n59547, n59548,
         n59549, n59550, n59551, n59552, n59553, n59554, n59555, n59556,
         n59557, n59558, n59559, n59560, n59561, n59562, n59563, n59564,
         n59565, n59566, n59567, n59568, n59569, n59570, n59571, n59572,
         n59573, n59574, n59575, n59576, n59577, n59578, n59579, n59580,
         n59581, n59582, n59583, n59584, n59585, n59586, n59587, n59588,
         n59589, n59590, n59591, n59592, n59593, n59594, n59595, n59596,
         n59597, n59598, n59599, n59600, n59601, n59602, n59603, n59604,
         n59605, n59606, n59607, n59608, n59609, n59610, n59611, n59612,
         n59613, n59614, n59615, n59616, n59617, n59618, n59619, n59620,
         n59621, n59622, n59623, n59624, n59625, n59626, n59627, n59628,
         n59629, n59630, n59631, n59632, n59633, n59634, n59635, n59636,
         n59637, n59638, n59639, n59640, n59641, n59642, n59643, n59644,
         n59645, n59646, n59647, n59648, n59649, n59650, n59651, n59652,
         n59653, n59654, n59655, n59656, n59657, n59658, n59659, n59660,
         n59661, n59662, n59663, n59664, n59665, n59666, n59667, n59668,
         n59669, n59670, n59671, n59672, n59673, n59674, n59675, n59676,
         n59677, n59678, n59679, n59680, n59681, n59682, n59683, n59684,
         n59685, n59686, n59687, n59688, n59689, n59690, n59691, n59692,
         n59693, n59694, n59695, n59696, n59697, n59698, n59699, n59700,
         n59701, n59702, n59703, n59704, n59705, n59706, n59707, n59708,
         n59709, n59710, n59711, n59712, n59713, n59714, n59715, n59716,
         n59717, n59718, n59719, n59720, n59721, n59722, n59723, n59724,
         n59725, n59726, n59727, n59728, n59729, n59730, n59731, n59732,
         n59733, n59734, n59735, n59736, n59737, n59738, n59739, n59740,
         n59741, n59742, n59743, n59744, n59745, n59746, n59747, n59748,
         n59749, n59750, n59751, n59752, n59753, n59754, n59755, n59756,
         n59757, n59758, n59759, n59760, n59761, n59762, n59763, n59764,
         n59765, n59766, n59767, n59768, n59769, n59770, n59771, n59772,
         n59773, n59774, n59775, n59776, n59777, n59778, n59779, n59780,
         n59781, n59782, n59783, n59784, n59785, n59786, n59787, n59788,
         n59789, n59790, n59791, n59792, n59793, n59794, n59795, n59796,
         n59797, n59798, n59799, n59800, n59801, n59802, n59803, n59804,
         n59805, n59806, n59807, n59808, n59809, n59810, n59811, n59812,
         n59813, n59814, n59815, n59816, n59817, n59818, n59819, n59820,
         n59821, n59822, n59823, n59824, n59825, n59826, n59827, n59828,
         n59829, n59830, n59831, n59832, n59833, n59834, n59835, n59836,
         n59837, n59838, n59839, n59840, n59841, n59842, n59843, n59844,
         n59845, n59846, n59847, n59848, n59849, n59850, n59851, n59852,
         n59853, n59854, n59855, n59856, n59857, n59858, n59859, n59860,
         n59861, n59862, n59863, n59864, n59865, n59866, n59867, n59868,
         n59869, n59870, n59871, n59872, n59873, n59874, n59875, n59876,
         n59877, n59878, n59879, n59880, n59881, n59882, n59883, n59884,
         n59885, n59886, n59887, n59888, n59889, n59890, n59891, n59892,
         n59893, n59894, n59895, n59896, n59897, n59898, n59899, n59900,
         n59901, n59902, n59903, n59904, n59905, n59906, n59907, n59908,
         n59909, n59910, n59911, n59912, n59913, n59914, n59915, n59916,
         n59917, n59918, n59919, n59920, n59921, n59922, n59923, n59924,
         n59925, n59926, n59927, n59928, n59929, n59930, n59931, n59932,
         n59933, n59934, n59935, n59936, n59937, n59938, n59939, n59940,
         n59941, n59942, n59943, n59944, n59945, n59946, n59947, n59948,
         n59949, n59950, n59951, n59952, n59953, n59954, n59955, n59956,
         n59957, n59958, n59959, n59960, n59961, n59962, n59963, n59964,
         n59965, n59966, n59967, n59968, n59969, n59970, n59971, n59972,
         n59973, n59974, n59975, n59976, n59977, n59978, n59979, n59980,
         n59981, n59982, n59983, n59984, n59985, n59986, n59987, n59988,
         n59989, n59990, n59991, n59992, n59993, n59994, n59995, n59996,
         n59997, n59998, n59999, n60000, n60001, n60002, n60003, n60004,
         n60005, n60006, n60007, n60008, n60009, n60010, n60011, n60012,
         n60013, n60014, n60015, n60016, n60017, n60018, n60019, n60020,
         n60021, n60022, n60023, n60024, n60025, n60026, n60027, n60028,
         n60029, n60030, n60031, n60032, n60033, n60034, n60035, n60036,
         n60037, n60038, n60039, n60040, n60041, n60042, n60043, n60044,
         n60045, n60046, n60047, n60048, n60049, n60050, n60051, n60052,
         n60053, n60054, n60055, n60056, n60057, n60058, n60059, n60060,
         n60061, n60062, n60063, n60064, n60065, n60066, n60067, n60068,
         n60069, n60070, n60071, n60072, n60073, n60074, n60075, n60076,
         n60077, n60078, n60079, n60080, n60081, n60082, n60083, n60084,
         n60085, n60086, n60087, n60088, n60089, n60090, n60091, n60092,
         n60093, n60094, n60095, n60096, n60097, n60098, n60099, n60100,
         n60101, n60102, n60103, n60104, n60105, n60106, n60107, n60108,
         n60109, n60110, n60111, n60112, n60113, n60114, n60115, n60116,
         n60117, n60118, n60119, n60120, n60121, n60122, n60123, n60124,
         n60125, n60126, n60127, n60128, n60129, n60130, n60131, n60132,
         n60133, n60134, n60135, n60136, n60137, n60138, n60139, n60140,
         n60141, n60142, n60143, n60144, n60145, n60146, n60147, n60148,
         n60149, n60150, n60151, n60152, n60153, n60154, n60155, n60156,
         n60157, n60158, n60159, n60160, n60161, n60162, n60163, n60164,
         n60165, n60166, n60167, n60168, n60169, n60170, n60171, n60172,
         n60173, n60174, n60175, n60176, n60177, n60178, n60179, n60180,
         n60181, n60182, n60183, n60184, n60185, n60186, n60187, n60188,
         n60189, n60190, n60191, n60192, n60193, n60194, n60195, n60196,
         n60197, n60198, n60199, n60200, n60201, n60202, n60203, n60204,
         n60205, n60206, n60207, n60208, n60209, n60210, n60211, n60212,
         n60213, n60214, n60215, n60216, n60217, n60218, n60219, n60220,
         n60221, n60222, n60223, n60224, n60225, n60226, n60227, n60228,
         n60229, n60230, n60231, n60232, n60233, n60234, n60235, n60236,
         n60237, n60238, n60239, n60240, n60241, n60242, n60243, n60244,
         n60245, n60246, n60247, n60248, n60249, n60250, n60251, n60252,
         n60253, n60254, n60255, n60256, n60257, n60258, n60259, n60260,
         n60261, n60262, n60263, n60264, n60265, n60266, n60267, n60268,
         n60269, n60270, n60271, n60272, n60273, n60274, n60275, n60276,
         n60277, n60278, n60279, n60280, n60281, n60282, n60283, n60284,
         n60285, n60286, n60287, n60288, n60289, n60290, n60291, n60292,
         n60293, n60294, n60295, n60296, n60297, n60298, n60299, n60300,
         n60301, n60302, n60303, n60304, n60305, n60306, n60307, n60308,
         n60309, n60310, n60311, n60312, n60313, n60314, n60315, n60316,
         n60317, n60318, n60319, n60320, n60321, n60322, n60323, n60324,
         n60325, n60326, n60327, n60328, n60329, n60330, n60331, n60332,
         n60333, n60334, n60335, n60336, n60337, n60338, n60339, n60340,
         n60341, n60342, n60343, n60344, n60345, n60346, n60347, n60348,
         n60349, n60350, n60351, n60352, n60353, n60354, n60355, n60356,
         n60357, n60358, n60359, n60360, n60361, n60362, n60363, n60364,
         n60365, n60366, n60367, n60368, n60369, n60370, n60371, n60372,
         n60373, n60374, n60375, n60376, n60377, n60378, n60379, n60380,
         n60381, n60382, n60383, n60384, n60385, n60386, n60387, n60388,
         n60389, n60390, n60391, n60392, n60393, n60394, n60395, n60396,
         n60397, n60398, n60399, n60400, n60401, n60402, n60403, n60404,
         n60405, n60406, n60407, n60408, n60409, n60410, n60411, n60412,
         n60413, n60414, n60415, n60416, n60417, n60418, n60419, n60420,
         n60421, n60422, n60423, n60424, n60425, n60426, n60427, n60428,
         n60429, n60430, n60431, n60432, n60433, n60434, n60435, n60436,
         n60437, n60438, n60439, n60440, n60441, n60442, n60443, n60444,
         n60445, n60446, n60447, n60448, n60449, n60450, n60451, n60452,
         n60453, n60454, n60455, n60456, n60457, n60458, n60459, n60460,
         n60461, n60462, n60463, n60464, n60465, n60466, n60467, n60468,
         n60469, n60470, n60471, n60472, n60473, n60474, n60475, n60476,
         n60477, n60478, n60479, n60480, n60481, n60482, n60483, n60484,
         n60485, n60486, n60487, n60488, n60489, n60490, n60491, n60492,
         n60493, n60494, n60495, n60496, n60497, n60498, n60499, n60500,
         n60501, n60502, n60503, n60504, n60505, n60506, n60507, n60508,
         n60509, n60510, n60511, n60512, n60513, n60514, n60515, n60516,
         n60517, n60518, n60519, n60520, n60521, n60522, n60523, n60524,
         n60525, n60526, n60527, n60528, n60529, n60530, n60531, n60532,
         n60533, n60534, n60535, n60536, n60537, n60538, n60539, n60540,
         n60541, n60542, n60543, n60544, n60545, n60546, n60547, n60548,
         n60549, n60550, n60551, n60552, n60553, n60554, n60555, n60556,
         n60557, n60558, n60559, n60560, n60561, n60562, n60563, n60564,
         n60565, n60566, n60567, n60568, n60569, n60570, n60571, n60572,
         n60573, n60574, n60575, n60576, n60577, n60578, n60579, n60580,
         n60581, n60582, n60583, n60584, n60585, n60586, n60587, n60588,
         n60589, n60590, n60591, n60592, n60593, n60594, n60595, n60596,
         n60597, n60598, n60599, n60600, n60601, n60602, n60603, n60604,
         n60605, n60606, n60607, n60608, n60609, n60610, n60611, n60612,
         n60613, n60614, n60615, n60616, n60617, n60618, n60619, n60620,
         n60621, n60622, n60623, n60624, n60625, n60626, n60627, n60628,
         n60629, n60630, n60631, n60632, n60633, n60634, n60635, n60636,
         n60637, n60638, n60639, n60640, n60641, n60642, n60643, n60644,
         n60645, n60646, n60647, n60648, n60649, n60650, n60651, n60652,
         n60653, n60654, n60655, n60656, n60657, n60658, n60659, n60660,
         n60661, n60662, n60663, n60664, n60665, n60666, n60667, n60668,
         n60669, n60670, n60671, n60672, n60673, n60674, n60675, n60676,
         n60677, n60678, n60679, n60680, n60681, n60682, n60683, n60684,
         n60685, n60686, n60687, n60688, n60689, n60690, n60691, n60692,
         n60693, n60694, n60695, n60696, n60697, n60698, n60699, n60700,
         n60701, n60702, n60703, n60704, n60705, n60706, n60707, n60708,
         n60709, n60710, n60711, n60712, n60713, n60714, n60715, n60716,
         n60717, n60718, n60719, n60720, n60721, n60722, n60723, n60724,
         n60725, n60726, n60727, n60728, n60729, n60730, n60731, n60732,
         n60733, n60734, n60735, n60736, n60737, n60738, n60739, n60740,
         n60741, n60742, n60743, n60744, n60745, n60746, n60747, n60748,
         n60749, n60750, n60751, n60752, n60753, n60754, n60755, n60756,
         n60757, n60758, n60759, n60760, n60761, n60762, n60763, n60764,
         n60765, n60766, n60767, n60768, n60769, n60770, n60771, n60772,
         n60773, n60774, n60775, n60776, n60777, n60778, n60779, n60780,
         n60781, n60782, n60783, n60784, n60785, n60786, n60787, n60788,
         n60789, n60790, n60791, n60792, n60793, n60794, n60795, n60796,
         n60797, n60798, n60799, n60800, n60801, n60802, n60803, n60804,
         n60805, n60806, n60807, n60808, n60809, n60810, n60811, n60812,
         n60813, n60814, n60815, n60816, n60817, n60818, n60819, n60820,
         n60821, n60822, n60823, n60824, n60825, n60826, n60827, n60828,
         n60829, n60830, n60831, n60832, n60833, n60834, n60835, n60836,
         n60837, n60838, n60839, n60840, n60841, n60842, n60843, n60844,
         n60845, n60846, n60847, n60848, n60849, n60850, n60851, n60852,
         n60853, n60854, n60855, n60856, n60857, n60858, n60859, n60860,
         n60861, n60862, n60863, n60864, n60865, n60866, n60867, n60868,
         n60869, n60870, n60871, n60872, n60873, n60874, n60875, n60876,
         n60877, n60878, n60879, n60880, n60881, n60882, n60883, n60884,
         n60885, n60886, n60887, n60888, n60889, n60890, n60891, n60892,
         n60893, n60894, n60895, n60896, n60897, n60898, n60899, n60900,
         n60901, n60902, n60903, n60904, n60905, n60906, n60907, n60908,
         n60909, n60910, n60911, n60912, n60913, n60914, n60915, n60916,
         n60917, n60918, n60919, n60920, n60921, n60922, n60923, n60924,
         n60925, n60926, n60927, n60928, n60929, n60930, n60931, n60932,
         n60933, n60934, n60935, n60936, n60937, n60938, n60939, n60940,
         n60941, n60942, n60943, n60944, n60945, n60946, n60947, n60948,
         n60949, n60950, n60951, n60952, n60953, n60954, n60955, n60956,
         n60957, n60958, n60959, n60960, n60961, n60962, n60963, n60964,
         n60965, n60966, n60967, n60968, n60969, n60970, n60971, n60972,
         n60973, n60974, n60975, n60976, n60977, n60978, n60979, n60980,
         n60981, n60982, n60983, n60984, n60985, n60986, n60987, n60988,
         n60989, n60990, n60991, n60992, n60993, n60994, n60995, n60996,
         n60997, n60998, n60999, n61000, n61001, n61002, n61003, n61004,
         n61005, n61006, n61007, n61008, n61009, n61010, n61011, n61012,
         n61013, n61014, n61015, n61016, n61017, n61018, n61019, n61020,
         n61021, n61022, n61023, n61024, n61025, n61026, n61027, n61028,
         n61029, n61030, n61031, n61032, n61033, n61034, n61035, n61036,
         n61037, n61038, n61039, n61040, n61041, n61042, n61043, n61044,
         n61045, n61046, n61047, n61048, n61049, n61050, n61051, n61052,
         n61053, n61054, n61055, n61056, n61057, n61058, n61059, n61060,
         n61061, n61062, n61063, n61064, n61065, n61066, n61067, n61068,
         n61069, n61070, n61071, n61072, n61073, n61074, n61075, n61076,
         n61077, n61078, n61079, n61080, n61081, n61082, n61083, n61084,
         n61085, n61086, n61087, n61088, n61089, n61090, n61091, n61092,
         n61093, n61094, n61095, n61096, n61097, n61098, n61099, n61100,
         n61101, n61102, n61103, n61104, n61105, n61106, n61107, n61108,
         n61109, n61110, n61111, n61112, n61113, n61114, n61115, n61116,
         n61117, n61118, n61119, n61120, n61121, n61122, n61123, n61124,
         n61125, n61126, n61127, n61128, n61129, n61130, n61131, n61132,
         n61133, n61134, n61135, n61136, n61137, n61138, n61139, n61140,
         n61141, n61142, n61143, n61144, n61145, n61146, n61147, n61148,
         n61149, n61150, n61151, n61152, n61153, n61154, n61155, n61156,
         n61157, n61158, n61159, n61160, n61161, n61162, n61163, n61164,
         n61165, n61166, n61167, n61168, n61169, n61170, n61171, n61172,
         n61173, n61174, n61175, n61176, n61177, n61178, n61179, n61180,
         n61181, n61182, n61183, n61184, n61185, n61186, n61187, n61188,
         n61189, n61190, n61191, n61192, n61193, n61194, n61195, n61196,
         n61197, n61198, n61199, n61200, n61201, n61202, n61203, n61204,
         n61205, n61206, n61207, n61208, n61209, n61210, n61211, n61212,
         n61213, n61214, n61215, n61216, n61217, n61218, n61219, n61220,
         n61221, n61222, n61223, n61224, n61225, n61226, n61227, n61228,
         n61229, n61230, n61231, n61232, n61233, n61234, n61235, n61236,
         n61237, n61238, n61239, n61240, n61241, n61242, n61243, n61244,
         n61245, n61246, n61247, n61248, n61249, n61250, n61251, n61252,
         n61253, n61254, n61255, n61256, n61257, n61258, n61259, n61260,
         n61261, n61262, n61263, n61264, n61265, n61266, n61267, n61268,
         n61269, n61270, n61271, n61272, n61273, n61274, n61275, n61276,
         n61277, n61278, n61279, n61280, n61281, n61282, n61283, n61284,
         n61285, n61286, n61287, n61288, n61289, n61290, n61291, n61292,
         n61293, n61294, n61295, n61296, n61297, n61298, n61299, n61300,
         n61301, n61302, n61303, n61304, n61305, n61306, n61307, n61308,
         n61309, n61310, n61311, n61312, n61313, n61314, n61315, n61316,
         n61317, n61318, n61319, n61320, n61321, n61322, n61323, n61324,
         n61325, n61326, n61327, n61328, n61329, n61330, n61331, n61332,
         n61333, n61334, n61335, n61336, n61337, n61338, n61339, n61340,
         n61341, n61342, n61343, n61344, n61345, n61346, n61347, n61348,
         n61349, n61350, n61351, n61352, n61353, n61354, n61355, n61356,
         n61357, n61358, n61359, n61360, n61361, n61362, n61363, n61364,
         n61365, n61366, n61367, n61368, n61369, n61370, n61371, n61372,
         n61373, n61374, n61375, n61376, n61377, n61378, n61379, n61380,
         n61381, n61382, n61383, n61384, n61385, n61386, n61387, n61388,
         n61389, n61390, n61391, n61392, n61393, n61394, n61395, n61396,
         n61397, n61398, n61399, n61400, n61401, n61402, n61403, n61404,
         n61405, n61406, n61407, n61408, n61409, n61410, n61411, n61412,
         n61413, n61414, n61415, n61416, n61417, n61418, n61419, n61420,
         n61421, n61422, n61423, n61424, n61425, n61426, n61427, n61428,
         n61429, n61430, n61431, n61432, n61433, n61434, n61435, n61436,
         n61437, n61438, n61439, n61440, n61441, n61442, n61443, n61444,
         n61445, n61446, n61447, n61448, n61449, n61450, n61451, n61452,
         n61453, n61454, n61455, n61456, n61457, n61458, n61459, n61460,
         n61461, n61462, n61463, n61464, n61465, n61466, n61467, n61468,
         n61469, n61470, n61471, n61472, n61473, n61474, n61475, n61476,
         n61477, n61478, n61479, n61480, n61481, n61482, n61483, n61484,
         n61485, n61486, n61487, n61488, n61489, n61490, n61491, n61492,
         n61493, n61494, n61495, n61496, n61497, n61498, n61499, n61500,
         n61501, n61502, n61503, n61504, n61505, n61506, n61507, n61508,
         n61509, n61510, n61511, n61512, n61513, n61514, n61515, n61516,
         n61517, n61518, n61519, n61520, n61521, n61522, n61523, n61524,
         n61525, n61526, n61527, n61528, n61529, n61530, n61531, n61532,
         n61533, n61534, n61535, n61536, n61537, n61538, n61539, n61540,
         n61541, n61542, n61543, n61544, n61545, n61546, n61547, n61548,
         n61549, n61550, n61551, n61552, n61553, n61554, n61555, n61556,
         n61557, n61558, n61559, n61560, n61561, n61562, n61563, n61564,
         n61565, n61566, n61567, n61568, n61569, n61570, n61571, n61572,
         n61573, n61574, n61575, n61576, n61577, n61578, n61579, n61580,
         n61581, n61582, n61583, n61584, n61585, n61586, n61587, n61588,
         n61589, n61590, n61591, n61592, n61593, n61594, n61595, n61596,
         n61597, n61598, n61599, n61600, n61601, n61602, n61603, n61604,
         n61605, n61606, n61607, n61608, n61609, n61610, n61611, n61612,
         n61613, n61614, n61615, n61616, n61617, n61618, n61619, n61620,
         n61621, n61622, n61623, n61624, n61625, n61626, n61627, n61628,
         n61629, n61630, n61631, n61632, n61633, n61634, n61635, n61636,
         n61637, n61638, n61639, n61640, n61641, n61642, n61643, n61644,
         n61645, n61646, n61647, n61648, n61649, n61650, n61651, n61652,
         n61653, n61654, n61655, n61656, n61657, n61658, n61659, n61660,
         n61661, n61662, n61663, n61664, n61665, n61666, n61667, n61668,
         n61669, n61670, n61671, n61672, n61673, n61674, n61675, n61676,
         n61677, n61678, n61679, n61680, n61681, n61682, n61683, n61684,
         n61685, n61686, n61687, n61688, n61689, n61690, n61691, n61692,
         n61693, n61694, n61695, n61696, n61697, n61698, n61699, n61700,
         n61701, n61702, n61703, n61704, n61705, n61706, n61707, n61708,
         n61709, n61710, n61711, n61712, n61713, n61714, n61715, n61716,
         n61717, n61718, n61719, n61720, n61721, n61722, n61723, n61724,
         n61725, n61726, n61727, n61728, n61729, n61730, n61731, n61732,
         n61733, n61734, n61735, n61736, n61737, n61738, n61739, n61740,
         n61741, n61742, n61743, n61744, n61745, n61746, n61747, n61748,
         n61749, n61750, n61751, n61752, n61753, n61754, n61755, n61756,
         n61757, n61758, n61759, n61760, n61761, n61762, n61763, n61764,
         n61765, n61766, n61767, n61768, n61769, n61770, n61771, n61772,
         n61773, n61774, n61775, n61776, n61777, n61778, n61779, n61780,
         n61781, n61782, n61783, n61784, n61785, n61786, n61787, n61788,
         n61789, n61790, n61791, n61792, n61793, n61794, n61795, n61796,
         n61797, n61798, n61799, n61800, n61801, n61802, n61803, n61804,
         n61805, n61806, n61807, n61808, n61809, n61810, n61811, n61812,
         n61813, n61814, n61815, n61816, n61817, n61818, n61819, n61820,
         n61821, n61822, n61823, n61824, n61825, n61826, n61827, n61828,
         n61829, n61830, n61831, n61832, n61833, n61834, n61835, n61836,
         n61837, n61838, n61839, n61840, n61841, n61842, n61843, n61844,
         n61845, n61846, n61847, n61848, n61849, n61850, n61851, n61852,
         n61853, n61854, n61855, n61856, n61857, n61858, n61859, n61860,
         n61861, n61862, n61863, n61864, n61865, n61866, n61867, n61868,
         n61869, n61870, n61871, n61872, n61873, n61874, n61875, n61876,
         n61877, n61878, n61879, n61880, n61881, n61882, n61883, n61884,
         n61885, n61886, n61887, n61888, n61889, n61890, n61891, n61892,
         n61893, n61894, n61895, n61896, n61897, n61898, n61899, n61900,
         n61901, n61902, n61903, n61904, n61905, n61906, n61907, n61908,
         n61909, n61910, n61911, n61912, n61913, n61914, n61915, n61916,
         n61917, n61918, n61919, n61920, n61921, n61922, n61923, n61924,
         n61925, n61926, n61927, n61928, n61929, n61930, n61931, n61932,
         n61933, n61934, n61935, n61936, n61937, n61938, n61939, n61940,
         n61941, n61942, n61943, n61944, n61945, n61946, n61947, n61948,
         n61949, n61950, n61951, n61952, n61953, n61954, n61955, n61956,
         n61957, n61958, n61959, n61960, n61961, n61962, n61963, n61964,
         n61965, n61966, n61967, n61968, n61969, n61970, n61971, n61972,
         n61973, n61974, n61975, n61976, n61977, n61978, n61979, n61980,
         n61981, n61982, n61983, n61984, n61985, n61986, n61987, n61988,
         n61989, n61990, n61991, n61992, n61993, n61994, n61995, n61996,
         n61997, n61998, n61999, n62000, n62001, n62002, n62003, n62004,
         n62005, n62006, n62007, n62008, n62009, n62010, n62011, n62012,
         n62013, n62014, n62015, n62016, n62017, n62018, n62019, n62020,
         n62021, n62022, n62023, n62024, n62025, n62026, n62027, n62028,
         n62029, n62030, n62031, n62032, n62033, n62034, n62035, n62036,
         n62037, n62038, n62039, n62040, n62041, n62042, n62043, n62044,
         n62045, n62046, n62047, n62048, n62049, n62050, n62051, n62052,
         n62053, n62054, n62055, n62056, n62057, n62058, n62059, n62060,
         n62061, n62062, n62063, n62064, n62065, n62066, n62067, n62068,
         n62069, n62070, n62071, n62072, n62073, n62074, n62075, n62076,
         n62077, n62078, n62079, n62080, n62081, n62082, n62083, n62084,
         n62085, n62086, n62087, n62088, n62089, n62090, n62091, n62092,
         n62093, n62094, n62095, n62096, n62097, n62098, n62099, n62100,
         n62101, n62102, n62103, n62104, n62105, n62106, n62107, n62108,
         n62109, n62110, n62111, n62112, n62113, n62114, n62115, n62116,
         n62117, n62118, n62119, n62120, n62121, n62122, n62123, n62124,
         n62125, n62126, n62127, n62128, n62129, n62130, n62131, n62132,
         n62133, n62134, n62135, n62136, n62137, n62138, n62139, n62140,
         n62141, n62142, n62143, n62144, n62145, n62146, n62147, n62148,
         n62149, n62150, n62151, n62152, n62153, n62154, n62155, n62156,
         n62157, n62158, n62159, n62160, n62161, n62162, n62163, n62164,
         n62165, n62166, n62167, n62168, n62169, n62170, n62171, n62172,
         n62173, n62174, n62175, n62176, n62177, n62178, n62179, n62180,
         n62181, n62182, n62183, n62184, n62185, n62186, n62187, n62188,
         n62189, n62190, n62191, n62192, n62193, n62194, n62195, n62196,
         n62197, n62198, n62199, n62200, n62201, n62202, n62203, n62204,
         n62205, n62206, n62207, n62208, n62209, n62210, n62211, n62212,
         n62213, n62214, n62215, n62216, n62217, n62218, n62219, n62220,
         n62221, n62222, n62223, n62224, n62225, n62226, n62227, n62228,
         n62229, n62230, n62231, n62232, n62233, n62234, n62235, n62236,
         n62237, n62238, n62239, n62240, n62241, n62242, n62243, n62244,
         n62245, n62246, n62247, n62248, n62249, n62250, n62251, n62252,
         n62253, n62254, n62255, n62256, n62257, n62258, n62259, n62260,
         n62261, n62262, n62263, n62264, n62265, n62266, n62267, n62268,
         n62269, n62270, n62271, n62272, n62273, n62274, n62275, n62276,
         n62277, n62278, n62279, n62280, n62281, n62282, n62283, n62284,
         n62285, n62286, n62287, n62288, n62289, n62290, n62291, n62292,
         n62293, n62294, n62295, n62296, n62297, n62298, n62299, n62300,
         n62301, n62302, n62303, n62304, n62305, n62306, n62307, n62308,
         n62309, n62310, n62311, n62312, n62313, n62314, n62315, n62316,
         n62317, n62318, n62319, n62320, n62321, n62322, n62323, n62324,
         n62325, n62326, n62327, n62328, n62329, n62330, n62331, n62332,
         n62333, n62334, n62335, n62336, n62337, n62338, n62339, n62340,
         n62341, n62342, n62343, n62344, n62345, n62346, n62347, n62348,
         n62349, n62350, n62351, n62352, n62353, n62354, n62355, n62356,
         n62357, n62358, n62359, n62360, n62361, n62362, n62363, n62364,
         n62365, n62366, n62367, n62368, n62369, n62370, n62371, n62372,
         n62373, n62374, n62375, n62376, n62377, n62378, n62379, n62380,
         n62381, n62382, n62383, n62384, n62385, n62386, n62387, n62388,
         n62389, n62390, n62391, n62392, n62393, n62394, n62395, n62396,
         n62397, n62398, n62399, n62400, n62401, n62402, n62403, n62404,
         n62405, n62406, n62407, n62408, n62409, n62410, n62411, n62412,
         n62413, n62414, n62415, n62416, n62417, n62418, n62419, n62420,
         n62421, n62422, n62423, n62424, n62425, n62426, n62427, n62428,
         n62429, n62430, n62431, n62432, n62433, n62434, n62435, n62436,
         n62437, n62438, n62439, n62440, n62441, n62442, n62443, n62444,
         n62445, n62446, n62447, n62448, n62449, n62450, n62451, n62452,
         n62453, n62454, n62455, n62456, n62457, n62458, n62459, n62460,
         n62461, n62462, n62463, n62464, n62465, n62466, n62467, n62468,
         n62469, n62470, n62471, n62472, n62473, n62474, n62475, n62476,
         n62477, n62478, n62479, n62480, n62481, n62482, n62483, n62484,
         n62485, n62486, n62487, n62488, n62489, n62490, n62491, n62492,
         n62493, n62494, n62495, n62496, n62497, n62498, n62499, n62500,
         n62501, n62502, n62503, n62504, n62505, n62506, n62507, n62508,
         n62509, n62510, n62511, n62512, n62513, n62514, n62515, n62516,
         n62517, n62518, n62519, n62520, n62521, n62522, n62523, n62524,
         n62525, n62526, n62527, n62528, n62529, n62530, n62531, n62532,
         n62533, n62534, n62535, n62536, n62537, n62538, n62539, n62540,
         n62541, n62542, n62543, n62544, n62545, n62546, n62547, n62548,
         n62549, n62550, n62551, n62552, n62553, n62554, n62555, n62556,
         n62557, n62558, n62559, n62560, n62561, n62562, n62563, n62564,
         n62565, n62566, n62567, n62568, n62569, n62570, n62571, n62572,
         n62573, n62574, n62575, n62576, n62577, n62578, n62579, n62580,
         n62581, n62582, n62583, n62584, n62585, n62586, n62587, n62588,
         n62589, n62590, n62591, n62592, n62593, n62594, n62595, n62596,
         n62597, n62598, n62599, n62600, n62601, n62602, n62603, n62604,
         n62605, n62606, n62607, n62608, n62609, n62610, n62611, n62612,
         n62613, n62614, n62615, n62616, n62617, n62618, n62619, n62620,
         n62621, n62622, n62623, n62624, n62625, n62626, n62627, n62628,
         n62629, n62630, n62631, n62632, n62633, n62634, n62635, n62636,
         n62637, n62638, n62639, n62640, n62641, n62642, n62643, n62644,
         n62645, n62646, n62647, n62648, n62649, n62650, n62651, n62652,
         n62653, n62654, n62655, n62656, n62657, n62658, n62659, n62660,
         n62661, n62662, n62663, n62664, n62665, n62666, n62667, n62668,
         n62669, n62670, n62671, n62672, n62673, n62674, n62675, n62676,
         n62677, n62678, n62679, n62680, n62681, n62682, n62683, n62684,
         n62685, n62686, n62687, n62688, n62689, n62690, n62691, n62692,
         n62693, n62694, n62695, n62696, n62697, n62698, n62699, n62700,
         n62701, n62702, n62703, n62704, n62705, n62706, n62707, n62708,
         n62709, n62710, n62711, n62712, n62713, n62714, n62715, n62716,
         n62717, n62718, n62719, n62720, n62721, n62722, n62723, n62724,
         n62725, n62726, n62727, n62728, n62729, n62730, n62731, n62732,
         n62733, n62734, n62735, n62736, n62737, n62738, n62739, n62740,
         n62741, n62742, n62743, n62744, n62745, n62746, n62747, n62748,
         n62749, n62750, n62751, n62752, n62753, n62754, n62755, n62756,
         n62757, n62758, n62759, n62760, n62761, n62762, n62763, n62764,
         n62765, n62766, n62767, n62768, n62769, n62770, n62771, n62772,
         n62773, n62774, n62775, n62776, n62777, n62778, n62779, n62780,
         n62781, n62782, n62783, n62784, n62785, n62786, n62787, n62788,
         n62789, n62790, n62791, n62792, n62793, n62794, n62795, n62796,
         n62797, n62798, n62799, n62800, n62801, n62802, n62803, n62804,
         n62805, n62806, n62807, n62808, n62809, n62810, n62811, n62812,
         n62813, n62814, n62815, n62816, n62817, n62818, n62819, n62820,
         n62821, n62822, n62823, n62824, n62825, n62826, n62827, n62828,
         n62829, n62830, n62831, n62832, n62833, n62834, n62835, n62836,
         n62837, n62838, n62839, n62840, n62841, n62842, n62843, n62844,
         n62845, n62846, n62847, n62848, n62849, n62850, n62851, n62852,
         n62853, n62854, n62855, n62856, n62857, n62858, n62859, n62860,
         n62861, n62862, n62863, n62864, n62865, n62866, n62867, n62868,
         n62869, n62870, n62871, n62872, n62873, n62874, n62875, n62876,
         n62877, n62878, n62879, n62880, n62881, n62882, n62883, n62884,
         n62885, n62886, n62887, n62888, n62889, n62890, n62891, n62892,
         n62893, n62894, n62895, n62896, n62897, n62898, n62899, n62900,
         n62901, n62902, n62903, n62904, n62905, n62906, n62907, n62908,
         n62909, n62910, n62911, n62912, n62913, n62914, n62915, n62916,
         n62917, n62918, n62919, n62920, n62921, n62922, n62923, n62924,
         n62925, n62926, n62927, n62928, n62929, n62930, n62931, n62932,
         n62933, n62934, n62935, n62936, n62937, n62938, n62939, n62940,
         n62941, n62942, n62943, n62944, n62945, n62946, n62947, n62948,
         n62949, n62950, n62951, n62952, n62953, n62954, n62955, n62956,
         n62957, n62958, n62959, n62960, n62961, n62962, n62963, n62964,
         n62965, n62966, n62967, n62968, n62969, n62970, n62971, n62972,
         n62973, n62974, n62975, n62976, n62977, n62978, n62979, n62980,
         n62981, n62982, n62983, n62984, n62985, n62986, n62987, n62988,
         n62989, n62990, n62991, n62992, n62993, n62994, n62995, n62996,
         n62997, n62998, n62999, n63000, n63001, n63002, n63003, n63004,
         n63005, n63006, n63007, n63008, n63009, n63010, n63011, n63012,
         n63013, n63014, n63015, n63016, n63017, n63018, n63019, n63020,
         n63021, n63022, n63023, n63024, n63025, n63026, n63027, n63028,
         n63029, n63030, n63031, n63032, n63033, n63034, n63035, n63036,
         n63037, n63038, n63039, n63040, n63041, n63042, n63043, n63044,
         n63045, n63046, n63047, n63048, n63049, n63050, n63051, n63052,
         n63053, n63054, n63055, n63056, n63057, n63058, n63059, n63060,
         n63061, n63062, n63063, n63064, n63065, n63066, n63067, n63068,
         n63069, n63070, n63071, n63072, n63073, n63074, n63075, n63076,
         n63077, n63078, n63079, n63080, n63081, n63082, n63083, n63084,
         n63085, n63086, n63087, n63088, n63089, n63090, n63091, n63092,
         n63093, n63094, n63095, n63096, n63097, n63098, n63099, n63100,
         n63101, n63102, n63103, n63104, n63105, n63106, n63107, n63108,
         n63109, n63110, n63111, n63112, n63113, n63114, n63115, n63116,
         n63117, n63118, n63119, n63120, n63121, n63122, n63123, n63124,
         n63125, n63126, n63127, n63128, n63129, n63130, n63131, n63132,
         n63133, n63134, n63135, n63136, n63137, n63138, n63139, n63140,
         n63141, n63142, n63143, n63144, n63145, n63146, n63147, n63148,
         n63149, n63150, n63151, n63152, n63153, n63154, n63155, n63156,
         n63157, n63158, n63159, n63160, n63161, n63162, n63163, n63164,
         n63165, n63166, n63167, n63168, n63169, n63170, n63171, n63172,
         n63173, n63174, n63175, n63176, n63177, n63178, n63179, n63180,
         n63181, n63182, n63183, n63184, n63185, n63186, n63187, n63188,
         n63189, n63190, n63191, n63192, n63193, n63194, n63195, n63196,
         n63197, n63198, n63199, n63200, n63201, n63202, n63203, n63204,
         n63205, n63206, n63207, n63208, n63209, n63210, n63211, n63212,
         n63213, n63214, n63215, n63216, n63217, n63218, n63219, n63220,
         n63221, n63222, n63223, n63224, n63225, n63226, n63227, n63228,
         n63229, n63230, n63231, n63232, n63233, n63234, n63235, n63236,
         n63237, n63238, n63239, n63240, n63241, n63242, n63243, n63244,
         n63245, n63246, n63247, n63248, n63249, n63250, n63251, n63252,
         n63253, n63254, n63255, n63256, n63257, n63258, n63259, n63260,
         n63261, n63262, n63263, n63264, n63265, n63266, n63267, n63268,
         n63269, n63270, n63271, n63272, n63273, n63274, n63275, n63276,
         n63277, n63278, n63279, n63280, n63281, n63282, n63283, n63284,
         n63285, n63286, n63287, n63288, n63289, n63290, n63291, n63292,
         n63293, n63294, n63295, n63296, n63297, n63298, n63299, n63300,
         n63301, n63302, n63303, n63304, n63305, n63306, n63307, n63308,
         n63309, n63310, n63311, n63312, n63313, n63314, n63315, n63316,
         n63317, n63318, n63319, n63320, n63321, n63322, n63323, n63324,
         n63325, n63326, n63327, n63328, n63329, n63330, n63331, n63332,
         n63333, n63334, n63335, n63336, n63337, n63338, n63339, n63340,
         n63341, n63342, n63343, n63344, n63345, n63346, n63347, n63348,
         n63349, n63350, n63351, n63352, n63353, n63354, n63355, n63356,
         n63357, n63358, n63359, n63360, n63361, n63362, n63363, n63364,
         n63365, n63366, n63367, n63368, n63369, n63370, n63371, n63372,
         n63373, n63374, n63375, n63376, n63377, n63378, n63379, n63380,
         n63381, n63382, n63383, n63384, n63385, n63386, n63387, n63388,
         n63389, n63390, n63391, n63392, n63393, n63394, n63395, n63396,
         n63397, n63398, n63399, n63400, n63401, n63402, n63403, n63404,
         n63405, n63406, n63407, n63408, n63409, n63410, n63411, n63412,
         n63413, n63414, n63415, n63416, n63417, n63418, n63419, n63420,
         n63421, n63422, n63423, n63424, n63425, n63426, n63427, n63428,
         n63429, n63430, n63431, n63432, n63433, n63434, n63435, n63436,
         n63437, n63438, n63439, n63440, n63441, n63442, n63443, n63444,
         n63445, n63446, n63447, n63448, n63449, n63450, n63451, n63452,
         n63453, n63454, n63455, n63456, n63457, n63458, n63459, n63460,
         n63461, n63462, n63463, n63464, n63465, n63466, n63467, n63468,
         n63469, n63470, n63471, n63472, n63473, n63474, n63475, n63476,
         n63477, n63478, n63479, n63480, n63481, n63482, n63483, n63484,
         n63485, n63486, n63487, n63488, n63489, n63490, n63491, n63492,
         n63493, n63494, n63495, n63496, n63497, n63498, n63499, n63500,
         n63501, n63502, n63503, n63504, n63505, n63506, n63507, n63508,
         n63509, n63510, n63511, n63512, n63513, n63514, n63515, n63516,
         n63517, n63518, n63519, n63520, n63521, n63522, n63523, n63524,
         n63525, n63526, n63527, n63528, n63529, n63530, n63531, n63532,
         n63533, n63534, n63535, n63536, n63537, n63538, n63539, n63540,
         n63541, n63542, n63543, n63544, n63545, n63546, n63547, n63548,
         n63549, n63550, n63551, n63552, n63553, n63554, n63555, n63556,
         n63557, n63558, n63559, n63560, n63561, n63562, n63563, n63564,
         n63565, n63566, n63567, n63568, n63569, n63570, n63571, n63572,
         n63573, n63574, n63575, n63576, n63577, n63578, n63579, n63580,
         n63581, n63582, n63583, n63584, n63585, n63586, n63587, n63588,
         n63589, n63590, n63591, n63592, n63593, n63594, n63595, n63596,
         n63597, n63598, n63599, n63600, n63601, n63602, n63603, n63604,
         n63605, n63606, n63607, n63608, n63609, n63610, n63611, n63612,
         n63613, n63614, n63615, n63616, n63617, n63618, n63619, n63620,
         n63621, n63622, n63623, n63624, n63625, n63626, n63627, n63628,
         n63629, n63630, n63631, n63632, n63633, n63634, n63635, n63636,
         n63637, n63638, n63639, n63640, n63641, n63642, n63643, n63644,
         n63645, n63646, n63647, n63648, n63649, n63650, n63651, n63652,
         n63653, n63654, n63655, n63656, n63657, n63658, n63659, n63660,
         n63661, n63662, n63663, n63664, n63665, n63666, n63667, n63668,
         n63669, n63670, n63671, n63672, n63673, n63674, n63675, n63676,
         n63677, n63678, n63679, n63680, n63681, n63682, n63683, n63684,
         n63685, n63686, n63687, n63688, n63689, n63690, n63691, n63692,
         n63693, n63694, n63695, n63696, n63697, n63698, n63699, n63700,
         n63701, n63702, n63703, n63704, n63705, n63706, n63707, n63708,
         n63709, n63710, n63711, n63712, n63713, n63714, n63715, n63716,
         n63717, n63718, n63719, n63720, n63721, n63722, n63723, n63724,
         n63725, n63726, n63727, n63728, n63729, n63730, n63731, n63732,
         n63733, n63734, n63735, n63736, n63737, n63738, n63739, n63740,
         n63741, n63742, n63743, n63744, n63745, n63746, n63747, n63748,
         n63749, n63750, n63751, n63752, n63753, n63754, n63755, n63756,
         n63757, n63758, n63759, n63760, n63761, n63762, n63763, n63764,
         n63765, n63766, n63767, n63768, n63769, n63770, n63771, n63772,
         n63773, n63774, n63775, n63776, n63777, n63778, n63779, n63780,
         n63781, n63782, n63783, n63784, n63785, n63786, n63787, n63788,
         n63789, n63790, n63791, n63792, n63793, n63794, n63795, n63796,
         n63797, n63798, n63799, n63800, n63801, n63802, n63803, n63804,
         n63805, n63806, n63807, n63808, n63809, n63810, n63811, n63812,
         n63813, n63814, n63815, n63816, n63817, n63818, n63819, n63820,
         n63821, n63822, n63823, n63824, n63825, n63826, n63827, n63828,
         n63829, n63830, n63831, n63832, n63833, n63834, n63835, n63836,
         n63837, n63838, n63839, n63840, n63841, n63842, n63843, n63844,
         n63845, n63846, n63847, n63848, n63849, n63850, n63851, n63852,
         n63853, n63854, n63855, n63856, n63857, n63858, n63859, n63860,
         n63861, n63862, n63863, n63864, n63865, n63866, n63867, n63868,
         n63869, n63870, n63871, n63872, n63873, n63874, n63875, n63876,
         n63877, n63878, n63879, n63880, n63881, n63882, n63883, n63884,
         n63885, n63886, n63887, n63888, n63889, n63890, n63891, n63892,
         n63893, n63894, n63895, n63896, n63897, n63898, n63899, n63900,
         n63901, n63902, n63903, n63904, n63905, n63906, n63907, n63908,
         n63909, n63910, n63911, n63912, n63913, n63914, n63915, n63916,
         n63917, n63918, n63919, n63920, n63921, n63922, n63923, n63924,
         n63925, n63926, n63927, n63928, n63929, n63930, n63931, n63932,
         n63933, n63934, n63935, n63936, n63937, n63938, n63939, n63940,
         n63941, n63942, n63943, n63944, n63945, n63946, n63947, n63948,
         n63949, n63950, n63951, n63952, n63953, n63954, n63955, n63956,
         n63957, n63958, n63959, n63960, n63961, n63962, n63963, n63964,
         n63965, n63966, n63967, n63968, n63969, n63970, n63971, n63972,
         n63973, n63974, n63975, n63976, n63977, n63978, n63979, n63980,
         n63981, n63982, n63983, n63984, n63985, n63986, n63987, n63988,
         n63989, n63990, n63991, n63992, n63993, n63994, n63995, n63996,
         n63997, n63998, n63999, n64000, n64001, n64002, n64003, n64004,
         n64005, n64006, n64007, n64008, n64009, n64010, n64011, n64012,
         n64013, n64014, n64015, n64016, n64017, n64018, n64019, n64020,
         n64021, n64022, n64023, n64024, n64025, n64026, n64027, n64028,
         n64029, n64030, n64031, n64032, n64033, n64034, n64035, n64036,
         n64037, n64038, n64039, n64040, n64041, n64042, n64043, n64044,
         n64045, n64046, n64047, n64048, n64049, n64050, n64051, n64052,
         n64053, n64054, n64055, n64056, n64057, n64058, n64059, n64060,
         n64061, n64062, n64063, n64064, n64065, n64066, n64067, n64068,
         n64069, n64070, n64071, n64072, n64073, n64074, n64075, n64076,
         n64077, n64078, n64079, n64080, n64081, n64082, n64083, n64084,
         n64085, n64086, n64087, n64088, n64089, n64090, n64091, n64092,
         n64093, n64094, n64095, n64096, n64097, n64098, n64099, n64100,
         n64101, n64102, n64103, n64104, n64105, n64106, n64107, n64108,
         n64109, n64110, n64111, n64112, n64113, n64114, n64115, n64116,
         n64117, n64118, n64119, n64120, n64121, n64122, n64123, n64124,
         n64125, n64126, n64127, n64128, n64129, n64130, n64131, n64132,
         n64133, n64134, n64135, n64136, n64137, n64138, n64139, n64140,
         n64141, n64142, n64143, n64144, n64145, n64146, n64147, n64148,
         n64149, n64150, n64151, n64152, n64153, n64154, n64155, n64156,
         n64157, n64158, n64159, n64160, n64161, n64162, n64163, n64164,
         n64165, n64166, n64167, n64168, n64169, n64170, n64171, n64172,
         n64173, n64174, n64175, n64176, n64177, n64178, n64179, n64180,
         n64181, n64182, n64183, n64184, n64185, n64186, n64187, n64188,
         n64189, n64190, n64191, n64192, n64193, n64194, n64195, n64196,
         n64197, n64198, n64199, n64200, n64201, n64202, n64203, n64204,
         n64205, n64206, n64207, n64208, n64209, n64210, n64211, n64212,
         n64213, n64214, n64215, n64216, n64217, n64218, n64219, n64220,
         n64221, n64222, n64223, n64224, n64225, n64226, n64227, n64228,
         n64229, n64230, n64231, n64232, n64233, n64234, n64235, n64236,
         n64237, n64238, n64239, n64240, n64241, n64242, n64243, n64244,
         n64245, n64246, n64247, n64248, n64249, n64250, n64251, n64252,
         n64253, n64254, n64255, n64256, n64257, n64258, n64259, n64260,
         n64261, n64262, n64263, n64264, n64265, n64266, n64267, n64268,
         n64269, n64270, n64271, n64272, n64273, n64274, n64275, n64276,
         n64277, n64278, n64279, n64280, n64281, n64282, n64283, n64284,
         n64285, n64286, n64287, n64288, n64289, n64290, n64291, n64292,
         n64293, n64294, n64295, n64296, n64297, n64298, n64299, n64300,
         n64301, n64302, n64303, n64304, n64305, n64306, n64307, n64308,
         n64309, n64310, n64311, n64312, n64313, n64314, n64315, n64316,
         n64317, n64318, n64319, n64320, n64321, n64322, n64323, n64324,
         n64325, n64326, n64327, n64328, n64329, n64330, n64331, n64332,
         n64333, n64334, n64335, n64336, n64337, n64338, n64339, n64340,
         n64341, n64342, n64343, n64344, n64345, n64346, n64347, n64348,
         n64349, n64350, n64351, n64352, n64353, n64354, n64355, n64356,
         n64357, n64358, n64359, n64360, n64361, n64362, n64363, n64364,
         n64365, n64366, n64367, n64368, n64369, n64370, n64371, n64372,
         n64373, n64374, n64375, n64376, n64377, n64378, n64379, n64380,
         n64381, n64382, n64383, n64384, n64385, n64386, n64387, n64388,
         n64389, n64390, n64391, n64392, n64393, n64394, n64395, n64396,
         n64397, n64398, n64399, n64400, n64401, n64402, n64403, n64404,
         n64405, n64406, n64407, n64408, n64409, n64410, n64411, n64412,
         n64413, n64414, n64415, n64416, n64417, n64418, n64419, n64420,
         n64421, n64422, n64423, n64424, n64425, n64426, n64427, n64428,
         n64429, n64430, n64431, n64432, n64433, n64434, n64435, n64436,
         n64437, n64438, n64439, n64440, n64441, n64442, n64443, n64444,
         n64445, n64446, n64447, n64448, n64449, n64450, n64451, n64452,
         n64453, n64454, n64455, n64456, n64457, n64458, n64459, n64460,
         n64461, n64462, n64463, n64464, n64465, n64466, n64467, n64468,
         n64469, n64470, n64471, n64472, n64473, n64474, n64475, n64476,
         n64477, n64478, n64479, n64480, n64481, n64482, n64483, n64484,
         n64485, n64486, n64487, n64488, n64489, n64490, n64491, n64492,
         n64493, n64494, n64495, n64496, n64497, n64498, n64499, n64500,
         n64501, n64502, n64503, n64504, n64505, n64506, n64507, n64508,
         n64509, n64510, n64511, n64512, n64513, n64514, n64515, n64516,
         n64517, n64518, n64519, n64520, n64521, n64522, n64523, n64524,
         n64525, n64526, n64527, n64528, n64529, n64530, n64531, n64532,
         n64533, n64534, n64535, n64536, n64537, n64538, n64539, n64540,
         n64541, n64542, n64543, n64544, n64545, n64546, n64547, n64548,
         n64549, n64550, n64551, n64552, n64553, n64554, n64555, n64556,
         n64557, n64558, n64559, n64560, n64561, n64562, n64563, n64564,
         n64565, n64566, n64567, n64568, n64569, n64570, n64571, n64572,
         n64573, n64574, n64575, n64576, n64577, n64578, n64579, n64580,
         n64581, n64582, n64583, n64584, n64585, n64586, n64587, n64588,
         n64589, n64590, n64591, n64592, n64593, n64594, n64595, n64596,
         n64597, n64598, n64599, n64600, n64601, n64602, n64603, n64604,
         n64605, n64606, n64607, n64608, n64609, n64610, n64611, n64612,
         n64613, n64614, n64615, n64616, n64617, n64618, n64619, n64620,
         n64621, n64622, n64623, n64624, n64625, n64626, n64627, n64628,
         n64629, n64630, n64631, n64632, n64633, n64634, n64635, n64636,
         n64637, n64638, n64639, n64640, n64641, n64642, n64643, n64644,
         n64645, n64646, n64647, n64648, n64649, n64650, n64651, n64652,
         n64653, n64654, n64655, n64656, n64657, n64658, n64659, n64660,
         n64661, n64662, n64663, n64664, n64665, n64666, n64667, n64668,
         n64669, n64670, n64671, n64672, n64673, n64674, n64675, n64676,
         n64677, n64678, n64679, n64680, n64681, n64682, n64683, n64684,
         n64685, n64686, n64687, n64688, n64689, n64690, n64691, n64692,
         n64693, n64694, n64695, n64696, n64697, n64698, n64699, n64700,
         n64701, n64702, n64703, n64704, n64705, n64706, n64707, n64708,
         n64709, n64710, n64711, n64712, n64713, n64714, n64715, n64716,
         n64717, n64718, n64719, n64720, n64721, n64722, n64723, n64724,
         n64725, n64726, n64727, n64728, n64729, n64730, n64731, n64732,
         n64733, n64734, n64735, n64736, n64737, n64738, n64739, n64740,
         n64741, n64742, n64743, n64744, n64745, n64746, n64747, n64748,
         n64749, n64750, n64751, n64752, n64753, n64754, n64755, n64756,
         n64757, n64758, n64759, n64760, n64761, n64762, n64763, n64764,
         n64765, n64766, n64767, n64768, n64769, n64770, n64771, n64772,
         n64773, n64774, n64775, n64776, n64777, n64778, n64779, n64780,
         n64781, n64782, n64783, n64784, n64785, n64786, n64787, n64788,
         n64789, n64790, n64791, n64792, n64793, n64794, n64795, n64796,
         n64797, n64798, n64799, n64800, n64801, n64802, n64803, n64804,
         n64805, n64806, n64807, n64808, n64809, n64810, n64811, n64812,
         n64813, n64814, n64815, n64816, n64817, n64818, n64819, n64820,
         n64821, n64822, n64823, n64824, n64825, n64826, n64827, n64828,
         n64829, n64830, n64831, n64832, n64833, n64834, n64835, n64836,
         n64837, n64838, n64839, n64840, n64841, n64842, n64843, n64844,
         n64845, n64846, n64847, n64848, n64849, n64850, n64851, n64852,
         n64853, n64854, n64855, n64856, n64857, n64858, n64859, n64860,
         n64861, n64862, n64863, n64864, n64865, n64866, n64867, n64868,
         n64869, n64870, n64871, n64872, n64873, n64874, n64875, n64876,
         n64877, n64878, n64879, n64880, n64881, n64882, n64883, n64884,
         n64885, n64886, n64887, n64888, n64889, n64890, n64891, n64892,
         n64893, n64894, n64895, n64896, n64897, n64898, n64899, n64900,
         n64901, n64902, n64903, n64904, n64905, n64906, n64907, n64908,
         n64909, n64910, n64911, n64912, n64913, n64914, n64915, n64916,
         n64917, n64918, n64919, n64920, n64921, n64922, n64923, n64924,
         n64925, n64926, n64927, n64928, n64929, n64930, n64931, n64932,
         n64933, n64934, n64935, n64936, n64937, n64938, n64939, n64940,
         n64941, n64942, n64943, n64944, n64945, n64946, n64947, n64948,
         n64949, n64950, n64951, n64952, n64953, n64954, n64955, n64956,
         n64957, n64958, n64959, n64960, n64961, n64962, n64963, n64964,
         n64965, n64966, n64967, n64968, n64969, n64970, n64971, n64972,
         n64973, n64974, n64975, n64976, n64977, n64978, n64979, n64980,
         n64981, n64982, n64983, n64984, n64985, n64986, n64987, n64988,
         n64989, n64990, n64991, n64992, n64993, n64994, n64995, n64996,
         n64997, n64998, n64999, n65000, n65001, n65002, n65003, n65004,
         n65005, n65006, n65007, n65008, n65009, n65010, n65011, n65012,
         n65013, n65014, n65015, n65016, n65017, n65018, n65019, n65020,
         n65021, n65022, n65023, n65024, n65025, n65026, n65027, n65028,
         n65029, n65030, n65031, n65032, n65033, n65034, n65035, n65036,
         n65037, n65038, n65039, n65040, n65041, n65042, n65043, n65044,
         n65045, n65046, n65047, n65048, n65049, n65050, n65051, n65052,
         n65053, n65054, n65055, n65056, n65057, n65058, n65059, n65060,
         n65061, n65062, n65063, n65064, n65065, n65066, n65067, n65068,
         n65069, n65070, n65071, n65072, n65073, n65074, n65075, n65076,
         n65077, n65078, n65079, n65080, n65081, n65082, n65083, n65084,
         n65085, n65086, n65087, n65088, n65089, n65090, n65091, n65092,
         n65093, n65094, n65095, n65096, n65097, n65098, n65099, n65100,
         n65101, n65102, n65103, n65104, n65105, n65106, n65107, n65108,
         n65109, n65110, n65111, n65112, n65113, n65114, n65115, n65116,
         n65117, n65118, n65119, n65120, n65121, n65122, n65123, n65124,
         n65125, n65126, n65127, n65128, n65129, n65130, n65131, n65132,
         n65133, n65134, n65135, n65136, n65137, n65138, n65139, n65140,
         n65141, n65142, n65143, n65144, n65145, n65146, n65147, n65148,
         n65149, n65150, n65151, n65152, n65153, n65154, n65155, n65156,
         n65157, n65158, n65159, n65160, n65161, n65162, n65163, n65164,
         n65165, n65166, n65167, n65168, n65169, n65170, n65171, n65172,
         n65173, n65174, n65175, n65176, n65177, n65178, n65179, n65180,
         n65181, n65182, n65183, n65184, n65185, n65186, n65187, n65188,
         n65189, n65190, n65191, n65192, n65193, n65194, n65195, n65196,
         n65197, n65198, n65199, n65200, n65201, n65202, n65203, n65204,
         n65205, n65206, n65207, n65208, n65209, n65210, n65211, n65212,
         n65213, n65214, n65215, n65216, n65217, n65218, n65219, n65220,
         n65221, n65222, n65223, n65224, n65225, n65226, n65227, n65228,
         n65229, n65230, n65231, n65232, n65233, n65234, n65235, n65236,
         n65237, n65238, n65239, n65240, n65241, n65242, n65243, n65244,
         n65245, n65246, n65247, n65248, n65249, n65250, n65251, n65252,
         n65253, n65254, n65255, n65256, n65257, n65258, n65259, n65260,
         n65261, n65262, n65263, n65264, n65265, n65266, n65267, n65268,
         n65269, n65270, n65271, n65272, n65273, n65274, n65275, n65276,
         n65277, n65278, n65279, n65280, n65281, n65282, n65283, n65284,
         n65285, n65286, n65287, n65288, n65289, n65290, n65291, n65292,
         n65293, n65294, n65295, n65296, n65297, n65298, n65299, n65300,
         n65301, n65302, n65303, n65304, n65305, n65306, n65307, n65308,
         n65309, n65310, n65311, n65312, n65313, n65314, n65315, n65316,
         n65317, n65318, n65319, n65320, n65321, n65322, n65323, n65324,
         n65325, n65326, n65327, n65328, n65329, n65330, n65331, n65332,
         n65333, n65334, n65335, n65336, n65337, n65338, n65339, n65340,
         n65341, n65342, n65343, n65344, n65345, n65346, n65347, n65348,
         n65349, n65350, n65351, n65352, n65353, n65354, n65355, n65356,
         n65357, n65358, n65359, n65360, n65361, n65362, n65363, n65364,
         n65365, n65366, n65367, n65368, n65369, n65370, n65371, n65372,
         n65373, n65374, n65375, n65376, n65377, n65378, n65379, n65380,
         n65381, n65382, n65383, n65384, n65385, n65386, n65387, n65388,
         n65389, n65390, n65391, n65392, n65393, n65394, n65395, n65396,
         n65397, n65398, n65399, n65400, n65401, n65402, n65403, n65404,
         n65405, n65406, n65407, n65408, n65409, n65410, n65411, n65412,
         n65413, n65414, n65415, n65416, n65417, n65418, n65419, n65420,
         n65421, n65422, n65423, n65424, n65425, n65426, n65427, n65428,
         n65429, n65430, n65431, n65432, n65433, n65434, n65435, n65436,
         n65437, n65438, n65439, n65440, n65441, n65442, n65443, n65444,
         n65445, n65446, n65447, n65448, n65449, n65450, n65451, n65452,
         n65453, n65454, n65455, n65456, n65457, n65458, n65459, n65460,
         n65461, n65462, n65463, n65464, n65465, n65466, n65467, n65468,
         n65469, n65470, n65471, n65472, n65473, n65474, n65475, n65476,
         n65477, n65478, n65479, n65480, n65481, n65482, n65483, n65484,
         n65485, n65486, n65487, n65488, n65489, n65490, n65491, n65492,
         n65493, n65494, n65495, n65496, n65497, n65498, n65499, n65500,
         n65501, n65502, n65503, n65504, n65505, n65506, n65507, n65508,
         n65509, n65510, n65511, n65512, n65513, n65514, n65515, n65516,
         n65517, n65518, n65519, n65520, n65521, n65522, n65523, n65524,
         n65525, n65526, n65527, n65528, n65529, n65530, n65531, n65532,
         n65533, n65534, n65535, n65536, n65537, n65538, n65539, n65540,
         n65541, n65542, n65543, n65544, n65545, n65546, n65547, n65548,
         n65549, n65550, n65551, n65552, n65553, n65554, n65555, n65556,
         n65557, n65558, n65559, n65560, n65561, n65562, n65563, n65564,
         n65565, n65566, n65567, n65568, n65569, n65570, n65571, n65572,
         n65573, n65574, n65575, n65576, n65577, n65578, n65579, n65580,
         n65581, n65582, n65583, n65584, n65585, n65586, n65587, n65588,
         n65589, n65590, n65591, n65592, n65593, n65594, n65595, n65596,
         n65597, n65598, n65599, n65600, n65601, n65602, n65603, n65604,
         n65605, n65606, n65607, n65608, n65609, n65610, n65611, n65612,
         n65613, n65614, n65615, n65616, n65617, n65618, n65619, n65620,
         n65621, n65622, n65623, n65624, n65625, n65626, n65627, n65628,
         n65629, n65630, n65631, n65632, n65633, n65634, n65635, n65636,
         n65637, n65638, n65639, n65640, n65641, n65642, n65643, n65644,
         n65645, n65646, n65647, n65648, n65649, n65650, n65651, n65652,
         n65653, n65654, n65655, n65656, n65657, n65658, n65659, n65660,
         n65661, n65662, n65663, n65664, n65665, n65666, n65667, n65668,
         n65669, n65670, n65671, n65672, n65673, n65674, n65675, n65676,
         n65677, n65678, n65679, n65680, n65681, n65682, n65683, n65684,
         n65685, n65686, n65687, n65688, n65689, n65690, n65691, n65692,
         n65693, n65694, n65695, n65696, n65697, n65698, n65699, n65700,
         n65701, n65702, n65703, n65704, n65705, n65706, n65707, n65708,
         n65709, n65710, n65711, n65712, n65713, n65714, n65715, n65716,
         n65717, n65718, n65719, n65720, n65721, n65722, n65723, n65724,
         n65725, n65726, n65727, n65728, n65729, n65730, n65731, n65732,
         n65733, n65734, n65735, n65736, n65737, n65738, n65739, n65740,
         n65741, n65742, n65743, n65744, n65745, n65746, n65747, n65748,
         n65749, n65750, n65751, n65752, n65753, n65754, n65755, n65756,
         n65757, n65758, n65759, n65760, n65761, n65762, n65763, n65764,
         n65765, n65766, n65767, n65768, n65769, n65770, n65771, n65772,
         n65773, n65774, n65775, n65776, n65777, n65778, n65779, n65780,
         n65781, n65782, n65783, n65784, n65785, n65786, n65787, n65788,
         n65789, n65790, n65791, n65792, n65793, n65794, n65795, n65796,
         n65797, n65798, n65799, n65800, n65801, n65802, n65803, n65804,
         n65805, n65806, n65807, n65808, n65809, n65810, n65811, n65812,
         n65813, n65814, n65815, n65816, n65817, n65818, n65819, n65820,
         n65821, n65822, n65823, n65824, n65825, n65826, n65827, n65828,
         n65829, n65830, n65831, n65832, n65833, n65834, n65835, n65836,
         n65837, n65838, n65839, n65840, n65841, n65842, n65843, n65844,
         n65845, n65846, n65847, n65848, n65849, n65850, n65851, n65852,
         n65853, n65854, n65855, n65856, n65857, n65858, n65859, n65860,
         n65861, n65862, n65863, n65864, n65865, n65866, n65867, n65868,
         n65869, n65870, n65871, n65872, n65873, n65874, n65875, n65876,
         n65877, n65878, n65879, n65880, n65881, n65882, n65883, n65884,
         n65885, n65886, n65887, n65888, n65889, n65890, n65891, n65892,
         n65893, n65894, n65895, n65896, n65897, n65898, n65899, n65900,
         n65901, n65902, n65903, n65904, n65905, n65906, n65907, n65908,
         n65909, n65910, n65911, n65912, n65913, n65914, n65915, n65916,
         n65917, n65918, n65919, n65920, n65921, n65922, n65923, n65924,
         n65925, n65926, n65927, n65928, n65929, n65930, n65931, n65932,
         n65933, n65934, n65935, n65936, n65937, n65938, n65939, n65940,
         n65941, n65942, n65943, n65944, n65945, n65946, n65947, n65948,
         n65949, n65950, n65951, n65952, n65953, n65954, n65955, n65956,
         n65957, n65958, n65959, n65960, n65961, n65962, n65963, n65964,
         n65965, n65966, n65967, n65968, n65969, n65970, n65971, n65972,
         n65973, n65974, n65975, n65976, n65977, n65978, n65979, n65980,
         n65981, n65982, n65983, n65984, n65985, n65986, n65987, n65988,
         n65989, n65990, n65991, n65992, n65993, n65994, n65995, n65996,
         n65997, n65998, n65999, n66000, n66001, n66002, n66003, n66004,
         n66005, n66006, n66007, n66008, n66009, n66010, n66011, n66012,
         n66013, n66014, n66015, n66016, n66017, n66018, n66019, n66020,
         n66021, n66022, n66023, n66024, n66025, n66026, n66027, n66028,
         n66029, n66030, n66031, n66032, n66033, n66034, n66035, n66036,
         n66037, n66038, n66039, n66040, n66041, n66042, n66043, n66044,
         n66045, n66046, n66047, n66048, n66049, n66050, n66051, n66052,
         n66053, n66054, n66055, n66056, n66057, n66058, n66059, n66060,
         n66061, n66062, n66063, n66064, n66065, n66066, n66067, n66068,
         n66069, n66070, n66071, n66072, n66073, n66074, n66075, n66076,
         n66077, n66078, n66079, n66080, n66081, n66082, n66083, n66084,
         n66085, n66086, n66087, n66088, n66089, n66090, n66091, n66092,
         n66093, n66094, n66095, n66096, n66097, n66098, n66099, n66100,
         n66101, n66102, n66103, n66104, n66105, n66106, n66107, n66108,
         n66109, n66110, n66111, n66112, n66113, n66114, n66115, n66116,
         n66117, n66118, n66119, n66120, n66121, n66122, n66123, n66124,
         n66125, n66126, n66127, n66128, n66129, n66130, n66131, n66132,
         n66133, n66134, n66135, n66136, n66137, n66138, n66139, n66140,
         n66141, n66142, n66143, n66144, n66145, n66146, n66147, n66148,
         n66149, n66150, n66151, n66152, n66153, n66154, n66155, n66156,
         n66157, n66158, n66159, n66160, n66161, n66162, n66163, n66164,
         n66165, n66166, n66167, n66168, n66169, n66170, n66171, n66172,
         n66173, n66174, n66175, n66176, n66177, n66178, n66179, n66180,
         n66181, n66182, n66183, n66184, n66185, n66186, n66187, n66188,
         n66189, n66190, n66191, n66192, n66193, n66194, n66195, n66196,
         n66197, n66198, n66199, n66200, n66201, n66202, n66203, n66204,
         n66205, n66206, n66207, n66208, n66209, n66210, n66211, n66212,
         n66213, n66214, n66215, n66216, n66217, n66218, n66219, n66220,
         n66221, n66222, n66223, n66224, n66225, n66226, n66227, n66228,
         n66229, n66230, n66231, n66232, n66233, n66234, n66235, n66236,
         n66237, n66238, n66239, n66240, n66241, n66242, n66243, n66244,
         n66245, n66246, n66247, n66248, n66249, n66250, n66251, n66252,
         n66253, n66254, n66255, n66256, n66257, n66258, n66259, n66260,
         n66261, n66262, n66263, n66264, n66265, n66266, n66267, n66268,
         n66269, n66270, n66271, n66272, n66273, n66274, n66275, n66276,
         n66277, n66278, n66279, n66280, n66281, n66282, n66283, n66284,
         n66285, n66286, n66287, n66288, n66289, n66290, n66291, n66292,
         n66293, n66294, n66295, n66296, n66297, n66298, n66299, n66300,
         n66301, n66302, n66303, n66304, n66305, n66306, n66307, n66308,
         n66309, n66310, n66311, n66312, n66313, n66314, n66315, n66316,
         n66317, n66318, n66319, n66320, n66321, n66322, n66323, n66324,
         n66325, n66326, n66327, n66328, n66329, n66330, n66331, n66332,
         n66333, n66334, n66335, n66336, n66337, n66338, n66339, n66340,
         n66341, n66342, n66343, n66344, n66345, n66346, n66347, n66348,
         n66349, n66350, n66351, n66352, n66353, n66354, n66355, n66356,
         n66357, n66358, n66359, n66360, n66361, n66362, n66363, n66364,
         n66365, n66366, n66367, n66368, n66369, n66370, n66371, n66372,
         n66373, n66374, n66375, n66376, n66377, n66378, n66379, n66380,
         n66381, n66382, n66383, n66384, n66385, n66386, n66387, n66388,
         n66389, n66390, n66391, n66392, n66393, n66394, n66395, n66396,
         n66397, n66398, n66399, n66400, n66401, n66402, n66403, n66404,
         n66405, n66406, n66407, n66408, n66409, n66410, n66411, n66412,
         n66413, n66414, n66415, n66416, n66417, n66418, n66419, n66420,
         n66421, n66422, n66423, n66424, n66425, n66426, n66427, n66428,
         n66429, n66430, n66431, n66432, n66433, n66434, n66435, n66436,
         n66437, n66438, n66439, n66440, n66441, n66442, n66443, n66444,
         n66445, n66446, n66447, n66448, n66449, n66450, n66451, n66452,
         n66453, n66454, n66455, n66456, n66457, n66458, n66459, n66460,
         n66461, n66462, n66463, n66464, n66465, n66466, n66467, n66468,
         n66469, n66470, n66471, n66472, n66473, n66474, n66475, n66476,
         n66477, n66478, n66479, n66480, n66481, n66482, n66483, n66484,
         n66485, n66486, n66487, n66488, n66489, n66490, n66491, n66492,
         n66493, n66494, n66495, n66496, n66497, n66498, n66499, n66500,
         n66501, n66502, n66503, n66504, n66505, n66506, n66507, n66508,
         n66509, n66510, n66511, n66512, n66513, n66514, n66515, n66516,
         n66517, n66518, n66519, n66520, n66521, n66522, n66523, n66524,
         n66525, n66526, n66527, n66528, n66529, n66530, n66531, n66532,
         n66533, n66534, n66535, n66536, n66537, n66538, n66539, n66540,
         n66541, n66542, n66543, n66544, n66545, n66546, n66547, n66548,
         n66549, n66550, n66551, n66552, n66553, n66554, n66555, n66556,
         n66557, n66558, n66559, n66560, n66561, n66562, n66563, n66564,
         n66565, n66566, n66567, n66568, n66569, n66570, n66571, n66572,
         n66573, n66574, n66575, n66576, n66577, n66578, n66579, n66580,
         n66581, n66582, n66583, n66584, n66585, n66586, n66587, n66588,
         n66589, n66590, n66591, n66592, n66593, n66594, n66595, n66596,
         n66597, n66598, n66599, n66600, n66601, n66602, n66603, n66604,
         n66605, n66606, n66607, n66608, n66609, n66610, n66611, n66612,
         n66613, n66614, n66615, n66616, n66617, n66618, n66619, n66620,
         n66621, n66622, n66623, n66624, n66625, n66626, n66627, n66628,
         n66629, n66630, n66631, n66632, n66633, n66634, n66635, n66636,
         n66637, n66638, n66639, n66640, n66641, n66642, n66643, n66644,
         n66645, n66646, n66647, n66648, n66649, n66650, n66651, n66652,
         n66653, n66654, n66655, n66656, n66657, n66658, n66659, n66660,
         n66661, n66662, n66663, n66664, n66665, n66666, n66667, n66668,
         n66669, n66670, n66671, n66672, n66673, n66674, n66675, n66676,
         n66677, n66678, n66679, n66680, n66681, n66682, n66683, n66684,
         n66685, n66686, n66687, n66688, n66689, n66690, n66691, n66692,
         n66693, n66694, n66695, n66696, n66697, n66698, n66699, n66700,
         n66701, n66702, n66703, n66704, n66705, n66706, n66707, n66708,
         n66709, n66710, n66711, n66712, n66713, n66714, n66715, n66716,
         n66717, n66718, n66719, n66720, n66721, n66722, n66723, n66724,
         n66725, n66726, n66727, n66728, n66729, n66730, n66731, n66732,
         n66733, n66734, n66735, n66736, n66737, n66738, n66739, n66740,
         n66741, n66742, n66743, n66744, n66745, n66746, n66747, n66748,
         n66749, n66750, n66751, n66752, n66753, n66754, n66755, n66756,
         n66757, n66758, n66759, n66760, n66761, n66762, n66763, n66764,
         n66765, n66766, n66767, n66768, n66769, n66770, n66771, n66772,
         n66773, n66774, n66775, n66776, n66777, n66778, n66779, n66780,
         n66781, n66782, n66783, n66784, n66785, n66786, n66787, n66788,
         n66789, n66790, n66791, n66792, n66793, n66794, n66795, n66796,
         n66797, n66798, n66799, n66800, n66801, n66802, n66803, n66804,
         n66805, n66806, n66807, n66808, n66809, n66810, n66811, n66812,
         n66813, n66814, n66815, n66816, n66817, n66818, n66819, n66820,
         n66821, n66822, n66823, n66824, n66825, n66826, n66827, n66828,
         n66829, n66830, n66831, n66832, n66833, n66834, n66835, n66836,
         n66837, n66838, n66839, n66840, n66841, n66842, n66843, n66844,
         n66845, n66846, n66847, n66848, n66849, n66850, n66851, n66852,
         n66853, n66854, n66855, n66856, n66857, n66858, n66859, n66860,
         n66861, n66862, n66863, n66864, n66865, n66866, n66867, n66868,
         n66869, n66870, n66871, n66872, n66873, n66874, n66875, n66876,
         n66877, n66878, n66879, n66880, n66881, n66882, n66883, n66884,
         n66885, n66886, n66887, n66888, n66889, n66890, n66891, n66892,
         n66893, n66894, n66895, n66896, n66897, n66898, n66899, n66900,
         n66901, n66902, n66903, n66904, n66905, n66906, n66907, n66908,
         n66909, n66910, n66911, n66912, n66913, n66914, n66915, n66916,
         n66917, n66918, n66919, n66920, n66921, n66922, n66923, n66924,
         n66925, n66926, n66927, n66928, n66929, n66930, n66931, n66932,
         n66933, n66934, n66935, n66936, n66937, n66938, n66939, n66940,
         n66941, n66942, n66943, n66944, n66945, n66946, n66947, n66948,
         n66949, n66950, n66951, n66952, n66953, n66954, n66955, n66956,
         n66957, n66958, n66959, n66960, n66961, n66962, n66963, n66964,
         n66965, n66966, n66967, n66968, n66969, n66970, n66971, n66972,
         n66973, n66974, n66975, n66976, n66977, n66978, n66979, n66980,
         n66981, n66982, n66983, n66984, n66985, n66986, n66987, n66988,
         n66989, n66990, n66991, n66992, n66993, n66994, n66995, n66996,
         n66997, n66998, n66999, n67000, n67001, n67002, n67003, n67004,
         n67005, n67006, n67007, n67008, n67009, n67010, n67011, n67012,
         n67013, n67014, n67015, n67016, n67017, n67018, n67019, n67020,
         n67021, n67022, n67023, n67024, n67025, n67026, n67027, n67028,
         n67029, n67030, n67031, n67032, n67033, n67034, n67035, n67036,
         n67037, n67038, n67039, n67040, n67041, n67042, n67043, n67044,
         n67045, n67046, n67047, n67048, n67049, n67050, n67051, n67052,
         n67053, n67054, n67055, n67056, n67057, n67058, n67059, n67060,
         n67061, n67062, n67063, n67064, n67065, n67066, n67067, n67068,
         n67069, n67070, n67071, n67072, n67073, n67074, n67075, n67076,
         n67077, n67078, n67079, n67080, n67081, n67082, n67083, n67084,
         n67085, n67086, n67087, n67088, n67089, n67090, n67091, n67092,
         n67093, n67094, n67095, n67096, n67097, n67098, n67099, n67100,
         n67101, n67102, n67103, n67104, n67105, n67106, n67107, n67108,
         n67109, n67110, n67111, n67112, n67113, n67114, n67115, n67116,
         n67117, n67118, n67119, n67120, n67121, n67122, n67123, n67124,
         n67125, n67126, n67127, n67128, n67129, n67130, n67131, n67132,
         n67133, n67134, n67135, n67136, n67137, n67138, n67139, n67140,
         n67141, n67142, n67143, n67144, n67145, n67146, n67147, n67148,
         n67149, n67150, n67151, n67152, n67153, n67154, n67155, n67156,
         n67157, n67158, n67159, n67160, n67161, n67162, n67163, n67164,
         n67165, n67166, n67167, n67168, n67169, n67170, n67171, n67172,
         n67173, n67174, n67175, n67176, n67177, n67178, n67179, n67180,
         n67181, n67182, n67183, n67184, n67185, n67186, n67187, n67188,
         n67189, n67190, n67191, n67192, n67193, n67194, n67195, n67196,
         n67197, n67198, n67199, n67200, n67201, n67202, n67203, n67204,
         n67205, n67206, n67207, n67208, n67209, n67210, n67211, n67212,
         n67213, n67214, n67215, n67216, n67217, n67218, n67219, n67220,
         n67221, n67222, n67223, n67224, n67225, n67226, n67227, n67228,
         n67229, n67230, n67231, n67232, n67233, n67234, n67235, n67236,
         n67237, n67238, n67239, n67240, n67241, n67242, n67243, n67244,
         n67245, n67246, n67247, n67248, n67249, n67250, n67251, n67252,
         n67253, n67254, n67255, n67256, n67257, n67258, n67259, n67260,
         n67261, n67262, n67263, n67264, n67265, n67266, n67267, n67268,
         n67269, n67270, n67271, n67272, n67273, n67274, n67275, n67276,
         n67277, n67278, n67279, n67280, n67281, n67282, n67283, n67284,
         n67285, n67286, n67287, n67288, n67289, n67290, n67291, n67292,
         n67293, n67294, n67295, n67296, n67297, n67298, n67299, n67300,
         n67301, n67302, n67303, n67304, n67305, n67306, n67307, n67308,
         n67309, n67310, n67311, n67312, n67313, n67314, n67315, n67316,
         n67317, n67318, n67319, n67320, n67321, n67322, n67323, n67324,
         n67325, n67326, n67327, n67328, n67329, n67330, n67331, n67332,
         n67333, n67334, n67335, n67336, n67337, n67338, n67339, n67340,
         n67341, n67342, n67343, n67344, n67345, n67346, n67347, n67348,
         n67349, n67350, n67351, n67352, n67353, n67354, n67355, n67356,
         n67357, n67358, n67359, n67360, n67361, n67362, n67363, n67364,
         n67365, n67366, n67367, n67368, n67369, n67370, n67371, n67372,
         n67373, n67374, n67375, n67376, n67377, n67378, n67379, n67380,
         n67381, n67382, n67383, n67384, n67385, n67386, n67387, n67388,
         n67389, n67390, n67391, n67392, n67393, n67394, n67395, n67396,
         n67397, n67398, n67399, n67400, n67401, n67402, n67403, n67404,
         n67405, n67406, n67407, n67408, n67409, n67410, n67411, n67412,
         n67413, n67414, n67415, n67416, n67417, n67418, n67419, n67420,
         n67421, n67422, n67423, n67424, n67425, n67426, n67427, n67428,
         n67429, n67430, n67431, n67432, n67433, n67434, n67435, n67436,
         n67437, n67438, n67439, n67440, n67441, n67442, n67443, n67444,
         n67445, n67446, n67447, n67448, n67449, n67450, n67451, n67452,
         n67453, n67454, n67455, n67456, n67457, n67458, n67459, n67460,
         n67461, n67462, n67463, n67464, n67465, n67466, n67467, n67468,
         n67469, n67470, n67471, n67472, n67473, n67474, n67475, n67476,
         n67477, n67478, n67479, n67480, n67481, n67482, n67483, n67484,
         n67485, n67486, n67487, n67488, n67489, n67490, n67491, n67492,
         n67493, n67494, n67495, n67496, n67497, n67498, n67499, n67500,
         n67501, n67502, n67503, n67504, n67505, n67506, n67507, n67508,
         n67509, n67510, n67511, n67512, n67513, n67514, n67515, n67516,
         n67517, n67518, n67519, n67520, n67521, n67522, n67523, n67524,
         n67525, n67526, n67527, n67528, n67529, n67530, n67531, n67532,
         n67533, n67534, n67535, n67536, n67537, n67538, n67539, n67540,
         n67541, n67542, n67543, n67544, n67545, n67546, n67547, n67548,
         n67549, n67550, n67551, n67552, n67553, n67554, n67555, n67556,
         n67557, n67558, n67559, n67560, n67561, n67562, n67563, n67564,
         n67565, n67566, n67567, n67568, n67569, n67570, n67571, n67572,
         n67573, n67574, n67575, n67576, n67577, n67578, n67579, n67580,
         n67581, n67582, n67583, n67584, n67585, n67586, n67587, n67588,
         n67589, n67590, n67591, n67592, n67593, n67594, n67595, n67596,
         n67597, n67598, n67599, n67600, n67601, n67602, n67603, n67604,
         n67605, n67606, n67607, n67608, n67609, n67610, n67611, n67612,
         n67613, n67614, n67615, n67616, n67617, n67618, n67619, n67620,
         n67621, n67622, n67623, n67624, n67625, n67626, n67627, n67628,
         n67629, n67630, n67631, n67632, n67633, n67634, n67635, n67636,
         n67637, n67638, n67639, n67640, n67641, n67642, n67643, n67644,
         n67645, n67646, n67647, n67648, n67649, n67650, n67651, n67652,
         n67653, n67654, n67655, n67656, n67657, n67658, n67659, n67660,
         n67661, n67662, n67663, n67664, n67665, n67666, n67667, n67668,
         n67669, n67670, n67671, n67672, n67673, n67674, n67675, n67676,
         n67677, n67678, n67679, n67680, n67681, n67682, n67683, n67684,
         n67685, n67686, n67687, n67688, n67689, n67690, n67691, n67692,
         n67693, n67694, n67695, n67696, n67697, n67698, n67699, n67700,
         n67701, n67702, n67703, n67704, n67705, n67706, n67707, n67708,
         n67709, n67710, n67711, n67712, n67713, n67714, n67715, n67716,
         n67717, n67718, n67719, n67720, n67721, n67722, n67723, n67724,
         n67725, n67726, n67727, n67728, n67729, n67730, n67731, n67732,
         n67733, n67734, n67735, n67736, n67737, n67738, n67739, n67740,
         n67741, n67742, n67743, n67744, n67745, n67746, n67747, n67748,
         n67749, n67750, n67751, n67752, n67753, n67754, n67755, n67756,
         n67757, n67758, n67759, n67760, n67761, n67762, n67763, n67764,
         n67765, n67766, n67767, n67768, n67769, n67770, n67771, n67772,
         n67773, n67774, n67775, n67776, n67777, n67778, n67779, n67780,
         n67781, n67782, n67783, n67784, n67785, n67786, n67787, n67788,
         n67789, n67790, n67791, n67792, n67793, n67794, n67795, n67796,
         n67797, n67798, n67799, n67800, n67801, n67802, n67803, n67804,
         n67805, n67806, n67807, n67808, n67809, n67810, n67811, n67812,
         n67813, n67814, n67815, n67816, n67817, n67818, n67819, n67820,
         n67821, n67822, n67823, n67824, n67825, n67826, n67827, n67828,
         n67829, n67830, n67831, n67832, n67833, n67834, n67835, n67836,
         n67837, n67838, n67839, n67840, n67841, n67842, n67843, n67844,
         n67845, n67846, n67847, n67848, n67849, n67850, n67851, n67852,
         n67853, n67854, n67855, n67856, n67857, n67858, n67859, n67860,
         n67861, n67862, n67863, n67864, n67865, n67866, n67867, n67868,
         n67869, n67870, n67871, n67872, n67873, n67874, n67875, n67876,
         n67877, n67878, n67879, n67880, n67881, n67882, n67883, n67884,
         n67885, n67886, n67887, n67888, n67889, n67890, n67891, n67892,
         n67893, n67894, n67895, n67896, n67897, n67898, n67899, n67900,
         n67901, n67902, n67903, n67904, n67905, n67906, n67907, n67908,
         n67909, n67910, n67911, n67912, n67913, n67914, n67915, n67916,
         n67917, n67918, n67919, n67920, n67921, n67922, n67923, n67924,
         n67925, n67926, n67927, n67928, n67929, n67930, n67931, n67932,
         n67933, n67934, n67935, n67936, n67937, n67938, n67939, n67940,
         n67941, n67942, n67943, n67944, n67945, n67946, n67947, n67948,
         n67949, n67950, n67951, n67952, n67953, n67954, n67955, n67956,
         n67957, n67958, n67959, n67960, n67961, n67962, n67963, n67964,
         n67965, n67966, n67967, n67968, n67969, n67970, n67971, n67972,
         n67973, n67974, n67975, n67976, n67977, n67978, n67979, n67980,
         n67981, n67982, n67983, n67984, n67985, n67986, n67987, n67988,
         n67989, n67990, n67991, n67992, n67993, n67994, n67995, n67996,
         n67997, n67998, n67999, n68000, n68001, n68002, n68003, n68004,
         n68005, n68006, n68007, n68008, n68009, n68010, n68011, n68012,
         n68013, n68014, n68015, n68016, n68017, n68018, n68019, n68020,
         n68021, n68022, n68023, n68024, n68025, n68026, n68027, n68028,
         n68029, n68030, n68031, n68032, n68033, n68034, n68035, n68036,
         n68037, n68038, n68039, n68040, n68041, n68042, n68043, n68044,
         n68045, n68046, n68047, n68048, n68049, n68050, n68051, n68052,
         n68053, n68054, n68055, n68056, n68057, n68058, n68059, n68060,
         n68061, n68062, n68063, n68064, n68065, n68066, n68067, n68068,
         n68069, n68070, n68071, n68072, n68073, n68074, n68075, n68076,
         n68077, n68078, n68079, n68080, n68081, n68082, n68083, n68084,
         n68085, n68086, n68087, n68088, n68089, n68090, n68091, n68092,
         n68093, n68094, n68095, n68096, n68097, n68098, n68099, n68100,
         n68101, n68102, n68103, n68104, n68105, n68106, n68107, n68108,
         n68109, n68110, n68111, n68112, n68113, n68114, n68115, n68116,
         n68117, n68118, n68119, n68120, n68121, n68122, n68123, n68124,
         n68125, n68126, n68127, n68128, n68129, n68130, n68131, n68132,
         n68133, n68134, n68135, n68136, n68137, n68138, n68139, n68140,
         n68141, n68142, n68143, n68144, n68145, n68146, n68147, n68148,
         n68149, n68150, n68151, n68152, n68153, n68154, n68155, n68156,
         n68157, n68158, n68159, n68160, n68161, n68162, n68163, n68164,
         n68165, n68166, n68167, n68168, n68169, n68170, n68171, n68172,
         n68173, n68174, n68175, n68176, n68177, n68178, n68179, n68180,
         n68181, n68182, n68183, n68184, n68185, n68186, n68187, n68188,
         n68189, n68190, n68191, n68192, n68193, n68194, n68195, n68196,
         n68197, n68198, n68199, n68200, n68201, n68202, n68203, n68204,
         n68205, n68206, n68207, n68208, n68209, n68210, n68211, n68212,
         n68213, n68214, n68215, n68216, n68217, n68218, n68219, n68220,
         n68221, n68222, n68223, n68224, n68225, n68226, n68227, n68228,
         n68229, n68230, n68231, n68232, n68233, n68234, n68235, n68236,
         n68237, n68238, n68239, n68240, n68241, n68242, n68243, n68244,
         n68245, n68246, n68247, n68248, n68249, n68250, n68251, n68252,
         n68253, n68254, n68255, n68256, n68257, n68258, n68259, n68260,
         n68261, n68262, n68263, n68264, n68265, n68266, n68267, n68268,
         n68269, n68270, n68271, n68272, n68273, n68274, n68275, n68276,
         n68277, n68278, n68279, n68280, n68281, n68282, n68283, n68284,
         n68285, n68286, n68287, n68288, n68289, n68290, n68291, n68292,
         n68293, n68294, n68295, n68296, n68297, n68298, n68299, n68300,
         n68301, n68302, n68303, n68304, n68305, n68306, n68307, n68308,
         n68309, n68310, n68311, n68312, n68313, n68314, n68315, n68316,
         n68317, n68318, n68319, n68320, n68321, n68322, n68323, n68324,
         n68325, n68326, n68327, n68328, n68329, n68330, n68331, n68332,
         n68333, n68334, n68335, n68336, n68337, n68338, n68339, n68340,
         n68341, n68342, n68343, n68344, n68345, n68346, n68347, n68348,
         n68349, n68350, n68351, n68352, n68353, n68354, n68355, n68356,
         n68357, n68358, n68359, n68360, n68361, n68362, n68363, n68364,
         n68365, n68366, n68367, n68368, n68369, n68370, n68371, n68372,
         n68373, n68374, n68375, n68376, n68377, n68378, n68379, n68380,
         n68381, n68382, n68383, n68384, n68385, n68386, n68387, n68388,
         n68389, n68390, n68391, n68392, n68393, n68394, n68395, n68396,
         n68397, n68398, n68399, n68400, n68401, n68402, n68403, n68404,
         n68405, n68406, n68407, n68408, n68409, n68410, n68411, n68412,
         n68413, n68414, n68415, n68416, n68417, n68418, n68419, n68420,
         n68421, n68422, n68423, n68424, n68425, n68426, n68427, n68428,
         n68429, n68430, n68431, n68432, n68433, n68434, n68435, n68436,
         n68437, n68438, n68439, n68440, n68441, n68442, n68443, n68444,
         n68445, n68446, n68447, n68448, n68449, n68450, n68451, n68452,
         n68453, n68454, n68455, n68456, n68457, n68458, n68459, n68460,
         n68461, n68462, n68463, n68464, n68465, n68466, n68467, n68468,
         n68469, n68470, n68471, n68472, n68473, n68474, n68475, n68476,
         n68477, n68478, n68479, n68480, n68481, n68482, n68483, n68484,
         n68485, n68486, n68487, n68488, n68489, n68490, n68491, n68492,
         n68493, n68494, n68495, n68496, n68497, n68498, n68499, n68500,
         n68501, n68502, n68503, n68504, n68505, n68506, n68507, n68508,
         n68509, n68510, n68511, n68512, n68513, n68514, n68515, n68516,
         n68517, n68518, n68519, n68520, n68521, n68522, n68523, n68524,
         n68525, n68526, n68527, n68528, n68529, n68530, n68531, n68532,
         n68533, n68534, n68535, n68536, n68537, n68538, n68539, n68540,
         n68541, n68542, n68543, n68544, n68545, n68546, n68547, n68548,
         n68549, n68550, n68551, n68552, n68553, n68554, n68555, n68556,
         n68557, n68558, n68559, n68560, n68561, n68562, n68563, n68564,
         n68565, n68566, n68567, n68568, n68569, n68570, n68571, n68572,
         n68573, n68574, n68575, n68576, n68577, n68578, n68579, n68580,
         n68581, n68582, n68583, n68584, n68585, n68586, n68587, n68588,
         n68589, n68590, n68591, n68592, n68593, n68594, n68595, n68596,
         n68597, n68598, n68599, n68600, n68601, n68602, n68603, n68604,
         n68605, n68606, n68607, n68608, n68609, n68610, n68611, n68612,
         n68613, n68614, n68615, n68616, n68617, n68618, n68619, n68620,
         n68621, n68622, n68623, n68624, n68625, n68626, n68627, n68628,
         n68629, n68630, n68631, n68632, n68633, n68634, n68635, n68636,
         n68637, n68638, n68639, n68640, n68641, n68642, n68643, n68644,
         n68645, n68646, n68647, n68648, n68649, n68650, n68651, n68652,
         n68653, n68654, n68655, n68656, n68657, n68658, n68659, n68660,
         n68661, n68662, n68663, n68664, n68665, n68666, n68667, n68668,
         n68669, n68670, n68671, n68672, n68673, n68674, n68675, n68676,
         n68677, n68678, n68679, n68680, n68681, n68682, n68683, n68684,
         n68685, n68686, n68687, n68688, n68689, n68690, n68691, n68692,
         n68693, n68694, n68695, n68696, n68697, n68698, n68699, n68700,
         n68701, n68702, n68703, n68704, n68705, n68706, n68707, n68708,
         n68709, n68710, n68711, n68712, n68713, n68714, n68715, n68716,
         n68717, n68718, n68719, n68720, n68721, n68722, n68723, n68724,
         n68725, n68726, n68727, n68728, n68729, n68730, n68731, n68732,
         n68733, n68734, n68735, n68736, n68737, n68738, n68739, n68740,
         n68741, n68742, n68743, n68744, n68745, n68746, n68747, n68748,
         n68749, n68750, n68751, n68752, n68753, n68754, n68755, n68756,
         n68757, n68758, n68759, n68760, n68761, n68762, n68763, n68764,
         n68765, n68766, n68767, n68768, n68769, n68770, n68771, n68772,
         n68773, n68774, n68775, n68776, n68777, n68778, n68779, n68780,
         n68781, n68782, n68783, n68784, n68785, n68786, n68787, n68788,
         n68789, n68790, n68791, n68792, n68793, n68794, n68795, n68796,
         n68797, n68798, n68799, n68800, n68801, n68802, n68803, n68804,
         n68805, n68806, n68807, n68808, n68809, n68810, n68811, n68812,
         n68813, n68814, n68815, n68816, n68817, n68818, n68819, n68820,
         n68821, n68822, n68823, n68824, n68825, n68826, n68827, n68828,
         n68829, n68830, n68831, n68832, n68833, n68834, n68835, n68836,
         n68837, n68838, n68839, n68840, n68841, n68842, n68843, n68844,
         n68845, n68846, n68847, n68848, n68849, n68850, n68851, n68852,
         n68853, n68854, n68855, n68856, n68857, n68858, n68859, n68860,
         n68861, n68862, n68863, n68864, n68865, n68866, n68867, n68868,
         n68869, n68870, n68871, n68872, n68873, n68874, n68875, n68876,
         n68877, n68878, n68879, n68880, n68881, n68882, n68883, n68884,
         n68885, n68886, n68887, n68888, n68889, n68890, n68891, n68892,
         n68893, n68894, n68895, n68896, n68897, n68898, n68899, n68900,
         n68901, n68902, n68903, n68904, n68905, n68906, n68907, n68908,
         n68909, n68910, n68911, n68912, n68913, n68914, n68915, n68916,
         n68917, n68918, n68919, n68920, n68921, n68922, n68923, n68924,
         n68925, n68926, n68927, n68928, n68929, n68930, n68931, n68932,
         n68933, n68934, n68935, n68936, n68937, n68938, n68939, n68940,
         n68941, n68942, n68943, n68944, n68945, n68946, n68947, n68948,
         n68949, n68950, n68951, n68952, n68953, n68954, n68955, n68956,
         n68957, n68958, n68959, n68960, n68961, n68962, n68963, n68964,
         n68965, n68966, n68967, n68968, n68969, n68970, n68971, n68972,
         n68973, n68974, n68975, n68976, n68977, n68978, n68979, n68980,
         n68981, n68982, n68983, n68984, n68985, n68986, n68987, n68988,
         n68989, n68990, n68991, n68992, n68993, n68994, n68995, n68996,
         n68997, n68998, n68999, n69000, n69001, n69002, n69003, n69004,
         n69005, n69006, n69007, n69008, n69009, n69010, n69011, n69012,
         n69013, n69014, n69015, n69016, n69017, n69018, n69019, n69020,
         n69021, n69022, n69023, n69024, n69025, n69026, n69027, n69028,
         n69029, n69030, n69031, n69032, n69033, n69034, n69035, n69036,
         n69037, n69038, n69039, n69040, n69041, n69042, n69043, n69044,
         n69045, n69046, n69047, n69048, n69049, n69050, n69051, n69052,
         n69053, n69054, n69055, n69056, n69057, n69058, n69059, n69060,
         n69061, n69062, n69063, n69064, n69065, n69066, n69067, n69068,
         n69069, n69070, n69071, n69072, n69073, n69074, n69075, n69076,
         n69077, n69078, n69079, n69080, n69081, n69082, n69083, n69084,
         n69085, n69086, n69087, n69088, n69089, n69090, n69091, n69092,
         n69093, n69094, n69095, n69096, n69097, n69098, n69099, n69100,
         n69101, n69102, n69103, n69104, n69105, n69106, n69107, n69108,
         n69109, n69110, n69111, n69112, n69113, n69114, n69115, n69116,
         n69117, n69118, n69119, n69120, n69121, n69122, n69123, n69124,
         n69125, n69126, n69127, n69128, n69129, n69130, n69131, n69132,
         n69133, n69134, n69135, n69136, n69137, n69138, n69139, n69140,
         n69141, n69142, n69143, n69144, n69145, n69146, n69147, n69148,
         n69149, n69150, n69151, n69152, n69153, n69154, n69155, n69156,
         n69157, n69158, n69159, n69160, n69161, n69162, n69163, n69164,
         n69165, n69166, n69167, n69168, n69169, n69170, n69171, n69172,
         n69173, n69174, n69175, n69176, n69177, n69178, n69179, n69180,
         n69181, n69182, n69183, n69184, n69185, n69186, n69187, n69188,
         n69189, n69190, n69191, n69192, n69193, n69194, n69195, n69196,
         n69197, n69198, n69199, n69200, n69201, n69202, n69203, n69204,
         n69205, n69206, n69207, n69208, n69209, n69210, n69211, n69212,
         n69213, n69214, n69215, n69216, n69217, n69218, n69219, n69220,
         n69221, n69222, n69223, n69224, n69225, n69226, n69227, n69228,
         n69229, n69230, n69231, n69232, n69233, n69234, n69235, n69236,
         n69237, n69238, n69239, n69240, n69241, n69242, n69243, n69244,
         n69245, n69246, n69247, n69248, n69249, n69250, n69251, n69252,
         n69253, n69254, n69255, n69256, n69257, n69258, n69259, n69260,
         n69261, n69262, n69263, n69264, n69265, n69266, n69267, n69268,
         n69269, n69270, n69271, n69272, n69273, n69274, n69275, n69276,
         n69277, n69278, n69279, n69280, n69281, n69282, n69283, n69284,
         n69285, n69286, n69287, n69288, n69289, n69290, n69291, n69292,
         n69293, n69294, n69295, n69296, n69297, n69298, n69299, n69300,
         n69301, n69302, n69303, n69304, n69305, n69306, n69307, n69308,
         n69309, n69310, n69311, n69312, n69313, n69314, n69315, n69316,
         n69317, n69318, n69319, n69320, n69321, n69322, n69323, n69324,
         n69325, n69326, n69327, n69328, n69329, n69330, n69331, n69332,
         n69333, n69334, n69335, n69336, n69337, n69338, n69339, n69340,
         n69341, n69342, n69343, n69344, n69345, n69346, n69347, n69348,
         n69349, n69350, n69351, n69352, n69353, n69354, n69355, n69356,
         n69357, n69358, n69359, n69360, n69361, n69362, n69363, n69364,
         n69365, n69366, n69367, n69368, n69369, n69370, n69371, n69372,
         n69373, n69374, n69375, n69376, n69377, n69378, n69379, n69380,
         n69381, n69382, n69383, n69384, n69385, n69386, n69387, n69388,
         n69389, n69390, n69391, n69392, n69393, n69394, n69395, n69396,
         n69397, n69398, n69399, n69400, n69401, n69402, n69403, n69404,
         n69405, n69406, n69407, n69408, n69409, n69410, n69411, n69412,
         n69413, n69414, n69415, n69416, n69417, n69418, n69419, n69420,
         n69421, n69422, n69423, n69424, n69425, n69426, n69427, n69428,
         n69429, n69430, n69431, n69432, n69433, n69434, n69435, n69436,
         n69437, n69438, n69439, n69440, n69441, n69442, n69443, n69444,
         n69445, n69446, n69447, n69448, n69449, n69450, n69451, n69452,
         n69453, n69454, n69455, n69456, n69457, n69458, n69459, n69460,
         n69461, n69462, n69463, n69464, n69465, n69466, n69467, n69468,
         n69469, n69470, n69471, n69472, n69473, n69474, n69475, n69476,
         n69477, n69478, n69479, n69480, n69481, n69482, n69483, n69484,
         n69485, n69486, n69487, n69488, n69489, n69490, n69491, n69492,
         n69493, n69494, n69495, n69496, n69497, n69498, n69499, n69500,
         n69501, n69502, n69503, n69504, n69505, n69506, n69507, n69508,
         n69509, n69510, n69511, n69512, n69513, n69514, n69515, n69516,
         n69517, n69518, n69519, n69520, n69521, n69522, n69523, n69524,
         n69525, n69526, n69527, n69528, n69529, n69530, n69531, n69532,
         n69533, n69534, n69535, n69536, n69537, n69538, n69539, n69540,
         n69541, n69542, n69543, n69544, n69545, n69546, n69547, n69548,
         n69549, n69550, n69551, n69552, n69553, n69554, n69555, n69556,
         n69557, n69558, n69559, n69560, n69561, n69562, n69563, n69564,
         n69565, n69566, n69567, n69568, n69569, n69570, n69571, n69572,
         n69573, n69574, n69575, n69576, n69577, n69578, n69579, n69580,
         n69581, n69582, n69583, n69584, n69585, n69586, n69587, n69588,
         n69589, n69590, n69591, n69592, n69593, n69594, n69595, n69596,
         n69597, n69598, n69599, n69600, n69601, n69602, n69603, n69604,
         n69605, n69606, n69607, n69608, n69609, n69610, n69611, n69612,
         n69613, n69614, n69615, n69616, n69617, n69618, n69619, n69620,
         n69621, n69622, n69623, n69624, n69625, n69626, n69627, n69628,
         n69629, n69630, n69631, n69632, n69633, n69634, n69635, n69636,
         n69637, n69638, n69639, n69640, n69641, n69642, n69643, n69644,
         n69645, n69646, n69647, n69648, n69649, n69650, n69651, n69652,
         n69653, n69654, n69655, n69656, n69657, n69658, n69659, n69660,
         n69661, n69662, n69663, n69664, n69665, n69666, n69667, n69668,
         n69669, n69670, n69671, n69672, n69673, n69674, n69675, n69676,
         n69677, n69678, n69679, n69680, n69681, n69682, n69683, n69684,
         n69685, n69686, n69687, n69688, n69689, n69690, n69691, n69692,
         n69693, n69694, n69695, n69696, n69697, n69698, n69699, n69700,
         n69701, n69702, n69703, n69704, n69705, n69706, n69707, n69708,
         n69709, n69710, n69711, n69712, n69713, n69714, n69715, n69716,
         n69717, n69718, n69719, n69720, n69721, n69722, n69723, n69724,
         n69725, n69726, n69727, n69728, n69729, n69730, n69731, n69732,
         n69733, n69734, n69735, n69736, n69737, n69738, n69739, n69740,
         n69741, n69742, n69743, n69744, n69745, n69746, n69747, n69748,
         n69749, n69750, n69751, n69752, n69753, n69754, n69755, n69756,
         n69757, n69758, n69759, n69760, n69761, n69762, n69763, n69764,
         n69765, n69766, n69767, n69768, n69769, n69770, n69771, n69772,
         n69773, n69774, n69775, n69776, n69777, n69778, n69779, n69780,
         n69781, n69782, n69783, n69784, n69785, n69786, n69787, n69788,
         n69789, n69790, n69791, n69792, n69793, n69794, n69795, n69796,
         n69797, n69798, n69799, n69800, n69801, n69802, n69803, n69804,
         n69805, n69806, n69807, n69808, n69809, n69810, n69811, n69812,
         n69813, n69814, n69815, n69816, n69817, n69818, n69819, n69820,
         n69821, n69822, n69823, n69824, n69825, n69826, n69827, n69828,
         n69829, n69830, n69831, n69832, n69833, n69834, n69835, n69836,
         n69837, n69838, n69839, n69840, n69841, n69842, n69843, n69844,
         n69845, n69846, n69847, n69848, n69849, n69850, n69851, n69852,
         n69853, n69854, n69855, n69856, n69857, n69858, n69859, n69860,
         n69861, n69862, n69863, n69864, n69865, n69866, n69867, n69868,
         n69869, n69870, n69871, n69872, n69873, n69874, n69875, n69876,
         n69877, n69878, n69879, n69880, n69881, n69882, n69883, n69884,
         n69885, n69886, n69887, n69888, n69889, n69890, n69891, n69892,
         n69893, n69894, n69895, n69896, n69897, n69898, n69899, n69900,
         n69901, n69902, n69903, n69904, n69905, n69906, n69907, n69908,
         n69909, n69910, n69911, n69912, n69913, n69914, n69915, n69916,
         n69917, n69918, n69919, n69920, n69921, n69922, n69923, n69924,
         n69925, n69926, n69927, n69928, n69929, n69930, n69931, n69932,
         n69933, n69934, n69935, n69936, n69937, n69938, n69939, n69940,
         n69941, n69942, n69943, n69944, n69945, n69946, n69947, n69948,
         n69949, n69950, n69951, n69952, n69953, n69954, n69955, n69956,
         n69957, n69958, n69959, n69960, n69961, n69962, n69963, n69964,
         n69965, n69966, n69967, n69968, n69969, n69970, n69971, n69972,
         n69973, n69974, n69975, n69976, n69977, n69978, n69979, n69980,
         n69981, n69982, n69983, n69984, n69985, n69986, n69987, n69988,
         n69989, n69990, n69991, n69992, n69993, n69994, n69995, n69996,
         n69997, n69998, n69999, n70000, n70001, n70002, n70003, n70004,
         n70005, n70006, n70007, n70008, n70009, n70010, n70011, n70012,
         n70013, n70014, n70015, n70016, n70017, n70018, n70019, n70020,
         n70021, n70022, n70023, n70024, n70025, n70026, n70027, n70028,
         n70029, n70030, n70031, n70032, n70033, n70034, n70035, n70036,
         n70037, n70038, n70039, n70040, n70041, n70042, n70043, n70044,
         n70045, n70046, n70047, n70048, n70049, n70050, n70051, n70052,
         n70053, n70054, n70055, n70056, n70057, n70058, n70059, n70060,
         n70061, n70062, n70063, n70064, n70065, n70066, n70067, n70068,
         n70069, n70070, n70071, n70072, n70073, n70074, n70075, n70076,
         n70077, n70078, n70079, n70080, n70081, n70082, n70083, n70084,
         n70085, n70086, n70087, n70088, n70089, n70090, n70091, n70092,
         n70093, n70094, n70095, n70096, n70097, n70098, n70099, n70100,
         n70101, n70102, n70103, n70104, n70105, n70106, n70107, n70108,
         n70109, n70110, n70111, n70112, n70113, n70114, n70115, n70116,
         n70117, n70118, n70119, n70120, n70121, n70122, n70123, n70124,
         n70125, n70126, n70127, n70128, n70129, n70130, n70131, n70132,
         n70133, n70134, n70135, n70136, n70137, n70138, n70139, n70140,
         n70141, n70142, n70143, n70144, n70145, n70146, n70147, n70148,
         n70149, n70150, n70151, n70152, n70153, n70154, n70155, n70156,
         n70157, n70158, n70159, n70160, n70161, n70162, n70163, n70164,
         n70165, n70166, n70167, n70168, n70169, n70170, n70171, n70172,
         n70173, n70174, n70175, n70176, n70177, n70178, n70179, n70180,
         n70181, n70182, n70183, n70184, n70185, n70186, n70187, n70188,
         n70189, n70190, n70191, n70192, n70193, n70194, n70195, n70196,
         n70197, n70198, n70199, n70200, n70201, n70202, n70203, n70204,
         n70205, n70206, n70207, n70208, n70209, n70210, n70211, n70212,
         n70213, n70214, n70215, n70216, n70217, n70218, n70219, n70220,
         n70221, n70222, n70223, n70224, n70225, n70226, n70227, n70228,
         n70229, n70230, n70231, n70232, n70233, n70234, n70235, n70236,
         n70237, n70238, n70239, n70240, n70241, n70242, n70243, n70244,
         n70245, n70246, n70247, n70248, n70249, n70250, n70251, n70252,
         n70253, n70254, n70255, n70256, n70257, n70258, n70259, n70260,
         n70261, n70262, n70263, n70264, n70265, n70266, n70267, n70268,
         n70269, n70270, n70271, n70272, n70273, n70274, n70275, n70276,
         n70277, n70278, n70279, n70280, n70281, n70282, n70283, n70284,
         n70285, n70286, n70287, n70288, n70289, n70290, n70291, n70292,
         n70293, n70294, n70295, n70296, n70297, n70298, n70299, n70300,
         n70301, n70302, n70303, n70304, n70305, n70306, n70307, n70308,
         n70309, n70310, n70311, n70312, n70313, n70314, n70315, n70316,
         n70317, n70318, n70319, n70320, n70321, n70322, n70323, n70324,
         n70325, n70326, n70327, n70328, n70329, n70330, n70331, n70332,
         n70333, n70334, n70335, n70336, n70337, n70338, n70339, n70340,
         n70341, n70342, n70343, n70344, n70345, n70346, n70347, n70348,
         n70349, n70350, n70351, n70352, n70353, n70354, n70355, n70356,
         n70357, n70358, n70359, n70360, n70361, n70362, n70363, n70364,
         n70365, n70366, n70367, n70368, n70369, n70370, n70371, n70372,
         n70373, n70374, n70375, n70376, n70377, n70378, n70379, n70380,
         n70381, n70382, n70383, n70384, n70385, n70386, n70387, n70388,
         n70389, n70390, n70391, n70392, n70393, n70394, n70395, n70396,
         n70397, n70398, n70399, n70400, n70401, n70402, n70403, n70404,
         n70405, n70406, n70407, n70408, n70409, n70410, n70411, n70412,
         n70413, n70414, n70415, n70416, n70417, n70418, n70419, n70420,
         n70421, n70422, n70423, n70424, n70425, n70426, n70427, n70428,
         n70429, n70430, n70431, n70432, n70433, n70434, n70435, n70436,
         n70437, n70438, n70439, n70440, n70441, n70442, n70443, n70444,
         n70445, n70446, n70447, n70448, n70449, n70450, n70451, n70452,
         n70453, n70454, n70455, n70456, n70457, n70458, n70459, n70460,
         n70461, n70462, n70463, n70464, n70465, n70466, n70467, n70468,
         n70469, n70470, n70471, n70472, n70473, n70474, n70475, n70476,
         n70477, n70478, n70479, n70480, n70481, n70482, n70483, n70484,
         n70485, n70486, n70487, n70488, n70489, n70490, n70491, n70492,
         n70493, n70494, n70495, n70496, n70497, n70498, n70499, n70500,
         n70501, n70502, n70503, n70504, n70505, n70506, n70507, n70508,
         n70509, n70510, n70511, n70512, n70513, n70514, n70515, n70516,
         n70517, n70518, n70519, n70520, n70521, n70522, n70523, n70524,
         n70525, n70526, n70527, n70528, n70529, n70530, n70531, n70532,
         n70533, n70534, n70535, n70536, n70537, n70538, n70539, n70540,
         n70541, n70542, n70543, n70544, n70545, n70546, n70547, n70548,
         n70549, n70550, n70551, n70552, n70553, n70554, n70555, n70556,
         n70557, n70558, n70559, n70560, n70561, n70562, n70563, n70564,
         n70565, n70566, n70567, n70568, n70569, n70570, n70571, n70572,
         n70573, n70574, n70575, n70576, n70577, n70578, n70579, n70580,
         n70581, n70582, n70583, n70584, n70585, n70586, n70587, n70588,
         n70589, n70590, n70591, n70592, n70593, n70594, n70595, n70596,
         n70597, n70598, n70599, n70600, n70601, n70602, n70603, n70604,
         n70605, n70606, n70607, n70608, n70609, n70610, n70611, n70612,
         n70613, n70614, n70615, n70616, n70617, n70618, n70619, n70620,
         n70621, n70622, n70623, n70624, n70625, n70626, n70627, n70628,
         n70629, n70630, n70631, n70632, n70633, n70634, n70635, n70636,
         n70637, n70638, n70639, n70640, n70641, n70642, n70643, n70644,
         n70645, n70646, n70647, n70648, n70649, n70650, n70651, n70652,
         n70653, n70654, n70655, n70656, n70657, n70658, n70659, n70660,
         n70661, n70662, n70663, n70664, n70665, n70666, n70667, n70668,
         n70669, n70670, n70671, n70672, n70673, n70674, n70675, n70676,
         n70677, n70678, n70679, n70680, n70681, n70682, n70683, n70684,
         n70685, n70686, n70687, n70688, n70689, n70690, n70691, n70692,
         n70693, n70694, n70695, n70696, n70697, n70698, n70699, n70700,
         n70701, n70702, n70703, n70704, n70705, n70706, n70707, n70708,
         n70709, n70710, n70711, n70712, n70713, n70714, n70715, n70716,
         n70717, n70718, n70719, n70720, n70721, n70722, n70723, n70724,
         n70725, n70726, n70727, n70728, n70729, n70730, n70731, n70732,
         n70733, n70734, n70735, n70736, n70737, n70738, n70739, n70740,
         n70741, n70742, n70743, n70744, n70745, n70746, n70747, n70748,
         n70749, n70750, n70751, n70752, n70753, n70754, n70755, n70756,
         n70757, n70758, n70759, n70760, n70761, n70762, n70763, n70764,
         n70765, n70766, n70767, n70768, n70769, n70770, n70771, n70772,
         n70773, n70774, n70775, n70776, n70777, n70778, n70779, n70780,
         n70781, n70782, n70783, n70784, n70785, n70786, n70787, n70788,
         n70789, n70790, n70791, n70792, n70793, n70794, n70795, n70796,
         n70797, n70798, n70799, n70800, n70801, n70802, n70803, n70804,
         n70805, n70806, n70807, n70808, n70809, n70810, n70811, n70812,
         n70813, n70814, n70815, n70816, n70817, n70818, n70819, n70820,
         n70821, n70822, n70823, n70824, n70825, n70826, n70827, n70828,
         n70829, n70830, n70831, n70832, n70833, n70834, n70835, n70836,
         n70837, n70838, n70839, n70840, n70841, n70842, n70843, n70844,
         n70845, n70846, n70847, n70848, n70849, n70850, n70851, n70852,
         n70853, n70854, n70855, n70856, n70857, n70858, n70859, n70860,
         n70861, n70862, n70863, n70864, n70865, n70866, n70867, n70868,
         n70869, n70870, n70871, n70872, n70873, n70874, n70875, n70876,
         n70877, n70878, n70879, n70880, n70881, n70882, n70883, n70884,
         n70885, n70886, n70887, n70888, n70889, n70890, n70891, n70892,
         n70893, n70894, n70895, n70896, n70897, n70898, n70899, n70900,
         n70901, n70902, n70903, n70904, n70905, n70906, n70907, n70908,
         n70909, n70910, n70911, n70912, n70913, n70914, n70915, n70916,
         n70917, n70918, n70919, n70920, n70921, n70922, n70923, n70924,
         n70925, n70926, n70927, n70928, n70929, n70930, n70931, n70932,
         n70933, n70934, n70935, n70936, n70937, n70938, n70939, n70940,
         n70941, n70942, n70943, n70944, n70945, n70946, n70947, n70948,
         n70949, n70950, n70951, n70952, n70953, n70954, n70955, n70956,
         n70957, n70958, n70959, n70960, n70961, n70962, n70963, n70964,
         n70965, n70966, n70967, n70968, n70969, n70970, n70971, n70972,
         n70973, n70974, n70975, n70976, n70977, n70978, n70979, n70980,
         n70981, n70982, n70983, n70984, n70985, n70986, n70987, n70988,
         n70989, n70990, n70991, n70992, n70993, n70994, n70995, n70996,
         n70997, n70998, n70999, n71000, n71001, n71002, n71003, n71004,
         n71005, n71006, n71007, n71008, n71009, n71010, n71011, n71012,
         n71013, n71014, n71015, n71016, n71017, n71018, n71019, n71020,
         n71021, n71022, n71023, n71024, n71025, n71026, n71027, n71028,
         n71029, n71030, n71031, n71032, n71033, n71034, n71035, n71036,
         n71037, n71038, n71039, n71040, n71041, n71042, n71043, n71044,
         n71045, n71046, n71047, n71048, n71049, n71050, n71051, n71052,
         n71053, n71054, n71055, n71056, n71057, n71058, n71059, n71060,
         n71061, n71062, n71063, n71064, n71065, n71066, n71067, n71068,
         n71069, n71070, n71071, n71072, n71073, n71074, n71075, n71076,
         n71077, n71078, n71079, n71080, n71081, n71082, n71083, n71084,
         n71085, n71086, n71087, n71088, n71089, n71090, n71091, n71092,
         n71093, n71094, n71095, n71096, n71097, n71098, n71099, n71100,
         n71101, n71102, n71103, n71104, n71105, n71106, n71107, n71108,
         n71109, n71110, n71111, n71112, n71113, n71114, n71115, n71116,
         n71117, n71118, n71119, n71120, n71121, n71122, n71123, n71124,
         n71125, n71126, n71127, n71128, n71129, n71130, n71131, n71132,
         n71133, n71134, n71135, n71136, n71137, n71138, n71139, n71140,
         n71141, n71142, n71143, n71144, n71145, n71146, n71147, n71148,
         n71149, n71150, n71151, n71152, n71153, n71154, n71155, n71156,
         n71157, n71158, n71159, n71160, n71161, n71162, n71163, n71164,
         n71165, n71166, n71167, n71168, n71169, n71170, n71171, n71172,
         n71173, n71174, n71175, n71176, n71177, n71178, n71179, n71180,
         n71181, n71182, n71183, n71184, n71185, n71186, n71187, n71188,
         n71189, n71190, n71191, n71192, n71193, n71194, n71195, n71196,
         n71197, n71198, n71199, n71200, n71201, n71202, n71203, n71204,
         n71205, n71206, n71207, n71208, n71209, n71210, n71211, n71212,
         n71213, n71214, n71215, n71216, n71217, n71218, n71219, n71220,
         n71221, n71222, n71223, n71224, n71225, n71226, n71227, n71228,
         n71229, n71230, n71231, n71232, n71233, n71234, n71235, n71236,
         n71237, n71238, n71239, n71240, n71241, n71242, n71243, n71244,
         n71245, n71246, n71247, n71248, n71249, n71250, n71251, n71252,
         n71253, n71254, n71255, n71256, n71257, n71258, n71259, n71260,
         n71261, n71262, n71263, n71264, n71265, n71266, n71267, n71268,
         n71269, n71270, n71271, n71272, n71273, n71274, n71275, n71276,
         n71277, n71278, n71279, n71280, n71281, n71282, n71283, n71284,
         n71285, n71286, n71287, n71288, n71289, n71290, n71291, n71292,
         n71293, n71294, n71295, n71296, n71297, n71298, n71299, n71300,
         n71301, n71302, n71303, n71304, n71305, n71306, n71307, n71308,
         n71309, n71310, n71311, n71312, n71313, n71314, n71315, n71316,
         n71317, n71318, n71319, n71320, n71321, n71322, n71323, n71324,
         n71325, n71326, n71327, n71328, n71329, n71330, n71331, n71332,
         n71333, n71334, n71335, n71336, n71337, n71338, n71339, n71340,
         n71341, n71342, n71343, n71344, n71345, n71346, n71347, n71348,
         n71349, n71350, n71351, n71352, n71353, n71354, n71355, n71356,
         n71357, n71358, n71359, n71360, n71361, n71362, n71363, n71364,
         n71365, n71366, n71367, n71368, n71369, n71370, n71371, n71372,
         n71373, n71374, n71375, n71376, n71377, n71378, n71379, n71380,
         n71381, n71382, n71383, n71384, n71385, n71386, n71387, n71388,
         n71389, n71390, n71391, n71392, n71393, n71394, n71395, n71396,
         n71397, n71398, n71399, n71400, n71401, n71402, n71403, n71404,
         n71405, n71406, n71407, n71408, n71409, n71410, n71411, n71412,
         n71413, n71414, n71415, n71416, n71417, n71418, n71419, n71420,
         n71421, n71422, n71423, n71424, n71425, n71426, n71427, n71428,
         n71429, n71430, n71431, n71432, n71433, n71434, n71435, n71436,
         n71437, n71438, n71439, n71440, n71441, n71442, n71443, n71444,
         n71445, n71446, n71447, n71448, n71449, n71450, n71451, n71452,
         n71453, n71454, n71455, n71456, n71457, n71458, n71459, n71460,
         n71461, n71462, n71463, n71464, n71465, n71466, n71467, n71468,
         n71469, n71470, n71471, n71472, n71473, n71474, n71475, n71476,
         n71477, n71478, n71479, n71480, n71481, n71482, n71483, n71484,
         n71485, n71486, n71487, n71488, n71489, n71490, n71491, n71492,
         n71493, n71494, n71495, n71496, n71497, n71498, n71499, n71500,
         n71501, n71502, n71503, n71504, n71505, n71506, n71507, n71508,
         n71509, n71510, n71511, n71512, n71513, n71514, n71515, n71516,
         n71517, n71518, n71519, n71520, n71521, n71522, n71523, n71524,
         n71525, n71526, n71527, n71528, n71529, n71530, n71531, n71532,
         n71533, n71534, n71535, n71536, n71537, n71538, n71539, n71540,
         n71541, n71542, n71543, n71544, n71545, n71546, n71547, n71548,
         n71549, n71550, n71551, n71552, n71553, n71554, n71555, n71556,
         n71557, n71558, n71559, n71560, n71561, n71562, n71563, n71564,
         n71565, n71566, n71567, n71568, n71569, n71570, n71571, n71572,
         n71573, n71574, n71575, n71576, n71577, n71578, n71579, n71580,
         n71581, n71582, n71583, n71584, n71585, n71586, n71587, n71588,
         n71589, n71590, n71591, n71592, n71593, n71594, n71595, n71596,
         n71597, n71598, n71599, n71600, n71601, n71602, n71603, n71604,
         n71605, n71606, n71607, n71608, n71609, n71610, n71611, n71612,
         n71613, n71614, n71615, n71616, n71617, n71618, n71619, n71620,
         n71621, n71622, n71623, n71624, n71625, n71626, n71627, n71628,
         n71629, n71630, n71631, n71632, n71633, n71634, n71635, n71636,
         n71637, n71638, n71639, n71640, n71641, n71642, n71643, n71644,
         n71645, n71646, n71647, n71648, n71649, n71650, n71651, n71652,
         n71653, n71654, n71655, n71656, n71657, n71658, n71659, n71660,
         n71661, n71662, n71663, n71664, n71665, n71666, n71667, n71668,
         n71669, n71670, n71671, n71672, n71673, n71674, n71675, n71676,
         n71677, n71678, n71679, n71680, n71681, n71682, n71683, n71684,
         n71685, n71686, n71687, n71688, n71689, n71690, n71691, n71692,
         n71693, n71694, n71695, n71696, n71697, n71698, n71699, n71700,
         n71701, n71702, n71703, n71704, n71705, n71706, n71707, n71708,
         n71709, n71710, n71711, n71712, n71713, n71714, n71715, n71716,
         n71717, n71718, n71719, n71720, n71721, n71722, n71723, n71724,
         n71725, n71726, n71727, n71728, n71729, n71730, n71731, n71732,
         n71733, n71734, n71735, n71736, n71737, n71738, n71739, n71740,
         n71741, n71742, n71743, n71744, n71745, n71746, n71747, n71748,
         n71749, n71750, n71751, n71752, n71753, n71754, n71755, n71756,
         n71757, n71758, n71759, n71760, n71761, n71762, n71763, n71764,
         n71765, n71766, n71767, n71768, n71769, n71770, n71771, n71772,
         n71773, n71774, n71775, n71776, n71777, n71778, n71779, n71780,
         n71781, n71782, n71783, n71784, n71785, n71786, n71787, n71788,
         n71789, n71790, n71791, n71792, n71793, n71794, n71795, n71796,
         n71797, n71798, n71799, n71800, n71801, n71802, n71803, n71804,
         n71805, n71806, n71807, n71808, n71809, n71810, n71811, n71812,
         n71813, n71814, n71815, n71816, n71817, n71818, n71819, n71820,
         n71821, n71822, n71823, n71824, n71825, n71826, n71827, n71828,
         n71829, n71830, n71831, n71832, n71833, n71834, n71835, n71836,
         n71837, n71838, n71839, n71840, n71841, n71842, n71843, n71844,
         n71845, n71846, n71847, n71848, n71849, n71850, n71851, n71852,
         n71853, n71854, n71855, n71856, n71857, n71858, n71859, n71860,
         n71861, n71862, n71863, n71864, n71865, n71866, n71867, n71868,
         n71869, n71870, n71871, n71872, n71873, n71874, n71875, n71876,
         n71877, n71878, n71879, n71880, n71881, n71882, n71883, n71884,
         n71885, n71886, n71887, n71888, n71889, n71890, n71891, n71892,
         n71893, n71894, n71895, n71896, n71897, n71898, n71899, n71900,
         n71901, n71902, n71903, n71904, n71905, n71906, n71907, n71908,
         n71909, n71910, n71911, n71912, n71913, n71914, n71915, n71916,
         n71917, n71918, n71919, n71920, n71921, n71922, n71923, n71924,
         n71925, n71926, n71927, n71928, n71929, n71930, n71931, n71932,
         n71933, n71934, n71935, n71936, n71937, n71938, n71939, n71940,
         n71941, n71942, n71943, n71944, n71945, n71946, n71947, n71948,
         n71949, n71950, n71951, n71952, n71953, n71954, n71955, n71956,
         n71957, n71958, n71959, n71960, n71961, n71962, n71963, n71964,
         n71965, n71966, n71967, n71968, n71969, n71970, n71971, n71972,
         n71973, n71974, n71975, n71976, n71977, n71978, n71979, n71980,
         n71981, n71982, n71983, n71984, n71985, n71986, n71987, n71988,
         n71989, n71990, n71991, n71992, n71993, n71994, n71995, n71996,
         n71997, n71998, n71999, n72000, n72001, n72002, n72003, n72004,
         n72005, n72006, n72007, n72008, n72009, n72010, n72011, n72012,
         n72013, n72014, n72015, n72016, n72017, n72018, n72019, n72020,
         n72021, n72022, n72023, n72024, n72025, n72026, n72027, n72028,
         n72029, n72030, n72031, n72032, n72033, n72034, n72035, n72036,
         n72037, n72038, n72039, n72040, n72041, n72042, n72043, n72044,
         n72045, n72046, n72047, n72048, n72049, n72050, n72051, n72052,
         n72053, n72054, n72055, n72056, n72057, n72058, n72059, n72060,
         n72061, n72062, n72063, n72064, n72065, n72066, n72067, n72068,
         n72069, n72070, n72071, n72072, n72073, n72074, n72075, n72076,
         n72077, n72078, n72079, n72080, n72081, n72082, n72083, n72084,
         n72085, n72086, n72087, n72088, n72089, n72090, n72091, n72092,
         n72093, n72094, n72095, n72096, n72097, n72098, n72099, n72100,
         n72101, n72102, n72103, n72104, n72105, n72106, n72107, n72108,
         n72109, n72110, n72111, n72112, n72113, n72114, n72115, n72116,
         n72117, n72118, n72119, n72120, n72121, n72122, n72123, n72124,
         n72125, n72126, n72127, n72128, n72129, n72130, n72131, n72132,
         n72133, n72134, n72135, n72136, n72137, n72138, n72139, n72140,
         n72141, n72142, n72143, n72144, n72145, n72146, n72147, n72148,
         n72149, n72150, n72151, n72152, n72153, n72154, n72155, n72156,
         n72157, n72158, n72159, n72160, n72161, n72162, n72163, n72164,
         n72165, n72166, n72167, n72168, n72169, n72170, n72171, n72172,
         n72173, n72174, n72175, n72176, n72177, n72178, n72179, n72180,
         n72181, n72182, n72183, n72184, n72185, n72186, n72187, n72188,
         n72189, n72190, n72191, n72192, n72193, n72194, n72195, n72196,
         n72197, n72198, n72199, n72200, n72201, n72202, n72203, n72204,
         n72205, n72206, n72207, n72208, n72209, n72210, n72211, n72212,
         n72213, n72214, n72215, n72216, n72217, n72218, n72219, n72220,
         n72221, n72222, n72223, n72224, n72225, n72226, n72227, n72228,
         n72229, n72230, n72231, n72232, n72233, n72234, n72235, n72236,
         n72237, n72238, n72239, n72240, n72241, n72242, n72243, n72244,
         n72245, n72246, n72247, n72248, n72249, n72250, n72251, n72252,
         n72253, n72254, n72255, n72256, n72257, n72258, n72259, n72260,
         n72261, n72262, n72263, n72264, n72265, n72266, n72267, n72268,
         n72269, n72270, n72271, n72272, n72273, n72274, n72275, n72276,
         n72277, n72278, n72279, n72280, n72281, n72282, n72283, n72284,
         n72285, n72286, n72287, n72288, n72289, n72290, n72291, n72292,
         n72293, n72294, n72295, n72296, n72297, n72298, n72299, n72300,
         n72301, n72302, n72303, n72304, n72305, n72306, n72307, n72308,
         n72309, n72310, n72311, n72312, n72313, n72314, n72315, n72316,
         n72317, n72318, n72319, n72320, n72321, n72322, n72323, n72324,
         n72325, n72326, n72327, n72328, n72329, n72330, n72331, n72332,
         n72333, n72334, n72335, n72336, n72337, n72338, n72339, n72340,
         n72341, n72342, n72343, n72344, n72345, n72346, n72347, n72348,
         n72349, n72350, n72351, n72352, n72353, n72354, n72355, n72356,
         n72357, n72358, n72359, n72360, n72361, n72362, n72363, n72364,
         n72365, n72366, n72367, n72368, n72369, n72370, n72371, n72372,
         n72373, n72374, n72375, n72376, n72377, n72378, n72379, n72380,
         n72381, n72382, n72383, n72384, n72385, n72386, n72387, n72388,
         n72389, n72390, n72391, n72392, n72393, n72394, n72395, n72396,
         n72397, n72398, n72399, n72400, n72401, n72402, n72403, n72404,
         n72405, n72406, n72407, n72408, n72409, n72410, n72411, n72412,
         n72413, n72414, n72415, n72416, n72417, n72418, n72419, n72420,
         n72421, n72422, n72423, n72424, n72425, n72426, n72427, n72428,
         n72429, n72430, n72431, n72432, n72433, n72434, n72435, n72436,
         n72437, n72438, n72439, n72440, n72441, n72442, n72443, n72444,
         n72445, n72446, n72447, n72448, n72449, n72450, n72451, n72452,
         n72453, n72454, n72455, n72456, n72457, n72458, n72459, n72460,
         n72461, n72462, n72463, n72464, n72465, n72466, n72467, n72468,
         n72469, n72470, n72471, n72472, n72473, n72474, n72475, n72476,
         n72477, n72478, n72479, n72480, n72481, n72482, n72483, n72484,
         n72485, n72486, n72487, n72488, n72489, n72490, n72491, n72492,
         n72493, n72494, n72495, n72496, n72497, n72498, n72499, n72500,
         n72501, n72502, n72503, n72504, n72505, n72506, n72507, n72508,
         n72509, n72510, n72511, n72512, n72513, n72514, n72515, n72516,
         n72517, n72518, n72519, n72520, n72521, n72522, n72523, n72524,
         n72525, n72526, n72527, n72528, n72529, n72530, n72531, n72532,
         n72533, n72534, n72535, n72536, n72537, n72538, n72539, n72540,
         n72541, n72542, n72543, n72544, n72545, n72546, n72547, n72548,
         n72549, n72550, n72551, n72552, n72553, n72554, n72555, n72556,
         n72557, n72558, n72559, n72560, n72561, n72562, n72563, n72564,
         n72565, n72566, n72567, n72568, n72569, n72570, n72571, n72572,
         n72573, n72574, n72575, n72576, n72577, n72578, n72579, n72580,
         n72581, n72582, n72583, n72584, n72585, n72586, n72587, n72588,
         n72589, n72590, n72591, n72592, n72593, n72594, n72595, n72596,
         n72597, n72598, n72599, n72600, n72601, n72602, n72603, n72604,
         n72605, n72606, n72607, n72608, n72609, n72610, n72611, n72612,
         n72613, n72614, n72615, n72616, n72617, n72618, n72619, n72620,
         n72621, n72622, n72623, n72624, n72625, n72626, n72627, n72628,
         n72629, n72630, n72631, n72632, n72633, n72634, n72635, n72636,
         n72637, n72638, n72639, n72640, n72641, n72642, n72643, n72644,
         n72645, n72646, n72647, n72648, n72649, n72650, n72651, n72652,
         n72653, n72654, n72655, n72656, n72657, n72658, n72659, n72660,
         n72661, n72662, n72663, n72664, n72665, n72666, n72667, n72668,
         n72669, n72670, n72671, n72672, n72673, n72674, n72675, n72676,
         n72677, n72678, n72679, n72680, n72681, n72682, n72683, n72684,
         n72685, n72686, n72687, n72688, n72689, n72690, n72691, n72692,
         n72693, n72694, n72695, n72696, n72697, n72698, n72699, n72700,
         n72701, n72702, n72703, n72704, n72705, n72706, n72707, n72708,
         n72709, n72710, n72711, n72712, n72713, n72714, n72715, n72716,
         n72717, n72718, n72719, n72720, n72721, n72722, n72723, n72724,
         n72725, n72726, n72727, n72728, n72729, n72730, n72731, n72732,
         n72733, n72734, n72735, n72736, n72737, n72738, n72739, n72740,
         n72741, n72742, n72743, n72744, n72745, n72746, n72747, n72748,
         n72749, n72750, n72751, n72752, n72753, n72754, n72755, n72756,
         n72757, n72758, n72759, n72760, n72761, n72762, n72763, n72764,
         n72765, n72766, n72767, n72768, n72769, n72770, n72771, n72772,
         n72773, n72774, n72775, n72776, n72777, n72778, n72779, n72780,
         n72781, n72782, n72783, n72784, n72785, n72786, n72787, n72788,
         n72789, n72790, n72791, n72792, n72793, n72794, n72795, n72796,
         n72797, n72798, n72799, n72800, n72801, n72802, n72803, n72804,
         n72805, n72806, n72807, n72808, n72809, n72810, n72811, n72812,
         n72813, n72814, n72815, n72816, n72817, n72818, n72819, n72820,
         n72821, n72822, n72823, n72824, n72825, n72826, n72827, n72828,
         n72829, n72830, n72831, n72832, n72833, n72834, n72835, n72836,
         n72837, n72838, n72839, n72840, n72841, n72842, n72843, n72844,
         n72845, n72846, n72847, n72848, n72849, n72850, n72851, n72852,
         n72853, n72854, n72855, n72856, n72857, n72858, n72859, n72860,
         n72861, n72862, n72863, n72864, n72865, n72866, n72867, n72868,
         n72869, n72870, n72871, n72872, n72873, n72874, n72875, n72876,
         n72877, n72878, n72879, n72880, n72881, n72882, n72883, n72884,
         n72885, n72886, n72887, n72888, n72889, n72890, n72891, n72892,
         n72893, n72894, n72895, n72896, n72897, n72898, n72899, n72900,
         n72901, n72902, n72903, n72904, n72905, n72906, n72907, n72908,
         n72909, n72910, n72911, n72912, n72913, n72914, n72915, n72916,
         n72917, n72918, n72919, n72920, n72921, n72922, n72923, n72924,
         n72925, n72926, n72927, n72928, n72929, n72930, n72931, n72932,
         n72933, n72934, n72935, n72936, n72937, n72938, n72939, n72940,
         n72941, n72942, n72943, n72944, n72945, n72946, n72947, n72948,
         n72949, n72950, n72951, n72952, n72953, n72954, n72955, n72956,
         n72957, n72958, n72959, n72960, n72961, n72962, n72963, n72964,
         n72965, n72966, n72967, n72968, n72969, n72970, n72971, n72972,
         n72973, n72974, n72975, n72976, n72977, n72978, n72979, n72980,
         n72981, n72982, n72983, n72984, n72985, n72986, n72987, n72988,
         n72989, n72990, n72991, n72992, n72993, n72994, n72995, n72996,
         n72997, n72998, n72999, n73000, n73001, n73002, n73003, n73004,
         n73005, n73006, n73007, n73008, n73009, n73010, n73011, n73012,
         n73013, n73014, n73015, n73016, n73017, n73018, n73019, n73020,
         n73021, n73022, n73023, n73024, n73025, n73026, n73027, n73028,
         n73029, n73030, n73031, n73032, n73033, n73034, n73035, n73036,
         n73037, n73038, n73039, n73040, n73041, n73042, n73043, n73044,
         n73045, n73046, n73047, n73048, n73049, n73050, n73051, n73052,
         n73053, n73054, n73055, n73056, n73057, n73058, n73059, n73060,
         n73061, n73062, n73063, n73064, n73065, n73066, n73067, n73068,
         n73069, n73070, n73071, n73072, n73073, n73074, n73075, n73076,
         n73077, n73078, n73079, n73080, n73081, n73082, n73083, n73084,
         n73085, n73086, n73087, n73088, n73089, n73090, n73091, n73092,
         n73093, n73094, n73095, n73096, n73097, n73098, n73099, n73100,
         n73101, n73102, n73103, n73104, n73105, n73106, n73107, n73108,
         n73109, n73110, n73111, n73112, n73113, n73114, n73115, n73116,
         n73117, n73118, n73119, n73120, n73121, n73122, n73123, n73124,
         n73125, n73126, n73127, n73128, n73129, n73130, n73131, n73132,
         n73133, n73134, n73135, n73136, n73137, n73138, n73139, n73140,
         n73141, n73142, n73143, n73144, n73145, n73146, n73147, n73148,
         n73149, n73150, n73151, n73152, n73153, n73154, n73155, n73156,
         n73157, n73158, n73159, n73160, n73161, n73162, n73163, n73164,
         n73165, n73166, n73167, n73168, n73169, n73170, n73171, n73172,
         n73173, n73174, n73175, n73176, n73177, n73178, n73179, n73180,
         n73181, n73182, n73183, n73184, n73185, n73186, n73187, n73188,
         n73189, n73190, n73191, n73192, n73193, n73194, n73195, n73196,
         n73197, n73198, n73199, n73200, n73201, n73202, n73203, n73204,
         n73205, n73206, n73207, n73208, n73209, n73210, n73211, n73212,
         n73213, n73214, n73215, n73216, n73217, n73218, n73219, n73220,
         n73221, n73222, n73223, n73224, n73225, n73226, n73227, n73228,
         n73229, n73230, n73231, n73232, n73233, n73234, n73235, n73236,
         n73237, n73238, n73239, n73240, n73241, n73242, n73243, n73244,
         n73245, n73246, n73247, n73248, n73249, n73250, n73251, n73252,
         n73253, n73254, n73255, n73256, n73257, n73258, n73259, n73260,
         n73261, n73262, n73263, n73264, n73265, n73266, n73267, n73268,
         n73269, n73270, n73271, n73272, n73273, n73274, n73275, n73276,
         n73277, n73278, n73279, n73280, n73281, n73282, n73283, n73284,
         n73285, n73286, n73287, n73288, n73289, n73290, n73291, n73292,
         n73293, n73294, n73295, n73296, n73297, n73298, n73299, n73300,
         n73301, n73302, n73303, n73304, n73305, n73306, n73307, n73308,
         n73309, n73310, n73311, n73312, n73313, n73314, n73315, n73316,
         n73317, n73318, n73319, n73320, n73321, n73322, n73323, n73324,
         n73325, n73326, n73327, n73328, n73329, n73330, n73331, n73332,
         n73333, n73334, n73335, n73336, n73337, n73338, n73339, n73340,
         n73341, n73342, n73343, n73344, n73345, n73346, n73347, n73348,
         n73349, n73350, n73351, n73352, n73353, n73354, n73355, n73356,
         n73357, n73358, n73359, n73360, n73361, n73362, n73363, n73364,
         n73365, n73366, n73367, n73368, n73369, n73370, n73371, n73372,
         n73373, n73374, n73375, n73376, n73377, n73378, n73379, n73380,
         n73381, n73382, n73383, n73384, n73385, n73386, n73387, n73388,
         n73389, n73390, n73391, n73392, n73393, n73394, n73395, n73396,
         n73397, n73398, n73399, n73400, n73401, n73402, n73403, n73404,
         n73405, n73406, n73407, n73408, n73409, n73410, n73411, n73412,
         n73413, n73414, n73415, n73416, n73417, n73418, n73419, n73420,
         n73421, n73422, n73423, n73424, n73425, n73426, n73427, n73428,
         n73429, n73430, n73431, n73432, n73433, n73434, n73435, n73436,
         n73437, n73438, n73439, n73440, n73441, n73442, n73443, n73444,
         n73445, n73446, n73447, n73448, n73449, n73450, n73451, n73452,
         n73453, n73454, n73455, n73456, n73457, n73458, n73459, n73460,
         n73461, n73462, n73463, n73464, n73465, n73466, n73467, n73468,
         n73469, n73470, n73471, n73472, n73473, n73474, n73475, n73476,
         n73477, n73478, n73479, n73480, n73481, n73482, n73483, n73484,
         n73485, n73486, n73487, n73488, n73489, n73490, n73491, n73492,
         n73493, n73494, n73495, n73496, n73497, n73498, n73499, n73500,
         n73501, n73502, n73503, n73504, n73505, n73506, n73507, n73508,
         n73509, n73510, n73511, n73512, n73513, n73514, n73515, n73516,
         n73517, n73518, n73519, n73520, n73521, n73522, n73523, n73524,
         n73525, n73526, n73527, n73528, n73529, n73530, n73531, n73532,
         n73533, n73534, n73535, n73536, n73537, n73538, n73539, n73540,
         n73541, n73542, n73543, n73544, n73545, n73546, n73547, n73548,
         n73549, n73550, n73551, n73552, n73553, n73554, n73555, n73556,
         n73557, n73558, n73559, n73560, n73561, n73562, n73563, n73564,
         n73565, n73566, n73567, n73568, n73569, n73570, n73571, n73572,
         n73573, n73574, n73575, n73576, n73577, n73578;
  wire   [31:1] u_csr_csr_mcycle_r;
  wire   [31:0] u_csr_csr_mcycle_q;
  wire   [1:0] u_mmu_state_q;
  wire   [31:12] u_mmu_pte_entry_q;
  wire   [27:12] u_mmu_request_addr_w;
  wire   [31:12] u_mmu_dtlb_va_addr_q;
  wire   [3:0] u_mmu_store_q;
  wire   [21:12] u_mmu_virt_addr_q;
  wire   [31:21] u_mmu_itlb_va_addr_q;
  wire   [31:1] opcode_pc_w;
  wire   [31:0] u_csr_csr_sepc_r;
  wire   [31:0] u_csr_csr_sepc_q;
  wire   [31:0] u_muldiv_dividend_q;
  wire   [62:1] u_muldiv_divisor_q;
  wire   [31:0] u_lsu_mem_addr_r;
  wire   [31:0] mmu_lsu_addr_w;
  wire   [31:0] u_csr_csr_stval_r;
  wire   [31:0] u_csr_csr_stval_q;
  wire   [31:0] u_muldiv_result_r;
  wire   [31:0] u_muldiv_mult_result_q;
  wire   [31:23] u_csr_csr_sr_r;
  wire   [17:0] u_csr_csr_sr_q;
  wire   [31:0] u_muldiv_q_mask_q;
  wire   [31:0] u_muldiv_quotient_q;
  wire   [4:0] writeback_muldiv_idx_w;
  wire   [31:1] u_decode_scoreboard_r;
  wire   [31:1] u_decode_scoreboard_q;
  wire   [63:0] u_fetch_skid_buffer_q;
  wire   [31:0] u_csr_csr_satp_r;
  wire   [31:12] u_mmu_itlb_entry_q;
  wire   [31:7] opcode_opcode_w;
  wire   [4:0] u_muldiv_rd_q;
  wire   [12:5] opcode_instr_w;
  wire   [31:0] u_csr_csr_mtvec_r;
  wire   [31:0] u_csr_csr_mtvec_q;
  wire   [31:0] u_csr_csr_mscratch_r;
  wire   [31:0] u_csr_csr_mscratch_q;
  wire   [31:27] u_csr_pc_m_q;
  wire   [4:0] u_csr_writeback_idx_q;
  wire   [15:0] u_csr_csr_medeleg_r;
  wire   [15:0] u_csr_csr_medeleg_q;
  wire   [15:0] u_csr_csr_mideleg_r;
  wire   [15:0] u_csr_csr_mideleg_q;
  wire   [31:0] u_csr_csr_sscratch_r;
  wire   [31:0] u_csr_csr_sscratch_q;
  wire   [31:0] u_csr_csr_stvec_r;
  wire   [31:0] u_csr_csr_stvec_q;
  wire   [4:0] writeback_exec_idx_w;
  wire   [3:0] u_csr_csr_scause_r;
  wire   [3:0] u_csr_csr_scause_q;
  wire   [3:0] u_csr_csr_mcause_r;
  wire   [3:0] u_csr_csr_mcause_q;
  wire   [31:0] u_csr_csr_mepc_r;
  wire   [31:0] u_csr_csr_mepc_q;
  wire   [31:2] arb_mmu_addr_w;
  wire   [31:0] u_exec_alu_p_w;
  wire   [31:0] writeback_exec_value_w;
  wire   [31:0] writeback_muldiv_value_w;
  wire   [31:0] u_csr_result_r;
  wire   [31:0] writeback_csr_value_w;
  assign mem_i_invalidate_o = 1'b0;

  DFFRX1 u_csr_csr_mcycle_q_reg_31_ ( .D(u_csr_csr_mcycle_r[31]), .CK(clk_i), 
        .RN(n44171), .QN(n37729) );
  DFFRX1 u_csr_csr_mcycle_q_reg_0_ ( .D(n8886), .CK(clk_i), .RN(n44171), .Q(
        u_csr_csr_mcycle_q[0]), .QN(n8886) );
  DFFRX1 u_csr_csr_mcycle_q_reg_1_ ( .D(u_csr_csr_mcycle_r[1]), .CK(clk_i), 
        .RN(n44171), .Q(u_csr_csr_mcycle_q[1]), .QN(n37343) );
  DFFRX1 u_csr_csr_mcycle_q_reg_2_ ( .D(u_csr_csr_mcycle_r[2]), .CK(clk_i), 
        .RN(n44170), .QN(n37563) );
  DFFRX1 u_csr_csr_mcycle_q_reg_3_ ( .D(u_csr_csr_mcycle_r[3]), .CK(clk_i), 
        .RN(n44170), .Q(u_csr_csr_mcycle_q[3]), .QN(n37693) );
  DFFRX1 u_csr_csr_mcycle_q_reg_4_ ( .D(u_csr_csr_mcycle_r[4]), .CK(clk_i), 
        .RN(n44170), .Q(u_csr_csr_mcycle_q[4]), .QN(n37721) );
  DFFRX1 u_csr_csr_mcycle_q_reg_5_ ( .D(u_csr_csr_mcycle_r[5]), .CK(clk_i), 
        .RN(n44170), .Q(u_csr_csr_mcycle_q[5]), .QN(n37345) );
  DFFRX1 u_csr_csr_mcycle_q_reg_6_ ( .D(u_csr_csr_mcycle_r[6]), .CK(clk_i), 
        .RN(n44170), .QN(n37569) );
  DFFRX1 u_csr_csr_mcycle_q_reg_7_ ( .D(u_csr_csr_mcycle_r[7]), .CK(clk_i), 
        .RN(n44170), .QN(n37346) );
  DFFRX1 u_csr_csr_mcycle_q_reg_8_ ( .D(u_csr_csr_mcycle_r[8]), .CK(clk_i), 
        .RN(n44170), .QN(n37571) );
  DFFRX1 u_csr_csr_mcycle_q_reg_9_ ( .D(u_csr_csr_mcycle_r[9]), .CK(clk_i), 
        .RN(n44170), .Q(u_csr_csr_mcycle_q[9]), .QN(n37694) );
  DFFRX1 u_csr_csr_mcycle_q_reg_10_ ( .D(u_csr_csr_mcycle_r[10]), .CK(clk_i), 
        .RN(n44170), .Q(u_csr_csr_mcycle_q[10]), .QN(n37711) );
  DFFRX1 u_csr_csr_mcycle_q_reg_11_ ( .D(u_csr_csr_mcycle_r[11]), .CK(clk_i), 
        .RN(n44170), .Q(u_csr_csr_mcycle_q[11]), .QN(n37347) );
  DFFRX1 u_csr_csr_mcycle_q_reg_12_ ( .D(u_csr_csr_mcycle_r[12]), .CK(clk_i), 
        .RN(n44170), .QN(n37574) );
  DFFRX1 u_csr_csr_mcycle_q_reg_13_ ( .D(u_csr_csr_mcycle_r[13]), .CK(clk_i), 
        .RN(n44170), .Q(u_csr_csr_mcycle_q[13]), .QN(n37692) );
  DFFRX1 u_csr_csr_mcycle_q_reg_14_ ( .D(u_csr_csr_mcycle_r[14]), .CK(clk_i), 
        .RN(n44170), .Q(u_csr_csr_mcycle_q[14]), .QN(n37712) );
  DFFRX1 u_csr_csr_mcycle_q_reg_15_ ( .D(u_csr_csr_mcycle_r[15]), .CK(clk_i), 
        .RN(n44170), .Q(u_csr_csr_mcycle_q[15]), .QN(n37348) );
  DFFRX1 u_csr_csr_mcycle_q_reg_16_ ( .D(u_csr_csr_mcycle_r[16]), .CK(clk_i), 
        .RN(n44170), .QN(n37578) );
  DFFRX1 u_csr_csr_mcycle_q_reg_17_ ( .D(u_csr_csr_mcycle_r[17]), .CK(clk_i), 
        .RN(n44170), .Q(u_csr_csr_mcycle_q[17]), .QN(n37689) );
  DFFRX1 u_csr_csr_mcycle_q_reg_18_ ( .D(u_csr_csr_mcycle_r[18]), .CK(clk_i), 
        .RN(n44170), .Q(u_csr_csr_mcycle_q[18]), .QN(n37696) );
  DFFRX1 u_csr_csr_mcycle_q_reg_19_ ( .D(u_csr_csr_mcycle_r[19]), .CK(clk_i), 
        .RN(n44170), .Q(u_csr_csr_mcycle_q[19]), .QN(n37349) );
  DFFRX1 u_csr_csr_mcycle_q_reg_20_ ( .D(u_csr_csr_mcycle_r[20]), .CK(clk_i), 
        .RN(n44169), .QN(n37585) );
  DFFRX1 u_csr_csr_mcycle_q_reg_21_ ( .D(u_csr_csr_mcycle_r[21]), .CK(clk_i), 
        .RN(n44169), .Q(u_csr_csr_mcycle_q[21]), .QN(n37690) );
  DFFRX1 u_csr_csr_mcycle_q_reg_22_ ( .D(u_csr_csr_mcycle_r[22]), .CK(clk_i), 
        .RN(n44169), .Q(u_csr_csr_mcycle_q[22]), .QN(n37697) );
  DFFRX1 u_csr_csr_mcycle_q_reg_23_ ( .D(u_csr_csr_mcycle_r[23]), .CK(clk_i), 
        .RN(n44169), .Q(u_csr_csr_mcycle_q[23]), .QN(n37350) );
  DFFRX1 u_csr_csr_mcycle_q_reg_24_ ( .D(u_csr_csr_mcycle_r[24]), .CK(clk_i), 
        .RN(n44169), .QN(n37588) );
  DFFRX1 u_csr_csr_mcycle_q_reg_25_ ( .D(u_csr_csr_mcycle_r[25]), .CK(clk_i), 
        .RN(n44169), .Q(u_csr_csr_mcycle_q[25]), .QN(n37691) );
  DFFRX1 u_csr_csr_mcycle_q_reg_26_ ( .D(u_csr_csr_mcycle_r[26]), .CK(clk_i), 
        .RN(n44169), .Q(u_csr_csr_mcycle_q[26]), .QN(n37698) );
  DFFRX1 u_csr_csr_mcycle_q_reg_27_ ( .D(u_csr_csr_mcycle_r[27]), .CK(clk_i), 
        .RN(n44169), .Q(u_csr_csr_mcycle_q[27]), .QN(n37352) );
  DFFRX1 u_csr_csr_mcycle_q_reg_28_ ( .D(u_csr_csr_mcycle_r[28]), .CK(clk_i), 
        .RN(n44169), .QN(n37598) );
  DFFRX1 u_csr_csr_mcycle_q_reg_29_ ( .D(u_csr_csr_mcycle_r[29]), .CK(clk_i), 
        .RN(n44169), .Q(u_csr_csr_mcycle_q[29]), .QN(n37695) );
  DFFRX1 u_csr_csr_mcycle_q_reg_30_ ( .D(u_csr_csr_mcycle_r[30]), .CK(clk_i), 
        .RN(n44169), .Q(u_csr_csr_mcycle_q[30]), .QN(n37699) );
  DFFRX1 u_mmu_state_q_reg_1_ ( .D(n8556), .CK(clk_i), .RN(n44250), .Q(
        u_mmu_state_q[1]), .QN(n37550) );
  DFFRX1 u_mmu_pte_entry_q_reg_1_ ( .D(u_mmu_N235), .CK(net1802), .RN(n44169), 
        .Q(u_mmu_pte_entry_q_1) );
  DFFRX1 u_mmu_pte_entry_q_reg_2_ ( .D(u_mmu_N236), .CK(net1802), .RN(n44169), 
        .Q(u_mmu_pte_entry_q_2) );
  DFFRX1 u_mmu_pte_entry_q_reg_3_ ( .D(u_mmu_N237), .CK(net1802), .RN(n44169), 
        .Q(u_mmu_pte_entry_q_3) );
  DFFRX1 u_mmu_pte_entry_q_reg_4_ ( .D(u_mmu_N238), .CK(net1802), .RN(n44169), 
        .Q(u_mmu_pte_entry_q_4) );
  DFFRX1 u_mmu_pte_entry_q_reg_22_ ( .D(u_mmu_N249), .CK(net1802), .RN(n44169), 
        .Q(u_mmu_pte_entry_q[22]) );
  DFFRX1 u_mmu_pte_entry_q_reg_23_ ( .D(u_mmu_N250), .CK(net1802), .RN(n44169), 
        .Q(u_mmu_pte_entry_q[23]) );
  DFFRX1 u_mmu_pte_entry_q_reg_24_ ( .D(n8550), .CK(clk_i), .RN(n44169), .Q(
        u_mmu_pte_entry_q[24]) );
  DFFRX1 u_mmu_pte_entry_q_reg_25_ ( .D(n8549), .CK(clk_i), .RN(n44168), .Q(
        u_mmu_pte_entry_q[25]) );
  DFFRX1 u_mmu_pte_entry_q_reg_26_ ( .D(n8548), .CK(clk_i), .RN(n44168), .Q(
        u_mmu_pte_entry_q[26]) );
  DFFRX1 u_mmu_pte_entry_q_reg_27_ ( .D(n8547), .CK(clk_i), .RN(n44168), .Q(
        u_mmu_pte_entry_q[27]) );
  DFFRX1 u_mmu_pte_entry_q_reg_28_ ( .D(n8546), .CK(clk_i), .RN(n44168), .Q(
        u_mmu_pte_entry_q[28]) );
  DFFRX1 u_mmu_pte_entry_q_reg_29_ ( .D(n8545), .CK(clk_i), .RN(n44168), .Q(
        u_mmu_pte_entry_q[29]) );
  DFFRX1 u_mmu_pte_entry_q_reg_30_ ( .D(n8544), .CK(clk_i), .RN(n44168), .Q(
        u_mmu_pte_entry_q[30]) );
  DFFRX1 u_mmu_pte_entry_q_reg_31_ ( .D(n8543), .CK(clk_i), .RN(n44168), .Q(
        u_mmu_pte_entry_q[31]) );
  DFFRX1 u_mmu_dtlb_va_addr_q_reg_27_ ( .D(n8445), .CK(clk_i), .RN(n44206), 
        .Q(u_mmu_dtlb_va_addr_q[27]) );
  DFFRX1 u_arb_read_hold_q_reg ( .D(n8558), .CK(clk_i), .RN(n44168), .Q(
        u_arb_read_hold_q), .QN(n37448) );
  DFFRX1 u_arb_src_mmu_q_reg ( .D(n8557), .CK(clk_i), .RN(n44168), .Q(
        u_arb_src_mmu_q) );
  DFFRX1 u_mmu_store_q_reg_3_ ( .D(n8539), .CK(clk_i), .RN(n44205), .Q(
        u_mmu_store_q[3]), .QN(n37430) );
  DFFRX1 u_mmu_itlb_va_addr_q_reg_29_ ( .D(n8444), .CK(clk_i), .RN(n44180), 
        .Q(u_mmu_itlb_va_addr_q[29]) );
  DFFRX1 u_fetch_fetch_pc_q_reg_31_ ( .D(u_fetch_N80), .CK(n37883), .RN(n44183), .QN(n1757) );
  DFFRX1 u_fetch_fetch_pc_q_reg_15_ ( .D(u_fetch_N64), .CK(n37882), .RN(n44107), .QN(n1773) );
  DFFRX1 u_fetch_fetch_pc_q_reg_16_ ( .D(u_fetch_N65), .CK(n37883), .RN(n44107), .QN(n1774) );
  DFFRX1 u_fetch_fetch_pc_q_reg_17_ ( .D(u_fetch_N66), .CK(n37883), .RN(n44108), .QN(n1775) );
  DFFRX1 u_fetch_fetch_pc_q_reg_18_ ( .D(u_fetch_N67), .CK(n37883), .RN(n44108), .QN(n1776) );
  DFFRX1 u_fetch_fetch_pc_q_reg_19_ ( .D(u_fetch_N68), .CK(n37883), .RN(n44109), .QN(n1777) );
  DFFRX1 u_fetch_fetch_pc_q_reg_20_ ( .D(u_fetch_N69), .CK(n37883), .RN(n44109), .QN(n1778) );
  DFFRX1 u_fetch_fetch_pc_q_reg_21_ ( .D(u_fetch_N70), .CK(n37883), .RN(n44110), .QN(n1779) );
  DFFRX1 u_fetch_fetch_pc_q_reg_22_ ( .D(u_fetch_N71), .CK(n37883), .RN(n44110), .QN(n1780) );
  DFFRX1 u_fetch_fetch_pc_q_reg_23_ ( .D(u_fetch_N72), .CK(n37883), .RN(n44111), .QN(n1781) );
  DFFRX1 u_fetch_fetch_pc_q_reg_24_ ( .D(u_fetch_N73), .CK(n37883), .RN(n44188), .QN(n1782) );
  DFFRX1 u_fetch_fetch_pc_q_reg_25_ ( .D(u_fetch_N74), .CK(n37883), .RN(n44188), .QN(n1783) );
  DFFRX1 u_fetch_fetch_pc_q_reg_26_ ( .D(u_fetch_N75), .CK(n37883), .RN(n44189), .QN(n1784) );
  DFFRX1 u_fetch_fetch_pc_q_reg_27_ ( .D(u_fetch_N76), .CK(n37883), .RN(n44191), .QN(n1785) );
  DFFRX1 u_fetch_fetch_pc_q_reg_28_ ( .D(u_fetch_N77), .CK(n37883), .RN(n44193), .QN(n1786) );
  DFFRX1 u_fetch_fetch_pc_q_reg_29_ ( .D(u_fetch_N78), .CK(n37883), .RN(n44196), .QN(n1787) );
  DFFRX1 u_fetch_fetch_pc_q_reg_30_ ( .D(u_fetch_N79), .CK(n37883), .RN(n44182), .QN(n1788) );
  DFFRX1 u_decode_u_regfile_reg_r24_q_reg_30_ ( .D(u_decode_u_regfile_N981), 
        .CK(n37881), .RN(n44180), .Q(n1789) );
  DFFRX1 u_decode_u_regfile_reg_r23_q_reg_30_ ( .D(u_decode_u_regfile_N944), 
        .CK(n37880), .RN(n44181), .Q(n1790) );
  DFFRX1 u_decode_u_regfile_reg_r25_q_reg_0_ ( .D(u_decode_u_regfile_N988), 
        .CK(n37879), .RN(n44205), .Q(n1791), .QN(n37303) );
  DFFRX1 u_muldiv_dividend_q_reg_0_ ( .D(u_muldiv_N232), .CK(net1908), .RN(
        n44168), .Q(u_muldiv_dividend_q[0]) );
  DFFRX1 u_decode_u_regfile_reg_r24_q_reg_31_ ( .D(u_decode_u_regfile_N982), 
        .CK(n37881), .RN(n44187), .Q(n1792), .QN(n36819) );
  DFFRX1 u_decode_u_regfile_reg_r24_q_reg_15_ ( .D(u_decode_u_regfile_N966), 
        .CK(n37878), .RN(n44124), .Q(n1793), .QN(n37163) );
  DFFRX1 u_muldiv_dividend_q_reg_15_ ( .D(u_muldiv_N247), .CK(net1908), .RN(
        n44168), .Q(u_muldiv_dividend_q[15]), .QN(n37446) );
  DFFRX1 u_decode_u_regfile_reg_r23_q_reg_15_ ( .D(u_decode_u_regfile_N929), 
        .CK(n37877), .RN(n44125), .Q(n1794) );
  DFFRX1 u_muldiv_divisor_q_reg_46_ ( .D(u_muldiv_N311), .CK(net1893), .RN(
        n44168), .Q(u_muldiv_divisor_q[46]) );
  DFFRX1 u_muldiv_divisor_q_reg_45_ ( .D(u_muldiv_N310), .CK(net1893), .RN(
        n44168), .Q(u_muldiv_divisor_q[45]) );
  DFFRX1 u_muldiv_divisor_q_reg_44_ ( .D(u_muldiv_N309), .CK(net1893), .RN(
        n44168), .Q(u_muldiv_divisor_q[44]) );
  DFFRX1 u_muldiv_divisor_q_reg_43_ ( .D(u_muldiv_N308), .CK(net1893), .RN(
        n44168), .Q(u_muldiv_divisor_q[43]), .QN(n37590) );
  DFFRX1 u_muldiv_divisor_q_reg_42_ ( .D(u_muldiv_N307), .CK(net1893), .RN(
        n44168), .Q(u_muldiv_divisor_q[42]) );
  DFFRX1 u_muldiv_divisor_q_reg_41_ ( .D(u_muldiv_N306), .CK(net1893), .RN(
        n44167), .Q(u_muldiv_divisor_q[41]) );
  DFFRX1 u_muldiv_divisor_q_reg_40_ ( .D(u_muldiv_N305), .CK(net1893), .RN(
        n44167), .Q(u_muldiv_divisor_q[40]) );
  DFFRX1 u_muldiv_divisor_q_reg_39_ ( .D(u_muldiv_N304), .CK(net1893), .RN(
        n44167), .Q(u_muldiv_divisor_q[39]) );
  DFFRX1 u_muldiv_divisor_q_reg_38_ ( .D(u_muldiv_N303), .CK(net1893), .RN(
        n44167), .Q(u_muldiv_divisor_q[38]) );
  DFFRX1 u_muldiv_divisor_q_reg_37_ ( .D(u_muldiv_N302), .CK(net1893), .RN(
        n44167), .Q(u_muldiv_divisor_q[37]) );
  DFFRX1 u_muldiv_divisor_q_reg_36_ ( .D(u_muldiv_N301), .CK(net1893), .RN(
        n44167), .Q(u_muldiv_divisor_q[36]) );
  DFFRX1 u_muldiv_divisor_q_reg_35_ ( .D(u_muldiv_N300), .CK(net1893), .RN(
        n44167), .Q(u_muldiv_divisor_q[35]) );
  DFFRX1 u_muldiv_divisor_q_reg_34_ ( .D(u_muldiv_N299), .CK(net1893), .RN(
        n44167), .Q(u_muldiv_divisor_q[34]) );
  DFFRX1 u_muldiv_divisor_q_reg_33_ ( .D(u_muldiv_N298), .CK(net1893), .RN(
        n44167), .Q(u_muldiv_divisor_q[33]) );
  DFFRX1 u_muldiv_divisor_q_reg_32_ ( .D(u_muldiv_N297), .CK(net1893), .RN(
        n44167), .Q(u_muldiv_divisor_q[32]), .QN(n37591) );
  DFFRX1 u_muldiv_divisor_q_reg_31_ ( .D(u_muldiv_N296), .CK(net1888), .RN(
        n44167), .Q(u_muldiv_divisor_q[31]) );
  DFFRX1 u_muldiv_divisor_q_reg_30_ ( .D(u_muldiv_N295), .CK(net1888), .RN(
        n44167), .Q(u_muldiv_divisor_q[30]), .QN(n37582) );
  DFFRX1 u_muldiv_divisor_q_reg_29_ ( .D(u_muldiv_N294), .CK(net1888), .RN(
        n44167), .Q(u_muldiv_divisor_q[29]), .QN(n37583) );
  DFFRX1 u_muldiv_divisor_q_reg_28_ ( .D(u_muldiv_N293), .CK(net1888), .RN(
        n44167), .Q(u_muldiv_divisor_q[28]), .QN(n37576) );
  DFFRX1 u_muldiv_divisor_q_reg_27_ ( .D(u_muldiv_N292), .CK(net1888), .RN(
        n44167), .Q(u_muldiv_divisor_q[27]), .QN(n37573) );
  DFFRX1 u_muldiv_divisor_q_reg_26_ ( .D(u_muldiv_N291), .CK(net1888), .RN(
        n44167), .Q(u_muldiv_divisor_q[26]), .QN(n42553) );
  DFFRX1 u_muldiv_divisor_q_reg_25_ ( .D(u_muldiv_N290), .CK(net1888), .RN(
        n44167), .Q(u_muldiv_divisor_q[25]), .QN(n37564) );
  DFFRX1 u_muldiv_divisor_q_reg_24_ ( .D(u_muldiv_N289), .CK(net1888), .RN(
        n44166), .Q(u_muldiv_divisor_q[24]), .QN(n37559) );
  DFFRX1 u_muldiv_divisor_q_reg_23_ ( .D(u_muldiv_N288), .CK(net1888), .RN(
        n44166), .Q(u_muldiv_divisor_q[23]), .QN(n37557) );
  DFFRX1 u_muldiv_divisor_q_reg_22_ ( .D(u_muldiv_N287), .CK(net1888), .RN(
        n44166), .Q(u_muldiv_divisor_q[22]), .QN(n42551) );
  DFFRX1 u_muldiv_divisor_q_reg_21_ ( .D(u_muldiv_N286), .CK(net1888), .RN(
        n44166), .Q(u_muldiv_divisor_q[21]), .QN(n37551) );
  DFFRX1 u_muldiv_divisor_q_reg_20_ ( .D(u_muldiv_N285), .CK(net1888), .RN(
        n44166), .Q(u_muldiv_divisor_q[20]), .QN(n37543) );
  DFFRX1 u_muldiv_divisor_q_reg_19_ ( .D(u_muldiv_N284), .CK(net1888), .RN(
        n44166), .Q(u_muldiv_divisor_q[19]), .QN(n37538) );
  DFFRX1 u_muldiv_divisor_q_reg_18_ ( .D(u_muldiv_N283), .CK(net1888), .RN(
        n44166), .Q(u_muldiv_divisor_q[18]), .QN(n42549) );
  DFFRX1 u_muldiv_divisor_q_reg_17_ ( .D(u_muldiv_N282), .CK(net1888), .RN(
        n44166), .Q(u_muldiv_divisor_q[17]), .QN(n37453) );
  DFFRX1 u_muldiv_divisor_q_reg_16_ ( .D(u_muldiv_N281), .CK(net1888), .RN(
        n44166), .Q(u_muldiv_divisor_q[16]), .QN(n37452) );
  DFFRX1 u_muldiv_divisor_q_reg_15_ ( .D(u_muldiv_N280), .CK(net1883), .RN(
        n44166), .Q(u_muldiv_divisor_q[15]), .QN(n37447) );
  DFFRX1 u_muldiv_divisor_q_reg_14_ ( .D(u_muldiv_N279), .CK(net1883), .RN(
        n44166), .Q(u_muldiv_divisor_q[14]), .QN(n42547) );
  DFFRX1 u_muldiv_divisor_q_reg_13_ ( .D(u_muldiv_N278), .CK(net1883), .RN(
        n44166), .Q(u_muldiv_divisor_q[13]), .QN(n37443) );
  DFFRX1 u_muldiv_divisor_q_reg_12_ ( .D(u_muldiv_N277), .CK(net1883), .RN(
        n44166), .Q(u_muldiv_divisor_q[12]), .QN(n37442) );
  DFFRX1 u_muldiv_divisor_q_reg_11_ ( .D(u_muldiv_N276), .CK(net1883), .RN(
        n44166), .Q(u_muldiv_divisor_q[11]), .QN(n37440) );
  DFFRX1 u_muldiv_divisor_q_reg_10_ ( .D(u_muldiv_N275), .CK(net1883), .RN(
        n44166), .Q(u_muldiv_divisor_q[10]), .QN(n42555) );
  DFFRX1 u_muldiv_divisor_q_reg_9_ ( .D(u_muldiv_N274), .CK(net1883), .RN(
        n44166), .Q(u_muldiv_divisor_q[9]), .QN(n37432) );
  DFFRX1 u_muldiv_divisor_q_reg_8_ ( .D(u_muldiv_N273), .CK(net1883), .RN(
        n44166), .Q(u_muldiv_divisor_q[8]), .QN(n37429) );
  DFFRX1 u_muldiv_divisor_q_reg_7_ ( .D(u_muldiv_N272), .CK(net1883), .RN(
        n44166), .Q(u_muldiv_divisor_q[7]), .QN(n37427) );
  DFFRX1 u_muldiv_divisor_q_reg_6_ ( .D(u_muldiv_N271), .CK(net1883), .RN(
        n44165), .Q(u_muldiv_divisor_q[6]), .QN(n37424) );
  DFFRX1 u_muldiv_divisor_q_reg_5_ ( .D(u_muldiv_N270), .CK(net1883), .RN(
        n44165), .Q(u_muldiv_divisor_q[5]), .QN(n37422) );
  DFFRX1 u_muldiv_divisor_q_reg_4_ ( .D(u_muldiv_N269), .CK(net1883), .RN(
        n44165), .Q(u_muldiv_divisor_q[4]), .QN(n37421) );
  DFFRX1 u_muldiv_divisor_q_reg_3_ ( .D(u_muldiv_N268), .CK(net1883), .RN(
        n44165), .Q(u_muldiv_divisor_q[3]), .QN(n37438) );
  DFFRX1 u_muldiv_divisor_q_reg_2_ ( .D(u_muldiv_N267), .CK(net1883), .RN(
        n44165), .Q(u_muldiv_divisor_q[2]), .QN(n37435) );
  DFFRX1 u_muldiv_divisor_q_reg_1_ ( .D(u_muldiv_N266), .CK(net1883), .RN(
        n44165), .QN(n37419) );
  DFFRX1 u_muldiv_divisor_q_reg_0_ ( .D(u_muldiv_N265), .CK(net1883), .RN(
        n44165), .QN(n37418) );
  DFFRX1 u_muldiv_dividend_q_reg_14_ ( .D(u_muldiv_N246), .CK(net1908), .RN(
        n44165), .Q(u_muldiv_dividend_q[14]), .QN(n37445) );
  DFFRX1 u_decode_u_regfile_reg_r24_q_reg_14_ ( .D(u_decode_u_regfile_N965), 
        .CK(n37878), .RN(n44140), .Q(n1796), .QN(n37179) );
  DFFRX1 u_lsu_mem_addr_q_reg_14_ ( .D(u_lsu_mem_addr_r[14]), .CK(n37876), 
        .RN(n44186), .Q(mmu_lsu_addr_w[14]), .QN(n8300) );
  DFFRX1 u_mmu_lsu_in_addr_q_reg_14_ ( .D(mmu_lsu_addr_w[14]), .CK(n37875), 
        .RN(n44186), .QN(n1797) );
  DFFRX1 u_decode_u_regfile_reg_r23_q_reg_14_ ( .D(u_decode_u_regfile_N928), 
        .CK(n37877), .RN(n44096), .Q(n1798) );
  DFFRX1 u_decode_u_regfile_reg_r23_q_reg_31_ ( .D(u_decode_u_regfile_N945), 
        .CK(n37880), .RN(n44204), .Q(n1799) );
  DFFRX1 u_decode_u_regfile_reg_r24_q_reg_29_ ( .D(u_decode_u_regfile_N980), 
        .CK(n37881), .RN(n44194), .Q(n1800), .QN(n37038) );
  DFFRX1 u_lsu_mem_addr_q_reg_29_ ( .D(u_lsu_mem_addr_r[29]), .CK(n37874), 
        .RN(n44184), .Q(n56367), .QN(n8332) );
  DFFRX1 u_mmu_lsu_in_addr_q_reg_29_ ( .D(n56367), .CK(n37873), .RN(n44206), 
        .QN(n1801) );
  DFFRX1 u_decode_u_regfile_reg_r23_q_reg_29_ ( .D(u_decode_u_regfile_N943), 
        .CK(n37880), .RN(n44195), .Q(n1802) );
  DFFRX1 u_decode_u_regfile_reg_r24_q_reg_28_ ( .D(u_decode_u_regfile_N979), 
        .CK(n37881), .RN(n44191), .Q(n1803), .QN(n37030) );
  DFFRX1 u_decode_u_regfile_reg_r23_q_reg_28_ ( .D(u_decode_u_regfile_N942), 
        .CK(n37880), .RN(n44193), .Q(n1804) );
  DFFRX1 u_decode_u_regfile_reg_r25_q_reg_5_ ( .D(u_decode_u_regfile_N993), 
        .CK(n37879), .RN(n44145), .Q(n1806), .QN(n37288) );
  DFFRX1 u_muldiv_dividend_q_reg_5_ ( .D(u_muldiv_N237), .CK(net1908), .RN(
        n44165), .Q(u_muldiv_dividend_q[5]) );
  DFFRX1 u_decode_u_regfile_reg_r24_q_reg_5_ ( .D(u_decode_u_regfile_N956), 
        .CK(n37878), .RN(n44145), .Q(n1807), .QN(n37289) );
  DFFRX1 u_csr_branch_target_q_reg_31_ ( .D(u_csr_N3696), .CK(clk_i), .RN(
        n44183), .Q(n56613) );
  DFFRX1 u_decode_u_regfile_reg_r24_q_reg_17_ ( .D(u_decode_u_regfile_N968), 
        .CK(n37881), .RN(n44098), .Q(n1808), .QN(n37166) );
  DFFRX1 u_decode_u_regfile_reg_r24_q_reg_24_ ( .D(u_decode_u_regfile_N975), 
        .CK(n37881), .RN(n44095), .Q(n1809), .QN(n42477) );
  DFFRX1 u_decode_u_regfile_reg_r24_q_reg_25_ ( .D(u_decode_u_regfile_N976), 
        .CK(n37881), .RN(n44113), .Q(n1810), .QN(n42488) );
  DFFRX1 u_decode_u_regfile_reg_r24_q_reg_27_ ( .D(u_decode_u_regfile_N978), 
        .CK(n37881), .RN(n44189), .Q(n1811), .QN(n37031) );
  DFFRX1 u_decode_u_regfile_reg_r24_q_reg_13_ ( .D(u_decode_u_regfile_N964), 
        .CK(n37878), .RN(n44122), .Q(n1812), .QN(n37191) );
  DFFRX1 u_decode_u_regfile_reg_r25_q_reg_1_ ( .D(u_decode_u_regfile_N989), 
        .CK(n37879), .RN(n44121), .QN(n36802) );
  DFFRX1 u_muldiv_dividend_q_reg_1_ ( .D(u_muldiv_N233), .CK(net1908), .RN(
        n44165), .Q(u_muldiv_dividend_q[1]) );
  DFFRX1 u_decode_u_regfile_reg_r24_q_reg_1_ ( .D(u_decode_u_regfile_N952), 
        .CK(n37878), .RN(n44121), .QN(n36860) );
  DFFRX1 u_decode_u_regfile_reg_r25_q_reg_4_ ( .D(u_decode_u_regfile_N992), 
        .CK(n37879), .RN(n44146), .Q(n1815), .QN(n37292) );
  DFFRX1 u_muldiv_dividend_q_reg_4_ ( .D(u_muldiv_N236), .CK(net1908), .RN(
        n44165), .Q(u_muldiv_dividend_q[4]), .QN(n37420) );
  DFFRX1 u_decode_u_regfile_reg_r24_q_reg_4_ ( .D(u_decode_u_regfile_N955), 
        .CK(n37878), .RN(n44146), .Q(n1816), .QN(n37293) );
  DFFRX1 u_decode_u_regfile_reg_r25_q_reg_8_ ( .D(u_decode_u_regfile_N996), 
        .CK(n37879), .RN(n44126), .Q(n1817), .QN(n37247) );
  DFFRX1 u_decode_u_regfile_reg_r24_q_reg_12_ ( .D(u_decode_u_regfile_N963), 
        .CK(n37878), .RN(n44138), .Q(n1818), .QN(n37213) );
  DFFRX1 u_decode_u_regfile_reg_r24_q_reg_18_ ( .D(u_decode_u_regfile_N969), 
        .CK(n37881), .RN(n44100), .Q(n1819), .QN(n37126) );
  DFFRX1 u_decode_u_regfile_reg_r24_q_reg_26_ ( .D(u_decode_u_regfile_N977), 
        .CK(n37881), .RN(n44114), .Q(n1820) );
  DFFRX1 u_decode_u_regfile_reg_r25_q_reg_7_ ( .D(u_decode_u_regfile_N995), 
        .CK(n37879), .RN(n44141), .Q(n1821), .QN(n37212) );
  DFFRX1 u_decode_u_regfile_reg_r24_q_reg_21_ ( .D(u_decode_u_regfile_N972), 
        .CK(n37881), .RN(n44089), .Q(n1822), .QN(n37133) );
  DFFRX1 u_decode_u_regfile_reg_r24_q_reg_16_ ( .D(u_decode_u_regfile_N967), 
        .CK(n37881), .RN(n44097), .Q(n1823), .QN(n37171) );
  DFFRX1 u_decode_u_regfile_reg_r24_q_reg_22_ ( .D(u_decode_u_regfile_N973), 
        .CK(n37881), .RN(n44091), .Q(n1824), .QN(n37098) );
  DFFRX1 u_decode_u_regfile_reg_r24_q_reg_23_ ( .D(u_decode_u_regfile_N974), 
        .CK(n37881), .RN(n44093), .Q(n1825) );
  DFFRX1 u_decode_u_regfile_reg_r25_q_reg_9_ ( .D(u_decode_u_regfile_N997), 
        .CK(n37879), .RN(n44133), .Q(n1826), .QN(n37267) );
  DFFRX1 u_decode_u_regfile_reg_r25_q_reg_3_ ( .D(u_decode_u_regfile_N991), 
        .CK(n37879), .RN(n44130), .QN(n37026) );
  DFFRX1 u_muldiv_dividend_q_reg_3_ ( .D(u_muldiv_N235), .CK(net1908), .RN(
        n44165), .Q(u_muldiv_dividend_q[3]), .QN(n37326) );
  DFFRX1 u_decode_u_regfile_reg_r24_q_reg_3_ ( .D(u_decode_u_regfile_N954), 
        .CK(n37878), .RN(n44130), .QN(n37091) );
  DFFRX1 u_decode_u_regfile_reg_r24_q_reg_20_ ( .D(u_decode_u_regfile_N971), 
        .CK(n37881), .RN(n44088), .Q(n1829) );
  DFFRX1 u_decode_u_regfile_reg_r25_q_reg_10_ ( .D(u_decode_u_regfile_N998), 
        .CK(n37879), .RN(n44135), .Q(n1830), .QN(n37260) );
  DFFRX1 u_decode_u_regfile_reg_r25_q_reg_2_ ( .D(u_decode_u_regfile_N990), 
        .CK(n37879), .RN(n44132), .Q(n1831), .QN(n37310) );
  DFFRX1 u_muldiv_dividend_q_reg_2_ ( .D(u_muldiv_N234), .CK(net1908), .RN(
        n44165), .Q(u_muldiv_dividend_q[2]), .QN(n37325) );
  DFFRX1 u_decode_u_regfile_reg_r24_q_reg_2_ ( .D(u_decode_u_regfile_N953), 
        .CK(n37878), .RN(n44132), .Q(n1832), .QN(n37312) );
  DFFRX1 u_decode_u_regfile_reg_r25_q_reg_6_ ( .D(u_decode_u_regfile_N994), 
        .CK(n37879), .RN(n44143), .Q(n1833), .QN(n37278) );
  DFFRX1 u_decode_u_regfile_reg_r24_q_reg_19_ ( .D(u_decode_u_regfile_N970), 
        .CK(n37881), .RN(n44102), .Q(n1834) );
  DFFRX1 u_decode_u_regfile_reg_r25_q_reg_11_ ( .D(u_decode_u_regfile_N999), 
        .CK(n37879), .RN(n44137), .Q(n1835), .QN(n37227) );
  DFFRX1 u_csr_csr_sr_q_reg_11_ ( .D(u_csr_csr_sr_r_11), .CK(clk_i), .RN(
        n44165), .Q(u_csr_csr_sr_q[11]), .QN(n37688) );
  DFFRX1 u_csr_csr_sr_q_reg_12_ ( .D(u_csr_csr_sr_r_12), .CK(clk_i), .RN(
        n44164), .Q(u_csr_csr_sr_q[12]), .QN(n37749) );
  DFFRX1 u_muldiv_div_busy_q_reg ( .D(u_muldiv_N264), .CK(clk_i), .RN(n44209), 
        .Q(u_muldiv_div_busy_q), .QN(n37436) );
  DFFRX1 u_muldiv_q_mask_q_reg_31_ ( .D(n8536), .CK(clk_i), .RN(n44164), .Q(
        u_muldiv_q_mask_q[31]) );
  DFFRX1 u_muldiv_q_mask_q_reg_30_ ( .D(n8522), .CK(clk_i), .RN(n44164), .Q(
        u_muldiv_q_mask_q[30]) );
  DFFRX1 u_muldiv_q_mask_q_reg_29_ ( .D(n8523), .CK(clk_i), .RN(n44164), .Q(
        u_muldiv_q_mask_q[29]) );
  DFFRX1 u_muldiv_q_mask_q_reg_28_ ( .D(n8524), .CK(clk_i), .RN(n44164), .Q(
        u_muldiv_q_mask_q[28]) );
  DFFRX1 u_muldiv_q_mask_q_reg_27_ ( .D(n8525), .CK(clk_i), .RN(n44164), .Q(
        u_muldiv_q_mask_q[27]) );
  DFFRX1 u_muldiv_q_mask_q_reg_26_ ( .D(n8526), .CK(clk_i), .RN(n44164), .Q(
        u_muldiv_q_mask_q[26]) );
  DFFRX1 u_muldiv_q_mask_q_reg_25_ ( .D(n8527), .CK(clk_i), .RN(n44164), .Q(
        u_muldiv_q_mask_q[25]) );
  DFFRX1 u_muldiv_q_mask_q_reg_24_ ( .D(n8528), .CK(clk_i), .RN(n44164), .Q(
        u_muldiv_q_mask_q[24]) );
  DFFRX1 u_muldiv_q_mask_q_reg_23_ ( .D(n8529), .CK(clk_i), .RN(n44164), .Q(
        u_muldiv_q_mask_q[23]) );
  DFFRX1 u_muldiv_q_mask_q_reg_22_ ( .D(n8530), .CK(clk_i), .RN(n44164), .Q(
        u_muldiv_q_mask_q[22]) );
  DFFRX1 u_muldiv_q_mask_q_reg_21_ ( .D(n8531), .CK(clk_i), .RN(n44164), .Q(
        u_muldiv_q_mask_q[21]) );
  DFFRX1 u_muldiv_q_mask_q_reg_20_ ( .D(n8532), .CK(clk_i), .RN(n44164), .Q(
        u_muldiv_q_mask_q[20]) );
  DFFRX1 u_muldiv_q_mask_q_reg_19_ ( .D(n8533), .CK(clk_i), .RN(n44164), .Q(
        u_muldiv_q_mask_q[19]) );
  DFFRX1 u_muldiv_q_mask_q_reg_18_ ( .D(n8534), .CK(clk_i), .RN(n44164), .Q(
        u_muldiv_q_mask_q[18]) );
  DFFRX1 u_muldiv_q_mask_q_reg_17_ ( .D(n8535), .CK(clk_i), .RN(n44164), .Q(
        u_muldiv_q_mask_q[17]) );
  DFFRX1 u_muldiv_q_mask_q_reg_16_ ( .D(n863), .CK(net1903), .RN(n44164), .Q(
        u_muldiv_q_mask_q[16]) );
  DFFRX1 u_muldiv_q_mask_q_reg_15_ ( .D(n862), .CK(net1903), .RN(n44164), .Q(
        u_muldiv_q_mask_q[15]) );
  DFFRX1 u_muldiv_q_mask_q_reg_14_ ( .D(n861), .CK(net1903), .RN(n44163), .Q(
        u_muldiv_q_mask_q[14]) );
  DFFRX1 u_muldiv_q_mask_q_reg_13_ ( .D(n860), .CK(net1903), .RN(n44163), .Q(
        u_muldiv_q_mask_q[13]) );
  DFFRX1 u_muldiv_q_mask_q_reg_12_ ( .D(n859), .CK(net1903), .RN(n44163), .Q(
        u_muldiv_q_mask_q[12]) );
  DFFRX1 u_muldiv_q_mask_q_reg_11_ ( .D(n858), .CK(net1903), .RN(n44163), .Q(
        u_muldiv_q_mask_q[11]) );
  DFFRX1 u_muldiv_q_mask_q_reg_10_ ( .D(n857), .CK(net1903), .RN(n44163), .Q(
        u_muldiv_q_mask_q[10]) );
  DFFRX1 u_muldiv_q_mask_q_reg_9_ ( .D(n856), .CK(net1903), .RN(n44167), .Q(
        u_muldiv_q_mask_q[9]) );
  DFFRX1 u_muldiv_q_mask_q_reg_8_ ( .D(n855), .CK(net1903), .RN(n44179), .Q(
        u_muldiv_q_mask_q[8]) );
  DFFRX1 u_muldiv_q_mask_q_reg_7_ ( .D(n854), .CK(net1903), .RN(n44179), .Q(
        u_muldiv_q_mask_q[7]) );
  DFFRX1 u_muldiv_q_mask_q_reg_6_ ( .D(n853), .CK(net1903), .RN(n44179), .Q(
        u_muldiv_q_mask_q[6]) );
  DFFRX1 u_muldiv_q_mask_q_reg_5_ ( .D(n852), .CK(net1903), .RN(n44179), .Q(
        u_muldiv_q_mask_q[5]) );
  DFFRX1 u_muldiv_q_mask_q_reg_4_ ( .D(n851), .CK(net1903), .RN(n44179), .Q(
        u_muldiv_q_mask_q[4]) );
  DFFRX1 u_muldiv_q_mask_q_reg_3_ ( .D(n850), .CK(net1903), .RN(n44179), .Q(
        u_muldiv_q_mask_q[3]) );
  DFFRX1 u_muldiv_q_mask_q_reg_2_ ( .D(n849), .CK(net1903), .RN(n44179), .Q(
        u_muldiv_q_mask_q[2]) );
  DFFRX1 u_muldiv_q_mask_q_reg_1_ ( .D(n848), .CK(net1903), .RN(n44179), .Q(
        u_muldiv_q_mask_q[1]) );
  DFFRX1 u_muldiv_q_mask_q_reg_0_ ( .D(n847), .CK(net1898), .RN(n44179), .Q(
        u_muldiv_q_mask_q[0]) );
  DFFRX1 u_muldiv_quotient_q_reg_0_ ( .D(u_muldiv_N328), .CK(net1918), .RN(
        n44179), .Q(u_muldiv_quotient_q[0]) );
  DFFRX1 u_muldiv_quotient_q_reg_1_ ( .D(u_muldiv_N329), .CK(net1918), .RN(
        n44179), .Q(u_muldiv_quotient_q[1]) );
  DFFRX1 u_muldiv_quotient_q_reg_2_ ( .D(u_muldiv_N330), .CK(net1918), .RN(
        n44179), .Q(u_muldiv_quotient_q[2]) );
  DFFRX1 u_muldiv_quotient_q_reg_3_ ( .D(u_muldiv_N331), .CK(net1918), .RN(
        n44179), .Q(u_muldiv_quotient_q[3]) );
  DFFRX1 u_muldiv_quotient_q_reg_4_ ( .D(u_muldiv_N332), .CK(net1918), .RN(
        n44179), .Q(u_muldiv_quotient_q[4]) );
  DFFRX1 u_muldiv_quotient_q_reg_5_ ( .D(u_muldiv_N333), .CK(net1918), .RN(
        n44179), .Q(u_muldiv_quotient_q[5]) );
  DFFRX1 u_muldiv_quotient_q_reg_6_ ( .D(u_muldiv_N334), .CK(net1918), .RN(
        n44179), .Q(u_muldiv_quotient_q[6]) );
  DFFRX1 u_muldiv_quotient_q_reg_7_ ( .D(u_muldiv_N335), .CK(net1918), .RN(
        n44179), .Q(u_muldiv_quotient_q[7]) );
  DFFRX1 u_muldiv_quotient_q_reg_8_ ( .D(u_muldiv_N336), .CK(net1918), .RN(
        n44178), .Q(u_muldiv_quotient_q[8]) );
  DFFRX1 u_muldiv_quotient_q_reg_9_ ( .D(u_muldiv_N337), .CK(net1918), .RN(
        n44178), .Q(u_muldiv_quotient_q[9]) );
  DFFRX1 u_muldiv_quotient_q_reg_10_ ( .D(u_muldiv_N338), .CK(net1918), .RN(
        n44178), .Q(u_muldiv_quotient_q[10]) );
  DFFRX1 u_muldiv_quotient_q_reg_11_ ( .D(u_muldiv_N339), .CK(net1918), .RN(
        n44178), .Q(u_muldiv_quotient_q[11]) );
  DFFRX1 u_muldiv_quotient_q_reg_12_ ( .D(u_muldiv_N340), .CK(net1918), .RN(
        n44178), .Q(u_muldiv_quotient_q[12]) );
  DFFRX1 u_muldiv_quotient_q_reg_13_ ( .D(u_muldiv_N341), .CK(net1918), .RN(
        n44178), .Q(u_muldiv_quotient_q[13]) );
  DFFRX1 u_muldiv_quotient_q_reg_14_ ( .D(u_muldiv_N342), .CK(net1918), .RN(
        n44178), .Q(u_muldiv_quotient_q[14]) );
  DFFRX1 u_muldiv_quotient_q_reg_15_ ( .D(u_muldiv_N343), .CK(net1918), .RN(
        n44178), .Q(u_muldiv_quotient_q[15]) );
  DFFRX1 u_muldiv_quotient_q_reg_16_ ( .D(u_muldiv_N344), .CK(net1923), .RN(
        n44178), .Q(u_muldiv_quotient_q[16]) );
  DFFRX1 u_muldiv_quotient_q_reg_17_ ( .D(u_muldiv_N345), .CK(net1923), .RN(
        n44178), .Q(u_muldiv_quotient_q[17]) );
  DFFRX1 u_muldiv_quotient_q_reg_18_ ( .D(u_muldiv_N346), .CK(net1923), .RN(
        n44178), .Q(u_muldiv_quotient_q[18]) );
  DFFRX1 u_muldiv_quotient_q_reg_19_ ( .D(u_muldiv_N347), .CK(net1923), .RN(
        n44178), .Q(u_muldiv_quotient_q[19]) );
  DFFRX1 u_muldiv_quotient_q_reg_20_ ( .D(u_muldiv_N348), .CK(net1923), .RN(
        n44178), .Q(u_muldiv_quotient_q[20]) );
  DFFRX1 u_muldiv_quotient_q_reg_21_ ( .D(u_muldiv_N349), .CK(net1923), .RN(
        n44178), .Q(u_muldiv_quotient_q[21]) );
  DFFRX1 u_muldiv_quotient_q_reg_22_ ( .D(u_muldiv_N350), .CK(net1923), .RN(
        n44178), .Q(u_muldiv_quotient_q[22]) );
  DFFRX1 u_muldiv_quotient_q_reg_23_ ( .D(u_muldiv_N351), .CK(net1923), .RN(
        n44178), .Q(u_muldiv_quotient_q[23]) );
  DFFRX1 u_muldiv_quotient_q_reg_24_ ( .D(u_muldiv_N352), .CK(net1923), .RN(
        n44178), .Q(u_muldiv_quotient_q[24]) );
  DFFRX1 u_muldiv_quotient_q_reg_25_ ( .D(u_muldiv_N353), .CK(net1923), .RN(
        n44178), .Q(u_muldiv_quotient_q[25]) );
  DFFRX1 u_muldiv_quotient_q_reg_26_ ( .D(u_muldiv_N354), .CK(net1923), .RN(
        n44177), .Q(u_muldiv_quotient_q[26]) );
  DFFRX1 u_muldiv_quotient_q_reg_27_ ( .D(u_muldiv_N355), .CK(net1923), .RN(
        n44177), .Q(u_muldiv_quotient_q[27]) );
  DFFRX1 u_muldiv_quotient_q_reg_28_ ( .D(u_muldiv_N356), .CK(net1923), .RN(
        n44177), .Q(u_muldiv_quotient_q[28]) );
  DFFRX1 u_muldiv_quotient_q_reg_29_ ( .D(u_muldiv_N357), .CK(net1923), .RN(
        n44177), .Q(u_muldiv_quotient_q[29]) );
  DFFRX1 u_muldiv_quotient_q_reg_30_ ( .D(u_muldiv_N358), .CK(net1923), .RN(
        n44177), .Q(u_muldiv_quotient_q[30]) );
  DFFRX1 u_muldiv_quotient_q_reg_31_ ( .D(u_muldiv_N359), .CK(net1923), .RN(
        n44177), .Q(u_muldiv_quotient_q[31]) );
  DFFRX1 u_muldiv_wb_rd_q_reg_0_ ( .D(u_muldiv_N513), .CK(clk_i), .RN(n44177), 
        .Q(writeback_muldiv_idx_w[0]), .QN(n37338) );
  DFFRX1 u_decode_scoreboard_q_reg_16_ ( .D(u_decode_scoreboard_r[16]), .CK(
        clk_i), .RN(n44177), .Q(u_decode_scoreboard_q[16]) );
  DFFRX1 u_muldiv_mult_busy_q_reg ( .D(n36344), .CK(clk_i), .RN(n44209), .Q(
        u_muldiv_mult_busy_q) );
  DFFRX1 u_csr_csr_satp_q_reg_31_ ( .D(u_csr_csr_satp_r[31]), .CK(clk_i), .RN(
        n44209), .Q(u_csr_csr_satp_q_31_), .QN(n42543) );
  DFFRX1 u_mmu_dtlb_entry_q_reg_25_ ( .D(u_mmu_pte_entry_q[25]), .CK(n37872), 
        .RN(n44177), .QN(n1838) );
  DFFRX1 u_mmu_dtlb_entry_q_reg_26_ ( .D(u_mmu_pte_entry_q[26]), .CK(n37872), 
        .RN(n44177), .QN(n1839) );
  DFFRX1 u_mmu_dtlb_entry_q_reg_27_ ( .D(u_mmu_pte_entry_q[27]), .CK(n37872), 
        .RN(n44177), .QN(n1840) );
  DFFRX1 u_mmu_dtlb_entry_q_reg_28_ ( .D(u_mmu_pte_entry_q[28]), .CK(n37872), 
        .RN(n44177), .QN(n1841) );
  DFFRX1 u_mmu_dtlb_entry_q_reg_29_ ( .D(u_mmu_pte_entry_q[29]), .CK(n37872), 
        .RN(n44177), .QN(n1842) );
  DFFRX1 u_mmu_dtlb_entry_q_reg_30_ ( .D(u_mmu_pte_entry_q[30]), .CK(n37872), 
        .RN(n44177), .QN(n1843) );
  DFFRX1 u_mmu_dtlb_entry_q_reg_31_ ( .D(u_mmu_pte_entry_q[31]), .CK(n37872), 
        .RN(n44177), .QN(n1844) );
  DFFRX1 u_mmu_dtlb_entry_q_reg_1_ ( .D(u_mmu_pte_entry_q_1), .CK(net1782), 
        .RN(n44177), .QN(n37433) );
  DFFRX1 u_mmu_dtlb_entry_q_reg_2_ ( .D(u_mmu_pte_entry_q_2), .CK(net1782), 
        .RN(n44177), .Q(n8417) );
  DFFRX1 u_mmu_dtlb_entry_q_reg_4_ ( .D(u_mmu_pte_entry_q_4), .CK(net1782), 
        .RN(n44177), .Q(u_mmu_dtlb_entry_q_4) );
  DFFRX1 u_mmu_dtlb_entry_q_reg_22_ ( .D(u_mmu_pte_entry_q[22]), .CK(net1782), 
        .RN(n44176), .QN(n1845) );
  DFFRX1 u_mmu_dtlb_entry_q_reg_23_ ( .D(u_mmu_pte_entry_q[23]), .CK(net1782), 
        .RN(n44176), .QN(n1846) );
  DFFRX1 u_mmu_dtlb_entry_q_reg_24_ ( .D(u_mmu_pte_entry_q[24]), .CK(net1782), 
        .RN(n44176), .QN(n1847) );
  DFFRX1 u_mmu_itlb_va_addr_q_reg_27_ ( .D(n8442), .CK(clk_i), .RN(n44183), 
        .Q(u_mmu_itlb_va_addr_q[27]) );
  DFFRX1 u_mmu_itlb_entry_q_reg_26_ ( .D(u_mmu_pte_entry_q[26]), .CK(n37871), 
        .RN(n44176), .Q(u_mmu_itlb_entry_q[26]) );
  DFFRX1 u_mmu_itlb_entry_q_reg_27_ ( .D(u_mmu_pte_entry_q[27]), .CK(n37871), 
        .RN(n44176), .Q(u_mmu_itlb_entry_q[27]) );
  DFFRX1 u_mmu_itlb_entry_q_reg_28_ ( .D(u_mmu_pte_entry_q[28]), .CK(n37871), 
        .RN(n44176), .Q(u_mmu_itlb_entry_q[28]) );
  DFFRX1 u_mmu_itlb_entry_q_reg_29_ ( .D(u_mmu_pte_entry_q[29]), .CK(n37871), 
        .RN(n44176), .Q(u_mmu_itlb_entry_q[29]) );
  DFFRX1 u_mmu_itlb_entry_q_reg_30_ ( .D(u_mmu_pte_entry_q[30]), .CK(n37871), 
        .RN(n44176), .Q(u_mmu_itlb_entry_q[30]) );
  DFFRX1 u_mmu_itlb_entry_q_reg_31_ ( .D(u_mmu_pte_entry_q[31]), .CK(n37871), 
        .RN(n44176), .Q(u_mmu_itlb_entry_q[31]) );
  DFFRX1 u_mmu_itlb_entry_q_reg_3_ ( .D(u_mmu_pte_entry_q_3), .CK(net1792), 
        .RN(n44176), .Q(u_mmu_itlb_entry_q_3) );
  DFFRX1 u_mmu_itlb_entry_q_reg_4_ ( .D(u_mmu_pte_entry_q_4), .CK(net1792), 
        .RN(n44176), .Q(u_mmu_itlb_entry_q_4) );
  DFFRX1 u_mmu_itlb_entry_q_reg_22_ ( .D(u_mmu_pte_entry_q[22]), .CK(net1792), 
        .RN(n44176), .Q(u_mmu_itlb_entry_q[22]) );
  DFFRX1 u_mmu_itlb_entry_q_reg_23_ ( .D(u_mmu_pte_entry_q[23]), .CK(net1792), 
        .RN(n44176), .Q(u_mmu_itlb_entry_q[23]) );
  DFFRX1 u_mmu_itlb_entry_q_reg_24_ ( .D(u_mmu_pte_entry_q[24]), .CK(net1792), 
        .RN(n44176), .Q(u_mmu_itlb_entry_q[24]) );
  DFFRX1 u_mmu_itlb_entry_q_reg_25_ ( .D(u_mmu_pte_entry_q[25]), .CK(net1792), 
        .RN(n44176), .Q(u_mmu_itlb_entry_q[25]) );
  DFFRX1 u_decode_inst_q_reg_19_ ( .D(u_decode_N341), .CK(n37870), .RN(n44251), 
        .Q(opcode_opcode_w[19]), .QN(n42791) );
  DFFRX1 u_decode_inst_q_reg_17_ ( .D(u_decode_N339), .CK(n37870), .RN(n44150), 
        .Q(opcode_opcode_w[17]), .QN(n42809) );
  DFFRX1 u_decode_inst_q_reg_16_ ( .D(u_decode_N338), .CK(n37870), .RN(n44201), 
        .Q(opcode_opcode_w[16]), .QN(n42721) );
  DFFRX1 u_muldiv_rd_q_reg_4_ ( .D(n8506), .CK(clk_i), .RN(n44176), .Q(
        u_muldiv_rd_q[4]), .QN(n37781) );
  DFFRX1 u_muldiv_wb_rd_q_reg_4_ ( .D(u_muldiv_N517), .CK(clk_i), .RN(n44176), 
        .Q(writeback_muldiv_idx_w[4]), .QN(n37339) );
  DFFRX1 u_muldiv_rd_q_reg_3_ ( .D(n8507), .CK(clk_i), .RN(n44176), .Q(
        u_muldiv_rd_q[3]), .QN(n37780) );
  DFFRX1 u_muldiv_wb_rd_q_reg_3_ ( .D(u_muldiv_N516), .CK(clk_i), .RN(n44175), 
        .Q(writeback_muldiv_idx_w[3]), .QN(n37542) );
  DFFRX1 u_muldiv_rd_q_reg_2_ ( .D(n8508), .CK(clk_i), .RN(n44175), .Q(
        u_muldiv_rd_q[2]), .QN(n37779) );
  DFFRX1 u_muldiv_wb_rd_q_reg_2_ ( .D(u_muldiv_N515), .CK(clk_i), .RN(n44175), 
        .Q(writeback_muldiv_idx_w[2]) );
  DFFRX1 u_muldiv_rd_q_reg_1_ ( .D(n8509), .CK(clk_i), .RN(n44175), .Q(
        u_muldiv_rd_q[1]), .QN(n37778) );
  DFFRX1 u_muldiv_wb_rd_q_reg_1_ ( .D(u_muldiv_N514), .CK(clk_i), .RN(n44175), 
        .Q(writeback_muldiv_idx_w[1]), .QN(n37541) );
  DFFRX1 u_muldiv_rd_q_reg_0_ ( .D(n8510), .CK(clk_i), .RN(n44175), .Q(
        u_muldiv_rd_q[0]), .QN(n37777) );
  DFFRX1 u_lsu_mem_rd_q_reg ( .D(u_lsu_N103), .CK(n37869), .RN(n44250), .Q(
        n42558), .QN(n8574) );
  DFFRX1 u_mmu_load_q_reg ( .D(n8441), .CK(clk_i), .RN(n44123), .Q(
        u_mmu_load_q), .QN(n37425) );
  DFFRX1 u_lsu_mem_invalidate_q_reg ( .D(u_lsu_N230), .CK(n37869), .RN(n44175), 
        .QN(n8647) );
  DFFRX1 u_lsu_mem_addr_q_reg_0_ ( .D(n73431), .CK(n37869), .RN(n44210), .Q(
        mmu_lsu_addr_w[0]), .QN(n1857) );
  DFFRX1 u_mmu_lsu_in_addr_q_reg_0_ ( .D(mmu_lsu_addr_w[0]), .CK(n37875), .RN(
        n44210), .Q(n57894), .QN(n1858) );
  DFFRX1 u_lsu_mem_addr_q_reg_1_ ( .D(n73430), .CK(n37869), .RN(n44197), .Q(
        mmu_lsu_addr_w[1]), .QN(n1859) );
  DFFRX1 u_mmu_lsu_in_addr_q_reg_1_ ( .D(mmu_lsu_addr_w[1]), .CK(n37875), .RN(
        n44197), .Q(n57992), .QN(n1860) );
  DFFRX1 u_lsu_mem_addr_q_reg_2_ ( .D(u_lsu_mem_addr_r[2]), .CK(n37869), .RN(
        n44198), .Q(mmu_lsu_addr_w[2]), .QN(n1861) );
  DFFRX1 u_mmu_lsu_in_addr_q_reg_2_ ( .D(mmu_lsu_addr_w[2]), .CK(n37875), .RN(
        n44198), .QN(n1862) );
  DFFRX1 u_lsu_mem_addr_q_reg_3_ ( .D(u_lsu_mem_addr_r[3]), .CK(n37869), .RN(
        n44198), .Q(mmu_lsu_addr_w[3]), .QN(n1863) );
  DFFRX1 u_mmu_lsu_in_addr_q_reg_3_ ( .D(mmu_lsu_addr_w[3]), .CK(n37875), .RN(
        n44198), .QN(n1864) );
  DFFRX1 u_lsu_mem_addr_q_reg_4_ ( .D(u_lsu_mem_addr_r[4]), .CK(n37869), .RN(
        n44199), .Q(mmu_lsu_addr_w[4]), .QN(n1865) );
  DFFRX1 u_mmu_lsu_in_addr_q_reg_4_ ( .D(mmu_lsu_addr_w[4]), .CK(n37875), .RN(
        n44199), .QN(n1866) );
  DFFRX1 u_lsu_mem_addr_q_reg_5_ ( .D(u_lsu_mem_addr_r[5]), .CK(n37869), .RN(
        n44199), .Q(mmu_lsu_addr_w[5]), .QN(n1867) );
  DFFRX1 u_mmu_lsu_in_addr_q_reg_5_ ( .D(mmu_lsu_addr_w[5]), .CK(n37875), .RN(
        n44199), .QN(n1868) );
  DFFRX1 u_lsu_mem_addr_q_reg_15_ ( .D(u_lsu_mem_addr_r[15]), .CK(n37876), 
        .RN(n44185), .Q(mmu_lsu_addr_w[15]), .QN(n8302) );
  DFFRX1 u_mmu_lsu_in_addr_q_reg_15_ ( .D(mmu_lsu_addr_w[15]), .CK(n37875), 
        .RN(n44185), .QN(n1869) );
  DFFRX1 u_lsu_mem_addr_q_reg_28_ ( .D(u_lsu_mem_addr_r[28]), .CK(n37876), 
        .RN(n44185), .Q(n56708), .QN(n8330) );
  DFFRX1 u_mmu_lsu_in_addr_q_reg_28_ ( .D(n56708), .CK(n37873), .RN(n44206), 
        .QN(n1870) );
  DFFRX1 u_lsu_mem_addr_q_reg_30_ ( .D(u_lsu_mem_addr_r[30]), .CK(n37874), 
        .RN(n44182), .Q(n56553), .QN(n8336) );
  DFFRX1 u_mmu_lsu_in_addr_q_reg_30_ ( .D(n56553), .CK(n37873), .RN(n44206), 
        .QN(n1871) );
  DFFRX1 u_lsu_mem_addr_q_reg_31_ ( .D(u_lsu_mem_addr_r[31]), .CK(n37874), 
        .RN(n44183), .Q(n56627), .QN(n8338) );
  DFFRX1 u_mmu_lsu_in_addr_q_reg_31_ ( .D(n56627), .CK(n37873), .RN(n44206), 
        .QN(n1872) );
  DFFRX1 u_lsu_mem_wr_q_reg_0_ ( .D(u_lsu_N226), .CK(n37868), .RN(n44205), .Q(
        n58194) );
  DFFRX1 u_lsu_mem_wr_q_reg_1_ ( .D(u_lsu_N227), .CK(n37868), .RN(n44205), .Q(
        n37328) );
  DFFRX1 u_lsu_mem_wr_q_reg_2_ ( .D(u_lsu_N228), .CK(n37868), .RN(n44205), .Q(
        n37327) );
  DFFRX1 u_lsu_mem_wr_q_reg_3_ ( .D(u_lsu_N229), .CK(n37868), .RN(n44205), .Q(
        n58184) );
  DFFRX1 u_mmu_store_q_reg_2_ ( .D(n8540), .CK(clk_i), .RN(n44205), .Q(
        u_mmu_store_q[2]), .QN(n37329) );
  DFFRX1 u_mmu_store_q_reg_1_ ( .D(n8541), .CK(clk_i), .RN(n44205), .Q(
        u_mmu_store_q[1]), .QN(n37431) );
  DFFRX1 u_mmu_store_q_reg_0_ ( .D(n8542), .CK(clk_i), .RN(n44205), .Q(
        u_mmu_store_q[0]), .QN(n42610) );
  DFFRX1 u_lsu_mem_unaligned_ld_q_reg ( .D(u_lsu_N98), .CK(n37868), .RN(n44209), .Q(n37353), .QN(n8810) );
  DFFRX1 u_lsu_mem_flush_q_reg ( .D(u_lsu_N231), .CK(n37868), .RN(n44175), 
        .QN(n8954) );
  DFFRX1 u_lsu_mem_req_tag_q_reg_0_ ( .D(opcode_opcode_w[7]), .CK(n37868), 
        .RN(n44171), .QN(n1877) );
  DFFRX1 u_lsu_mem_req_tag_q_reg_1_ ( .D(opcode_opcode_w[8]), .CK(n37868), 
        .RN(n44200), .QN(n1878) );
  DFFRX1 u_lsu_mem_req_tag_q_reg_2_ ( .D(opcode_opcode_w[9]), .CK(n37868), 
        .RN(n44200), .QN(n1879) );
  DFFRX1 u_lsu_mem_req_tag_q_reg_3_ ( .D(opcode_opcode_w[10]), .CK(n37868), 
        .RN(n44179), .QN(n1880) );
  DFFRX1 u_lsu_mem_req_tag_q_reg_4_ ( .D(opcode_opcode_w[11]), .CK(n37868), 
        .RN(n44087), .QN(n1881) );
  DFFRX1 u_lsu_mem_req_tag_q_reg_5_ ( .D(n73431), .CK(n37868), .RN(n44200), 
        .QN(n1882) );
  DFFRX1 u_lsu_mem_req_tag_q_reg_6_ ( .D(n8498), .CK(clk_i), .RN(n44175), .QN(
        n1883) );
  DFFRX1 u_lsu_mem_req_tag_q_reg_8_ ( .D(n8496), .CK(clk_i), .RN(n44175), .QN(
        n1884) );
  DFFRX1 u_lsu_mem_req_tag_q_reg_9_ ( .D(n8495), .CK(clk_i), .RN(n44175), .QN(
        n1885) );
  DFFRX1 u_lsu_mem_req_tag_q_reg_10_ ( .D(n8494), .CK(clk_i), .RN(n44175), 
        .QN(n1886) );
  DFFRX1 u_lsu_mem_unaligned_st_q_reg ( .D(u_lsu_N99), .CK(n37868), .RN(n44209), .QN(n1887) );
  DFFRX1 u_lsu_mem_req_tag_q_reg_7_ ( .D(n4705), .CK(n37869), .RN(n44175), 
        .QN(n8255) );
  DFFRX1 u_csr_csr_satp_q_reg_8_ ( .D(u_csr_csr_satp_r[8]), .CK(clk_i), .RN(
        n44197), .Q(n73414) );
  DFFRX1 u_csr_csr_mtvec_q_reg_8_ ( .D(u_csr_csr_mtvec_r[8]), .CK(clk_i), .RN(
        n44175), .Q(u_csr_csr_mtvec_q[8]), .QN(n37710) );
  DFFRX1 u_csr_csr_satp_q_reg_7_ ( .D(u_csr_csr_satp_r[7]), .CK(clk_i), .RN(
        n44196), .Q(n73415) );
  DFFRX1 u_csr_csr_mtvec_q_reg_7_ ( .D(u_csr_csr_mtvec_r[7]), .CK(clk_i), .RN(
        n44175), .Q(u_csr_csr_mtvec_q[7]), .QN(n37715) );
  DFFRX1 u_csr_csr_satp_q_reg_5_ ( .D(u_csr_csr_satp_r[5]), .CK(clk_i), .RN(
        n44196), .Q(n73416) );
  DFFRX1 u_csr_csr_mtvec_q_reg_5_ ( .D(u_csr_csr_mtvec_r[5]), .CK(clk_i), .RN(
        n44174), .Q(u_csr_csr_mtvec_q[5]), .QN(n37714) );
  DFFRX1 u_csr_csr_satp_q_reg_3_ ( .D(u_csr_csr_satp_r[3]), .CK(clk_i), .RN(
        n44211), .Q(n57946), .QN(n1895) );
  DFFRX1 u_csr_csr_mtvec_q_reg_3_ ( .D(u_csr_csr_mtvec_r[3]), .CK(clk_i), .RN(
        n44174), .Q(u_csr_csr_mtvec_q[3]), .QN(n37700) );
  DFFRX1 u_csr_csr_mscratch_q_reg_3_ ( .D(u_csr_csr_mscratch_r[3]), .CK(clk_i), 
        .RN(n44174), .Q(u_csr_csr_mscratch_q[3]) );
  DFFRX1 u_csr_csr_mtvec_q_reg_31_ ( .D(u_csr_csr_mtvec_r[31]), .CK(clk_i), 
        .RN(n44174), .Q(u_csr_csr_mtvec_q[31]), .QN(n37745) );
  DFFRX1 u_csr_csr_mtvec_q_reg_30_ ( .D(u_csr_csr_mtvec_r[30]), .CK(clk_i), 
        .RN(n44174), .Q(u_csr_csr_mtvec_q[30]), .QN(n37744) );
  DFFRX1 u_csr_csr_mtvec_q_reg_29_ ( .D(u_csr_csr_mtvec_r[29]), .CK(clk_i), 
        .RN(n44174), .Q(u_csr_csr_mtvec_q[29]), .QN(n37743) );
  DFFRX1 u_csr_csr_mtvec_q_reg_28_ ( .D(u_csr_csr_mtvec_r[28]), .CK(clk_i), 
        .RN(n44174), .Q(u_csr_csr_mtvec_q[28]), .QN(n37742) );
  DFFRX1 u_csr_csr_mtvec_q_reg_27_ ( .D(u_csr_csr_mtvec_r[27]), .CK(clk_i), 
        .RN(n44174), .Q(u_csr_csr_mtvec_q[27]), .QN(n37741) );
  DFFRX1 u_csr_csr_mtvec_q_reg_26_ ( .D(u_csr_csr_mtvec_r[26]), .CK(clk_i), 
        .RN(n44174), .Q(u_csr_csr_mtvec_q[26]), .QN(n37740) );
  DFFRX1 u_csr_csr_mtvec_q_reg_25_ ( .D(u_csr_csr_mtvec_r[25]), .CK(clk_i), 
        .RN(n44174), .Q(u_csr_csr_mtvec_q[25]), .QN(n37739) );
  DFFRX1 u_csr_csr_mtvec_q_reg_24_ ( .D(u_csr_csr_mtvec_r[24]), .CK(clk_i), 
        .RN(n44173), .Q(u_csr_csr_mtvec_q[24]), .QN(n37738) );
  DFFRX1 u_csr_csr_mtvec_q_reg_23_ ( .D(u_csr_csr_mtvec_r[23]), .CK(clk_i), 
        .RN(n44173), .Q(u_csr_csr_mtvec_q[23]), .QN(n37737) );
  DFFRX1 u_csr_csr_mtvec_q_reg_1_ ( .D(u_csr_csr_mtvec_r[1]), .CK(clk_i), .RN(
        n44173), .Q(u_csr_csr_mtvec_q[1]), .QN(n37713) );
  DFFRX1 u_csr_csr_mscratch_q_reg_1_ ( .D(u_csr_csr_mscratch_r[1]), .CK(clk_i), 
        .RN(n44173), .Q(u_csr_csr_mscratch_q[1]) );
  DFFRX1 u_csr_csr_mtvec_q_reg_11_ ( .D(u_csr_csr_mtvec_r[11]), .CK(clk_i), 
        .RN(n44173), .Q(u_csr_csr_mtvec_q[11]), .QN(n37708) );
  DFFRX1 u_csr_csr_mtvec_q_reg_12_ ( .D(u_csr_csr_mtvec_r[12]), .CK(clk_i), 
        .RN(n44173), .Q(u_csr_csr_mtvec_q[12]), .QN(n37720) );
  DFFRX1 u_csr_csr_mtvec_q_reg_22_ ( .D(u_csr_csr_mtvec_r[22]), .CK(clk_i), 
        .RN(n44173), .Q(u_csr_csr_mtvec_q[22]), .QN(n37736) );
  DFFRX1 u_csr_csr_mtvec_q_reg_21_ ( .D(u_csr_csr_mtvec_r[21]), .CK(clk_i), 
        .RN(n44173), .Q(u_csr_csr_mtvec_q[21]), .QN(n37735) );
  DFFRX1 u_csr_csr_mtvec_q_reg_20_ ( .D(u_csr_csr_mtvec_r[20]), .CK(clk_i), 
        .RN(n44173), .Q(u_csr_csr_mtvec_q[20]), .QN(n37734) );
  DFFRX1 u_csr_csr_mtvec_q_reg_19_ ( .D(u_csr_csr_mtvec_r[19]), .CK(clk_i), 
        .RN(n44173), .Q(u_csr_csr_mtvec_q[19]), .QN(n37733) );
  DFFRX1 u_csr_csr_mtvec_q_reg_18_ ( .D(u_csr_csr_mtvec_r[18]), .CK(clk_i), 
        .RN(n44172), .Q(u_csr_csr_mtvec_q[18]), .QN(n37732) );
  DFFRX1 u_csr_csr_sr_q_reg_18_ ( .D(u_csr_N2391), .CK(net1878), .RN(n44172), 
        .Q(n37776), .QN(n8835) );
  DFFRX1 u_csr_pc_m_q_reg_30_ ( .D(n8499), .CK(clk_i), .RN(n44182), .Q(
        u_csr_pc_m_q[30]), .QN(n37760) );
  DFFRX1 u_csr_pc_m_q_reg_31_ ( .D(n8537), .CK(clk_i), .RN(n44182), .Q(
        u_csr_pc_m_q[31]), .QN(n37761) );
  DFFRX1 u_csr_writeback_idx_q_reg_0_ ( .D(opcode_opcode_w[7]), .CK(net1867), 
        .RN(n44200), .Q(u_csr_writeback_idx_q[0]), .QN(n37537) );
  DFFRX1 u_csr_writeback_idx_q_reg_1_ ( .D(opcode_opcode_w[8]), .CK(net1867), 
        .RN(n44200), .Q(u_csr_writeback_idx_q[1]), .QN(n37336) );
  DFFRX1 u_csr_writeback_idx_q_reg_2_ ( .D(opcode_opcode_w[9]), .CK(net1867), 
        .RN(n44200), .Q(u_csr_writeback_idx_q[2]), .QN(n37483) );
  DFFRX1 u_csr_writeback_idx_q_reg_3_ ( .D(opcode_opcode_w[10]), .CK(net1867), 
        .RN(n44207), .Q(u_csr_writeback_idx_q[3]), .QN(n37351) );
  DFFRX1 u_csr_writeback_idx_q_reg_4_ ( .D(opcode_opcode_w[11]), .CK(net1867), 
        .RN(n44207), .Q(u_csr_writeback_idx_q[4]), .QN(n37592) );
  DFFRX1 u_csr_pc_m_q_reg_15_ ( .D(opcode_pc_w[15]), .CK(net1872), .RN(n44107), 
        .Q(n1896) );
  DFFRX1 u_csr_writeback_en_q_reg ( .D(u_csr_N3471), .CK(clk_i), .RN(n44208), 
        .Q(u_csr_writeback_en_q), .QN(n37589) );
  DFFRX1 u_csr_csr_mtvec_q_reg_17_ ( .D(u_csr_csr_mtvec_r[17]), .CK(clk_i), 
        .RN(n44172), .Q(u_csr_csr_mtvec_q[17]), .QN(n37731) );
  DFFRX1 u_csr_csr_mtvec_q_reg_16_ ( .D(u_csr_csr_mtvec_r[16]), .CK(clk_i), 
        .RN(n44172), .Q(u_csr_csr_mtvec_q[16]), .QN(n37730) );
  DFFRX1 u_csr_csr_mtvec_q_reg_15_ ( .D(u_csr_csr_mtvec_r[15]), .CK(clk_i), 
        .RN(n44172), .Q(u_csr_csr_mtvec_q[15]), .QN(n37719) );
  DFFRX1 u_csr_csr_mtvec_q_reg_14_ ( .D(u_csr_csr_mtvec_r[14]), .CK(clk_i), 
        .RN(n44172), .Q(u_csr_csr_mtvec_q[14]), .QN(n37718) );
  DFFRX1 u_csr_csr_mtvec_q_reg_13_ ( .D(u_csr_csr_mtvec_r[13]), .CK(clk_i), 
        .RN(n44172), .Q(u_csr_csr_mtvec_q[13]), .QN(n37717) );
  DFFRX1 u_csr_csr_mtvec_q_reg_10_ ( .D(u_csr_csr_mtvec_r[10]), .CK(clk_i), 
        .RN(n44172), .Q(u_csr_csr_mtvec_q[10]), .QN(n37704) );
  DFFRX1 u_csr_csr_mscratch_q_reg_10_ ( .D(u_csr_csr_mscratch_r[10]), .CK(
        clk_i), .RN(n44172), .Q(u_csr_csr_mscratch_q[10]) );
  DFFRX1 u_csr_csr_satp_q_reg_9_ ( .D(u_csr_csr_satp_r[9]), .CK(clk_i), .RN(
        n44197), .Q(n73413) );
  DFFRX1 u_csr_csr_mtvec_q_reg_9_ ( .D(u_csr_csr_mtvec_r[9]), .CK(clk_i), .RN(
        n44172), .Q(u_csr_csr_mtvec_q[9]), .QN(n37716) );
  DFFRX1 u_csr_csr_mscratch_q_reg_9_ ( .D(u_csr_csr_mscratch_r[9]), .CK(clk_i), 
        .RN(n44172), .Q(u_csr_csr_mscratch_q[9]) );
  DFFRX1 u_csr_csr_satp_q_reg_6_ ( .D(u_csr_csr_satp_r[6]), .CK(clk_i), .RN(
        n44196), .Q(n57977), .QN(n1898) );
  DFFRX1 u_csr_csr_mtvec_q_reg_6_ ( .D(u_csr_csr_mtvec_r[6]), .CK(clk_i), .RN(
        n44171), .Q(u_csr_csr_mtvec_q[6]), .QN(n37706) );
  DFFRX1 u_csr_csr_mscratch_q_reg_6_ ( .D(u_csr_csr_mscratch_r[6]), .CK(clk_i), 
        .RN(n44171), .Q(u_csr_csr_mscratch_q[6]) );
  DFFRX1 u_csr_csr_satp_q_reg_4_ ( .D(u_csr_csr_satp_r[4]), .CK(clk_i), .RN(
        n44211), .Q(n57957), .QN(n1899) );
  DFFRX1 u_csr_csr_mtvec_q_reg_4_ ( .D(u_csr_csr_mtvec_r[4]), .CK(clk_i), .RN(
        n44171), .Q(u_csr_csr_mtvec_q[4]), .QN(n37705) );
  DFFRX1 u_csr_csr_mscratch_q_reg_4_ ( .D(u_csr_csr_mscratch_r[4]), .CK(clk_i), 
        .RN(n44175), .Q(u_csr_csr_mscratch_q[4]) );
  DFFRX1 u_csr_csr_sr_q_reg_4_ ( .D(u_csr_N2377), .CK(net1878), .RN(n44155), 
        .Q(u_csr_csr_sr_q[4]) );
  DFFRX1 u_csr_csr_mtvec_q_reg_2_ ( .D(u_csr_csr_mtvec_r[2]), .CK(clk_i), .RN(
        n44155), .Q(u_csr_csr_mtvec_q[2]), .QN(n37709) );
  DFFRX1 u_csr_csr_mscratch_q_reg_2_ ( .D(u_csr_csr_mscratch_r[2]), .CK(clk_i), 
        .RN(n44155), .Q(u_csr_csr_mscratch_q[2]) );
  DFFRX1 u_csr_csr_mip_q_reg_7_ ( .D(u_csr_csr_mip_r_7), .CK(clk_i), .RN(
        n44155), .Q(u_csr_csr_mip_q_7), .QN(n37545) );
  DFFRX1 u_csr_csr_mie_q_reg_1_ ( .D(u_csr_csr_mie_r_1), .CK(clk_i), .RN(
        n44155), .Q(u_csr_csr_mie_q_1) );
  DFFRX1 u_csr_csr_mie_q_reg_3_ ( .D(u_csr_csr_mie_r_3), .CK(clk_i), .RN(
        n44155), .Q(u_csr_csr_mie_q_3), .QN(n37544) );
  DFFRX1 u_csr_csr_medeleg_q_reg_0_ ( .D(u_csr_csr_medeleg_r[0]), .CK(clk_i), 
        .RN(n44155), .Q(u_csr_csr_medeleg_q[0]) );
  DFFRX1 u_csr_csr_medeleg_q_reg_10_ ( .D(u_csr_csr_medeleg_r[10]), .CK(clk_i), 
        .RN(n44155), .Q(u_csr_csr_medeleg_q[10]) );
  DFFRX1 u_csr_csr_medeleg_q_reg_11_ ( .D(u_csr_csr_medeleg_r[11]), .CK(clk_i), 
        .RN(n44155), .Q(u_csr_csr_medeleg_q[11]) );
  DFFRX1 u_csr_csr_medeleg_q_reg_12_ ( .D(u_csr_csr_medeleg_r[12]), .CK(clk_i), 
        .RN(n44155), .Q(u_csr_csr_medeleg_q[12]) );
  DFFRX1 u_csr_csr_medeleg_q_reg_13_ ( .D(u_csr_csr_medeleg_r[13]), .CK(clk_i), 
        .RN(n44123), .Q(u_csr_csr_medeleg_q[13]) );
  DFFRX1 u_csr_csr_medeleg_q_reg_14_ ( .D(u_csr_csr_medeleg_r[14]), .CK(clk_i), 
        .RN(n44154), .Q(u_csr_csr_medeleg_q[14]) );
  DFFRX1 u_csr_csr_medeleg_q_reg_15_ ( .D(u_csr_csr_medeleg_r[15]), .CK(clk_i), 
        .RN(n44125), .Q(u_csr_csr_medeleg_q[15]) );
  DFFRX1 u_csr_csr_medeleg_q_reg_1_ ( .D(u_csr_csr_medeleg_r[1]), .CK(clk_i), 
        .RN(n44154), .Q(u_csr_csr_medeleg_q[1]) );
  DFFRX1 u_csr_csr_medeleg_q_reg_2_ ( .D(u_csr_csr_medeleg_r[2]), .CK(clk_i), 
        .RN(n44154), .Q(u_csr_csr_medeleg_q[2]) );
  DFFRX1 u_csr_csr_medeleg_q_reg_3_ ( .D(u_csr_csr_medeleg_r[3]), .CK(clk_i), 
        .RN(n44154), .Q(u_csr_csr_medeleg_q[3]) );
  DFFRX1 u_csr_csr_medeleg_q_reg_4_ ( .D(u_csr_csr_medeleg_r[4]), .CK(clk_i), 
        .RN(n44154), .Q(u_csr_csr_medeleg_q[4]), .QN(n40932) );
  DFFRX1 u_csr_csr_medeleg_q_reg_5_ ( .D(u_csr_csr_medeleg_r[5]), .CK(clk_i), 
        .RN(n44154), .Q(u_csr_csr_medeleg_q[5]) );
  DFFRX1 u_csr_csr_medeleg_q_reg_6_ ( .D(u_csr_csr_medeleg_r[6]), .CK(clk_i), 
        .RN(n44154), .Q(u_csr_csr_medeleg_q[6]), .QN(n40933) );
  DFFRX1 u_csr_csr_medeleg_q_reg_7_ ( .D(u_csr_csr_medeleg_r[7]), .CK(clk_i), 
        .RN(n44154), .Q(u_csr_csr_medeleg_q[7]), .QN(n37566) );
  DFFRX1 u_csr_csr_medeleg_q_reg_8_ ( .D(u_csr_csr_medeleg_r[8]), .CK(clk_i), 
        .RN(n44154), .Q(u_csr_csr_medeleg_q[8]) );
  DFFRX1 u_csr_csr_medeleg_q_reg_9_ ( .D(u_csr_csr_medeleg_r[9]), .CK(clk_i), 
        .RN(n44154), .Q(u_csr_csr_medeleg_q[9]) );
  DFFRX1 u_csr_csr_mideleg_q_reg_0_ ( .D(u_csr_csr_mideleg_r[0]), .CK(clk_i), 
        .RN(n44154), .Q(u_csr_csr_mideleg_q[0]) );
  DFFRX1 u_csr_csr_mideleg_q_reg_10_ ( .D(u_csr_csr_mideleg_r[10]), .CK(clk_i), 
        .RN(n44154), .Q(u_csr_csr_mideleg_q[10]) );
  DFFRX1 u_csr_csr_mideleg_q_reg_11_ ( .D(u_csr_csr_mideleg_r[11]), .CK(clk_i), 
        .RN(n44154), .Q(u_csr_csr_mideleg_q[11]) );
  DFFRX1 u_csr_csr_mideleg_q_reg_12_ ( .D(u_csr_csr_mideleg_r[12]), .CK(clk_i), 
        .RN(n44154), .Q(u_csr_csr_mideleg_q[12]) );
  DFFRX1 u_csr_csr_mideleg_q_reg_13_ ( .D(u_csr_csr_mideleg_r[13]), .CK(clk_i), 
        .RN(n44154), .Q(u_csr_csr_mideleg_q[13]) );
  DFFRX1 u_csr_csr_mideleg_q_reg_14_ ( .D(u_csr_csr_mideleg_r[14]), .CK(clk_i), 
        .RN(n44154), .Q(u_csr_csr_mideleg_q[14]) );
  DFFRX1 u_csr_csr_mideleg_q_reg_15_ ( .D(u_csr_csr_mideleg_r[15]), .CK(clk_i), 
        .RN(n44154), .Q(u_csr_csr_mideleg_q[15]) );
  DFFRX1 u_csr_csr_mideleg_q_reg_1_ ( .D(u_csr_csr_mideleg_r[1]), .CK(clk_i), 
        .RN(n44154), .Q(u_csr_csr_mideleg_q[1]), .QN(n40923) );
  DFFRX1 u_csr_csr_mideleg_q_reg_2_ ( .D(u_csr_csr_mideleg_r[2]), .CK(clk_i), 
        .RN(n44153), .Q(u_csr_csr_mideleg_q[2]) );
  DFFRX1 u_csr_csr_mideleg_q_reg_3_ ( .D(u_csr_csr_mideleg_r[3]), .CK(clk_i), 
        .RN(n44153), .Q(u_csr_csr_mideleg_q[3]), .QN(n37533) );
  DFFRX1 u_csr_csr_mideleg_q_reg_4_ ( .D(u_csr_csr_mideleg_r[4]), .CK(clk_i), 
        .RN(n44153), .Q(u_csr_csr_mideleg_q[4]) );
  DFFRX1 u_csr_csr_mideleg_q_reg_5_ ( .D(u_csr_csr_mideleg_r[5]), .CK(clk_i), 
        .RN(n44153), .Q(u_csr_csr_mideleg_q[5]) );
  DFFRX1 u_csr_csr_mideleg_q_reg_6_ ( .D(u_csr_csr_mideleg_r[6]), .CK(clk_i), 
        .RN(n44153), .Q(u_csr_csr_mideleg_q[6]) );
  DFFRX1 u_csr_csr_mideleg_q_reg_7_ ( .D(u_csr_csr_mideleg_r[7]), .CK(clk_i), 
        .RN(n44153), .Q(u_csr_csr_mideleg_q[7]) );
  DFFRX1 u_csr_csr_mideleg_q_reg_8_ ( .D(u_csr_csr_mideleg_r[8]), .CK(clk_i), 
        .RN(n44153), .Q(u_csr_csr_mideleg_q[8]) );
  DFFRX1 u_csr_csr_mideleg_q_reg_9_ ( .D(u_csr_csr_mideleg_r[9]), .CK(clk_i), 
        .RN(n44153), .Q(u_csr_csr_mideleg_q[9]), .QN(n37531) );
  DFFRX1 u_csr_csr_mie_q_reg_11_ ( .D(\u_csr_csr_mie_r[11] ), .CK(clk_i), .RN(
        n44153), .Q(\u_csr_csr_mie_q[11] ), .QN(n37485) );
  DFFRX1 u_csr_csr_mie_q_reg_5_ ( .D(u_csr_csr_mie_r_5), .CK(clk_i), .RN(
        n44153), .Q(u_csr_csr_mie_q_5), .QN(n37331) );
  DFFRX1 u_csr_csr_mie_q_reg_7_ ( .D(u_csr_csr_mie_r_7), .CK(clk_i), .RN(
        n44153), .Q(u_csr_csr_mie_q_7), .QN(n37330) );
  DFFRX1 u_csr_csr_mie_q_reg_9_ ( .D(u_csr_csr_mie_r_9), .CK(clk_i), .RN(
        n44153), .Q(u_csr_csr_mie_q_9), .QN(n37549) );
  DFFRX1 u_csr_csr_mip_q_reg_11_ ( .D(\u_csr_csr_mip_r[11] ), .CK(clk_i), .RN(
        n44153), .Q(\u_csr_csr_mip_q[11] ), .QN(n37553) );
  DFFRX1 u_csr_csr_mip_q_reg_1_ ( .D(u_csr_csr_mip_r_1), .CK(clk_i), .RN(
        n44153), .Q(u_csr_csr_mip_q_1) );
  DFFRX1 u_csr_csr_mip_q_reg_3_ ( .D(u_csr_csr_mip_r_3), .CK(clk_i), .RN(
        n44153), .Q(u_csr_csr_mip_q_3), .QN(n37335) );
  DFFRX1 u_csr_csr_mip_q_reg_5_ ( .D(u_csr_csr_mip_r_5), .CK(clk_i), .RN(
        n44153), .Q(u_csr_csr_mip_q_5), .QN(n37546) );
  DFFRX1 u_csr_csr_mip_q_reg_9_ ( .D(u_csr_csr_mip_r_9), .CK(clk_i), .RN(
        n44153), .QN(n37334) );
  DFFRX1 u_csr_csr_sr_q_reg_22_ ( .D(u_csr_N2395), .CK(net1878), .RN(n44153), 
        .Q(u_csr_csr_sr_q_22) );
  DFFRX1 u_csr_csr_sr_q_reg_21_ ( .D(u_csr_N2394), .CK(net1878), .RN(n44152), 
        .Q(u_csr_csr_sr_q_21) );
  DFFRX1 u_csr_csr_sr_q_reg_20_ ( .D(u_csr_N2393), .CK(net1878), .RN(n44152), 
        .Q(u_csr_csr_sr_q_20) );
  DFFRX1 u_csr_csr_sr_q_reg_19_ ( .D(u_csr_N2392), .CK(net1878), .RN(n44152), 
        .Q(u_csr_csr_sr_q_19) );
  DFFRX1 u_csr_csr_sr_q_reg_17_ ( .D(u_csr_N2390), .CK(net1878), .RN(n44152), 
        .Q(u_csr_csr_sr_q[17]) );
  DFFRX1 u_csr_csr_sr_q_reg_16_ ( .D(u_csr_N2389), .CK(net1878), .RN(n44152), 
        .Q(u_csr_csr_sr_q[16]) );
  DFFRX1 u_csr_csr_sr_q_reg_15_ ( .D(u_csr_N2388), .CK(net1878), .RN(n44152), 
        .Q(u_csr_csr_sr_q[15]) );
  DFFRX1 u_csr_csr_sr_q_reg_14_ ( .D(u_csr_N2387), .CK(net1878), .RN(n44152), 
        .Q(u_csr_csr_sr_q[14]) );
  DFFRX1 u_csr_csr_sr_q_reg_13_ ( .D(u_csr_N2386), .CK(net1878), .RN(n44152), 
        .Q(u_csr_csr_sr_q[13]) );
  DFFRX1 u_csr_csr_sr_q_reg_10_ ( .D(u_csr_N2383), .CK(net1878), .RN(n44152), 
        .Q(u_csr_csr_sr_q[10]) );
  DFFRX1 u_csr_csr_sr_q_reg_9_ ( .D(u_csr_N2382), .CK(net1878), .RN(n44152), 
        .Q(u_csr_csr_sr_q[9]) );
  DFFRX1 u_csr_csr_sr_q_reg_6_ ( .D(u_csr_N2379), .CK(net1878), .RN(n44152), 
        .Q(u_csr_csr_sr_q[6]) );
  DFFRX1 u_csr_csr_sr_q_reg_2_ ( .D(u_csr_N2375), .CK(net1878), .RN(n44152), 
        .Q(u_csr_csr_sr_q[2]) );
  DFFRX1 u_csr_csr_mtvec_q_reg_0_ ( .D(u_csr_csr_mtvec_r[0]), .CK(clk_i), .RN(
        n44152), .Q(u_csr_csr_mtvec_q[0]), .QN(n37707) );
  DFFRX1 u_csr_csr_mscratch_q_reg_0_ ( .D(u_csr_csr_mscratch_r[0]), .CK(clk_i), 
        .RN(n44152), .Q(u_csr_csr_mscratch_q[0]) );
  DFFRX1 u_csr_csr_sr_q_reg_0_ ( .D(u_csr_N2373), .CK(net1878), .RN(n44152), 
        .Q(u_csr_csr_sr_q[0]) );
  DFFRX1 u_csr_csr_satp_q_reg_30_ ( .D(u_csr_csr_satp_r[30]), .CK(clk_i), .RN(
        n44152), .Q(n73062), .QN(n1902) );
  DFFRX1 u_csr_csr_satp_q_reg_2_ ( .D(u_csr_csr_satp_r[2]), .CK(clk_i), .RN(
        n44211), .Q(n57937), .QN(n1903) );
  DFFRX1 u_csr_csr_satp_q_reg_29_ ( .D(u_csr_csr_satp_r[29]), .CK(clk_i), .RN(
        n44152), .Q(n73559) );
  DFFRX1 u_csr_csr_satp_q_reg_28_ ( .D(u_csr_csr_satp_r[28]), .CK(clk_i), .RN(
        n44152), .Q(n73560) );
  DFFRX1 u_csr_csr_satp_q_reg_27_ ( .D(u_csr_csr_satp_r[27]), .CK(clk_i), .RN(
        n44151), .Q(n73561) );
  DFFRX1 u_csr_csr_satp_q_reg_26_ ( .D(u_csr_csr_satp_r[26]), .CK(clk_i), .RN(
        n44151), .Q(n73562) );
  DFFRX1 u_csr_csr_satp_q_reg_25_ ( .D(u_csr_csr_satp_r[25]), .CK(clk_i), .RN(
        n44151), .Q(n73563) );
  DFFRX1 u_csr_csr_satp_q_reg_24_ ( .D(u_csr_csr_satp_r[24]), .CK(clk_i), .RN(
        n44151), .Q(n73564) );
  DFFRX1 u_csr_csr_satp_q_reg_23_ ( .D(u_csr_csr_satp_r[23]), .CK(clk_i), .RN(
        n44151), .Q(n73565) );
  DFFRX1 u_csr_csr_satp_q_reg_22_ ( .D(u_csr_csr_satp_r[22]), .CK(clk_i), .RN(
        n44151), .Q(n73566) );
  DFFRX1 u_csr_csr_satp_q_reg_21_ ( .D(u_csr_csr_satp_r[21]), .CK(clk_i), .RN(
        n44151), .Q(n73567) );
  DFFRX1 u_csr_csr_satp_q_reg_20_ ( .D(u_csr_csr_satp_r[20]), .CK(clk_i), .RN(
        n44151), .Q(n73031), .QN(n1913) );
  DFFRX1 u_csr_csr_satp_q_reg_1_ ( .D(u_csr_csr_satp_r[1]), .CK(clk_i), .RN(
        n44210), .Q(n73417) );
  DFFRX1 u_csr_csr_satp_q_reg_19_ ( .D(u_csr_csr_satp_r[19]), .CK(clk_i), .RN(
        n44198), .Q(n73408) );
  DFFRX1 u_csr_csr_satp_q_reg_18_ ( .D(u_csr_csr_satp_r[18]), .CK(clk_i), .RN(
        n44198), .Q(n58074), .QN(n1916) );
  DFFRX1 u_csr_csr_satp_q_reg_17_ ( .D(u_csr_csr_satp_r[17]), .CK(clk_i), .RN(
        n44198), .Q(n73409) );
  DFFRX1 u_csr_csr_satp_q_reg_16_ ( .D(u_csr_csr_satp_r[16]), .CK(clk_i), .RN(
        n44198), .Q(n73410) );
  DFFRX1 u_csr_csr_satp_q_reg_15_ ( .D(u_csr_csr_satp_r[15]), .CK(clk_i), .RN(
        n44198), .Q(n58049), .QN(n1919) );
  DFFRX1 u_csr_csr_satp_q_reg_14_ ( .D(u_csr_csr_satp_r[14]), .CK(clk_i), .RN(
        n44198), .Q(n58041), .QN(n1920) );
  DFFRX1 u_csr_csr_satp_q_reg_13_ ( .D(u_csr_csr_satp_r[13]), .CK(clk_i), .RN(
        n44197), .Q(n58035), .QN(n1921) );
  DFFRX1 u_csr_csr_satp_q_reg_12_ ( .D(u_csr_csr_satp_r[12]), .CK(clk_i), .RN(
        n44197), .Q(n73411) );
  DFFRX1 u_csr_csr_satp_q_reg_11_ ( .D(u_csr_csr_satp_r[11]), .CK(clk_i), .RN(
        n44197), .Q(n73412) );
  DFFRX1 u_csr_csr_satp_q_reg_10_ ( .D(u_csr_csr_satp_r[10]), .CK(clk_i), .RN(
        n44197), .Q(n58014), .QN(n1924) );
  DFFRX1 u_csr_csr_satp_q_reg_0_ ( .D(u_csr_csr_satp_r[0]), .CK(clk_i), .RN(
        n44210), .Q(n57910), .QN(n1925) );
  DFFRX1 u_csr_csr_sr_q_reg_31_ ( .D(u_csr_csr_sr_r[31]), .CK(clk_i), .RN(
        n44151), .Q(u_csr_csr_sr_q_31) );
  DFFRX1 u_csr_csr_sr_q_reg_30_ ( .D(u_csr_csr_sr_r[30]), .CK(clk_i), .RN(
        n44151), .Q(u_csr_csr_sr_q_30) );
  DFFRX1 u_csr_csr_sr_q_reg_29_ ( .D(u_csr_csr_sr_r[29]), .CK(clk_i), .RN(
        n44151), .Q(u_csr_csr_sr_q_29) );
  DFFRX1 u_csr_csr_sr_q_reg_28_ ( .D(u_csr_csr_sr_r[28]), .CK(clk_i), .RN(
        n44151), .Q(u_csr_csr_sr_q_28) );
  DFFRX1 u_csr_csr_sr_q_reg_27_ ( .D(u_csr_csr_sr_r[27]), .CK(clk_i), .RN(
        n44151), .Q(u_csr_csr_sr_q_27) );
  DFFRX1 u_csr_csr_sr_q_reg_26_ ( .D(u_csr_csr_sr_r[26]), .CK(clk_i), .RN(
        n44151), .Q(u_csr_csr_sr_q_26) );
  DFFRX1 u_csr_csr_sr_q_reg_25_ ( .D(u_csr_csr_sr_r[25]), .CK(clk_i), .RN(
        n44151), .Q(u_csr_csr_sr_q_25) );
  DFFRX1 u_csr_csr_sr_q_reg_24_ ( .D(u_csr_csr_sr_r[24]), .CK(clk_i), .RN(
        n44151), .Q(u_csr_csr_sr_q_24) );
  DFFRX1 u_csr_csr_sr_q_reg_23_ ( .D(u_csr_csr_sr_r[23]), .CK(clk_i), .RN(
        n44151), .Q(u_csr_csr_sr_q_23) );
  DFFRX1 u_csr_csr_sscratch_q_reg_9_ ( .D(u_csr_csr_sscratch_r[9]), .CK(clk_i), 
        .RN(n44150), .Q(u_csr_csr_sscratch_q[9]), .QN(n37726) );
  DFFRX1 u_csr_csr_sscratch_q_reg_8_ ( .D(u_csr_csr_sscratch_r[8]), .CK(clk_i), 
        .RN(n44150), .Q(u_csr_csr_sscratch_q[8]), .QN(n37725) );
  DFFRX1 u_csr_csr_sscratch_q_reg_7_ ( .D(u_csr_csr_sscratch_r[7]), .CK(clk_i), 
        .RN(n44150), .Q(u_csr_csr_sscratch_q[7]), .QN(n37724) );
  DFFRX1 u_csr_csr_stvec_q_reg_4_ ( .D(u_csr_csr_stvec_r[4]), .CK(clk_i), .RN(
        n44149), .Q(u_csr_csr_stvec_q[4]), .QN(n37701) );
  DFFRX1 u_csr_csr_stvec_q_reg_3_ ( .D(u_csr_csr_stvec_r[3]), .CK(clk_i), .RN(
        n44149), .Q(u_csr_csr_stvec_q[3]), .QN(n37723) );
  DFFRX1 u_csr_csr_stvec_q_reg_2_ ( .D(u_csr_csr_stvec_r[2]), .CK(clk_i), .RN(
        n44149), .Q(u_csr_csr_stvec_q[2]), .QN(n37703) );
  DFFRX1 u_csr_csr_stvec_q_reg_1_ ( .D(u_csr_csr_stvec_r[1]), .CK(clk_i), .RN(
        n44149), .Q(u_csr_csr_stvec_q[1]), .QN(n37722) );
  DFFRX1 u_csr_csr_stvec_q_reg_0_ ( .D(u_csr_csr_stvec_r[0]), .CK(clk_i), .RN(
        n44148), .Q(u_csr_csr_stvec_q[0]), .QN(n37702) );
  DFFRX1 u_mmu_dtlb_valid_q_reg ( .D(n8504), .CK(clk_i), .RN(n44205), .Q(
        u_mmu_dtlb_valid_q) );
  DFFRX1 u_mmu_itlb_valid_q_reg ( .D(n8505), .CK(clk_i), .RN(n44145), .Q(
        u_mmu_itlb_valid_q) );
  DFFRX1 u_exec_rd_x_q_reg_3_ ( .D(u_exec_N241), .CK(clk_i), .RN(n44128), .Q(
        writeback_exec_idx_w[3]), .QN(n39766) );
  DFFRX1 u_csr_writeback_squash_q_reg ( .D(u_csr_N3472), .CK(clk_i), .RN(
        n44148), .QN(n37332) );
  DFFRX1 u_decode_scoreboard_q_reg_24_ ( .D(u_decode_scoreboard_r[24]), .CK(
        clk_i), .RN(n44148), .Q(u_decode_scoreboard_q[24]) );
  DFFRX1 u_decode_scoreboard_q_reg_25_ ( .D(u_decode_scoreboard_r[25]), .CK(
        clk_i), .RN(n44151), .Q(u_decode_scoreboard_q[25]) );
  DFFRX1 u_decode_scoreboard_q_reg_1_ ( .D(u_decode_scoreboard_r[1]), .CK(
        clk_i), .RN(n44163), .Q(u_decode_scoreboard_q[1]) );
  DFFRX1 u_decode_scoreboard_q_reg_17_ ( .D(u_decode_scoreboard_r[17]), .CK(
        clk_i), .RN(n44163), .Q(u_decode_scoreboard_q[17]) );
  DFFRX1 u_decode_scoreboard_q_reg_5_ ( .D(u_decode_scoreboard_r[5]), .CK(
        clk_i), .RN(n44208), .Q(u_decode_scoreboard_q[5]) );
  DFFRX1 u_decode_scoreboard_q_reg_29_ ( .D(u_decode_scoreboard_r[29]), .CK(
        clk_i), .RN(n44208), .Q(u_decode_scoreboard_q[29]) );
  DFFRX1 u_decode_scoreboard_q_reg_21_ ( .D(u_decode_scoreboard_r[21]), .CK(
        clk_i), .RN(n44208), .Q(u_decode_scoreboard_q[21]), .QN(n37434) );
  DFFRX1 u_decode_scoreboard_q_reg_4_ ( .D(u_decode_scoreboard_r[4]), .CK(
        clk_i), .RN(n44208), .Q(u_decode_scoreboard_q[4]) );
  DFFRX1 u_decode_scoreboard_q_reg_28_ ( .D(u_decode_scoreboard_r[28]), .CK(
        clk_i), .RN(n44208), .Q(u_decode_scoreboard_q[28]) );
  DFFRX1 u_decode_scoreboard_q_reg_20_ ( .D(u_decode_scoreboard_r[20]), .CK(
        clk_i), .RN(n44208), .Q(u_decode_scoreboard_q[20]) );
  DFFRX1 u_decode_scoreboard_q_reg_7_ ( .D(u_decode_scoreboard_r[7]), .CK(
        clk_i), .RN(n44209), .Q(u_decode_scoreboard_q[7]) );
  DFFRX1 u_decode_scoreboard_q_reg_31_ ( .D(u_decode_scoreboard_r[31]), .CK(
        clk_i), .RN(n44209), .Q(u_decode_scoreboard_q[31]) );
  DFFRX1 u_decode_scoreboard_q_reg_23_ ( .D(u_decode_scoreboard_r[23]), .CK(
        clk_i), .RN(n44208), .Q(u_decode_scoreboard_q[23]) );
  DFFRX1 u_decode_scoreboard_q_reg_6_ ( .D(u_decode_scoreboard_r[6]), .CK(
        clk_i), .RN(n44209), .Q(u_decode_scoreboard_q[6]) );
  DFFRX1 u_decode_scoreboard_q_reg_30_ ( .D(u_decode_scoreboard_r[30]), .CK(
        clk_i), .RN(n44208), .Q(u_decode_scoreboard_q[30]), .QN(n40921) );
  DFFRX1 u_decode_scoreboard_q_reg_22_ ( .D(u_decode_scoreboard_r[22]), .CK(
        clk_i), .RN(n44209), .Q(u_decode_scoreboard_q[22]) );
  DFFRX1 u_decode_scoreboard_q_reg_3_ ( .D(u_decode_scoreboard_r[3]), .CK(
        clk_i), .RN(n44207), .Q(u_decode_scoreboard_q[3]) );
  DFFRX1 u_decode_scoreboard_q_reg_27_ ( .D(u_decode_scoreboard_r[27]), .CK(
        clk_i), .RN(n44208), .Q(u_decode_scoreboard_q[27]) );
  DFFRX1 u_decode_scoreboard_q_reg_19_ ( .D(u_decode_scoreboard_r[19]), .CK(
        clk_i), .RN(n44207), .Q(u_decode_scoreboard_q[19]) );
  DFFRX1 u_decode_scoreboard_q_reg_2_ ( .D(u_decode_scoreboard_r[2]), .CK(
        clk_i), .RN(n44208), .Q(u_decode_scoreboard_q[2]), .QN(n37752) );
  DFFRX1 u_decode_scoreboard_q_reg_26_ ( .D(u_decode_scoreboard_r[26]), .CK(
        clk_i), .RN(n44208), .Q(u_decode_scoreboard_q[26]), .QN(n37753) );
  DFFRX1 u_decode_scoreboard_q_reg_18_ ( .D(u_decode_scoreboard_r[18]), .CK(
        clk_i), .RN(n44209), .Q(u_decode_scoreboard_q[18]), .QN(n37756) );
  DFFRX1 u_decode_scoreboard_q_reg_9_ ( .D(u_decode_scoreboard_r[9]), .CK(
        clk_i), .RN(n44163), .Q(u_decode_scoreboard_q[9]) );
  DFFRX1 u_decode_scoreboard_q_reg_15_ ( .D(u_decode_scoreboard_r[15]), .CK(
        clk_i), .RN(n44208), .Q(u_decode_scoreboard_q[15]) );
  DFFRX1 u_decode_scoreboard_q_reg_14_ ( .D(u_decode_scoreboard_r[14]), .CK(
        clk_i), .RN(n44208), .Q(u_decode_scoreboard_q[14]) );
  DFFRX1 u_decode_scoreboard_q_reg_13_ ( .D(u_decode_scoreboard_r[13]), .CK(
        clk_i), .RN(n44208), .Q(u_decode_scoreboard_q[13]) );
  DFFRX1 u_decode_scoreboard_q_reg_12_ ( .D(u_decode_scoreboard_r[12]), .CK(
        clk_i), .RN(n44208), .Q(u_decode_scoreboard_q[12]) );
  DFFRX1 u_decode_scoreboard_q_reg_11_ ( .D(u_decode_scoreboard_r[11]), .CK(
        clk_i), .RN(n44208), .Q(u_decode_scoreboard_q[11]), .QN(n37754) );
  DFFRX1 u_decode_scoreboard_q_reg_10_ ( .D(u_decode_scoreboard_r[10]), .CK(
        clk_i), .RN(n44208), .Q(u_decode_scoreboard_q[10]), .QN(n37755) );
  DFFRX1 u_decode_scoreboard_q_reg_8_ ( .D(u_decode_scoreboard_r[8]), .CK(
        clk_i), .RN(n44163), .Q(u_decode_scoreboard_q[8]) );
  DFFRX1 u_muldiv_div_inst_q_reg ( .D(n8521), .CK(clk_i), .RN(n44163), .Q(
        u_muldiv_div_inst_q), .QN(n37586) );
  DFFRX1 u_csr_csr_sr_q_reg_7_ ( .D(u_csr_csr_sr_r_7), .CK(clk_i), .RN(n44163), 
        .Q(u_csr_csr_sr_q[7]), .QN(n37750) );
  DFFRX1 u_csr_csr_sr_q_reg_3_ ( .D(u_csr_csr_sr_r_3), .CK(clk_i), .RN(n44163), 
        .Q(u_csr_csr_sr_q[3]), .QN(n37748) );
  DFFRX1 u_csr_csr_scause_q_reg_3_ ( .D(u_csr_csr_scause_r[3]), .CK(clk_i), 
        .RN(n44163), .Q(u_csr_csr_scause_q[3]) );
  DFFRX1 u_csr_csr_scause_q_reg_31_ ( .D(u_csr_csr_scause_r_31), .CK(clk_i), 
        .RN(n44163), .Q(u_csr_csr_scause_q_31) );
  DFFRX1 u_csr_csr_mcause_q_reg_31_ ( .D(u_csr_csr_mcause_r_31), .CK(clk_i), 
        .RN(n44163), .Q(u_csr_csr_mcause_q_31) );
  DFFRX1 u_csr_csr_scause_q_reg_2_ ( .D(u_csr_csr_scause_r[2]), .CK(clk_i), 
        .RN(n44163), .QN(n37728) );
  DFFRX1 u_csr_csr_mcause_q_reg_2_ ( .D(u_csr_csr_mcause_r[2]), .CK(clk_i), 
        .RN(n44163), .Q(u_csr_csr_mcause_q[2]), .QN(n37775) );
  DFFRX1 u_csr_csr_sr_q_reg_8_ ( .D(u_csr_csr_sr_r_8), .CK(clk_i), .RN(n44162), 
        .Q(u_csr_csr_sr_q[8]), .QN(n37663) );
  DFFRX1 u_csr_csr_sr_q_reg_1_ ( .D(u_csr_csr_sr_r_1), .CK(clk_i), .RN(n44162), 
        .Q(u_csr_csr_sr_q[1]), .QN(n37540) );
  DFFRX1 u_csr_csr_sr_q_reg_5_ ( .D(u_csr_csr_sr_r_5), .CK(clk_i), .RN(n44162), 
        .Q(u_csr_csr_sr_q[5]), .QN(n37751) );
  DFFRX1 u_csr_csr_mcause_q_reg_3_ ( .D(u_csr_csr_mcause_r[3]), .CK(clk_i), 
        .RN(n44162), .Q(u_csr_csr_mcause_q[3]) );
  DFFRX1 u_csr_csr_scause_q_reg_1_ ( .D(u_csr_csr_scause_r[1]), .CK(clk_i), 
        .RN(n44162), .Q(u_csr_csr_scause_q[1]), .QN(n37762) );
  DFFRX1 u_csr_csr_mcause_q_reg_1_ ( .D(u_csr_csr_mcause_r[1]), .CK(clk_i), 
        .RN(n44162), .Q(u_csr_csr_mcause_q[1]) );
  DFFRX1 u_csr_csr_scause_q_reg_0_ ( .D(u_csr_csr_scause_r[0]), .CK(clk_i), 
        .RN(n44162), .QN(n37727) );
  DFFRX1 u_csr_csr_mcause_q_reg_0_ ( .D(u_csr_csr_mcause_r[0]), .CK(clk_i), 
        .RN(n44162), .Q(u_csr_csr_mcause_q[0]) );
  DFFRX1 u_csr_branch_target_q_reg_11_ ( .D(u_csr_N3676), .CK(clk_i), .RN(
        n44104), .Q(n55016) );
  DFFRX1 u_fetch_branch_pc_q_reg_11_ ( .D(net2292), .CK(n37867), .RN(n44105), 
        .QN(n1931) );
  DFFRX1 u_csr_pc_m_q_reg_11_ ( .D(opcode_pc_w[11]), .CK(net1872), .RN(n44104), 
        .QN(n37769) );
  DFFRX1 u_csr_branch_target_q_reg_29_ ( .D(u_csr_N3694), .CK(clk_i), .RN(
        n44196), .Q(n56349) );
  DFFRX1 u_csr_branch_target_q_reg_28_ ( .D(u_csr_N3693), .CK(clk_i), .RN(
        n44193), .Q(n56166) );
  DFFRX1 u_fetch_branch_pc_q_reg_28_ ( .D(net2314), .CK(n37866), .RN(n44193), 
        .QN(n1936) );
  DFFRX1 u_csr_branch_target_q_reg_27_ ( .D(u_csr_N3692), .CK(clk_i), .RN(
        n44191), .Q(n55989) );
  DFFRX1 u_fetch_branch_pc_q_reg_27_ ( .D(net2313), .CK(n37866), .RN(n44191), 
        .QN(n1938) );
  DFFRX1 u_csr_branch_target_q_reg_0_ ( .D(u_csr_N3665), .CK(clk_i), .RN(
        n44204), .Q(n57273), .QN(n8848) );
  DFFRX1 u_csr_pc_m_q_reg_0_ ( .D(u_csr_N184), .CK(net1867), .RN(n44204), .QN(
        n37747) );
  DFFRX1 u_csr_csr_stval_q_reg_0_ ( .D(u_csr_csr_stval_r[0]), .CK(clk_i), .RN(
        n44162), .Q(u_csr_csr_stval_q[0]) );
  DFFRX1 u_decode_u_regfile_reg_r1_q_reg_0_ ( .D(u_decode_u_regfile_N100), 
        .CK(n37865), .RN(n44123), .Q(n1943), .QN(n37304) );
  DFFRX1 u_decode_u_regfile_reg_r26_q_reg_0_ ( .D(u_decode_u_regfile_N1025), 
        .CK(n37864), .RN(n44130), .Q(n1944) );
  DFFRX1 u_decode_u_regfile_reg_r27_q_reg_0_ ( .D(u_decode_u_regfile_N1062), 
        .CK(n37863), .RN(n44131), .Q(n1945) );
  DFFRX1 u_decode_u_regfile_reg_r28_q_reg_0_ ( .D(u_decode_u_regfile_N1099), 
        .CK(n37862), .RN(n44130), .Q(n1946), .QN(n37226) );
  DFFRX1 u_decode_u_regfile_reg_r29_q_reg_0_ ( .D(u_decode_u_regfile_N1136), 
        .CK(n37861), .RN(n44131), .Q(n1947), .QN(n36812) );
  DFFRX1 u_decode_u_regfile_reg_r30_q_reg_0_ ( .D(u_decode_u_regfile_N1173), 
        .CK(n37860), .RN(n44131), .Q(n1948), .QN(n37218) );
  DFFRX1 u_decode_u_regfile_reg_r31_q_reg_0_ ( .D(u_decode_u_regfile_N1210), 
        .CK(n37859), .RN(n44130), .Q(n1949), .QN(n37219) );
  DFFRX1 u_decode_u_regfile_reg_r2_q_reg_0_ ( .D(u_decode_u_regfile_N137), 
        .CK(n37858), .RN(n44130), .Q(n1950) );
  DFFRX1 u_decode_u_regfile_reg_r3_q_reg_0_ ( .D(u_decode_u_regfile_N174), 
        .CK(n37857), .RN(n44131), .Q(n1951), .QN(n37299) );
  DFFRX1 u_decode_u_regfile_reg_r4_q_reg_0_ ( .D(u_decode_u_regfile_N211), 
        .CK(n37856), .RN(n44130), .Q(n1952) );
  DFFRX1 u_decode_u_regfile_reg_r6_q_reg_0_ ( .D(u_decode_u_regfile_N285), 
        .CK(n37855), .RN(n44130), .Q(n1954) );
  DFFRX1 u_decode_u_regfile_reg_r7_q_reg_0_ ( .D(u_decode_u_regfile_N322), 
        .CK(n37854), .RN(n44130), .Q(n1955), .QN(n37222) );
  DFFRX1 u_decode_u_regfile_reg_r9_q_reg_0_ ( .D(u_decode_u_regfile_N396), 
        .CK(n37853), .RN(n44131), .Q(n1957), .QN(n37301) );
  DFFRX1 u_decode_u_regfile_reg_r10_q_reg_0_ ( .D(u_decode_u_regfile_N433), 
        .CK(n37852), .RN(n44131), .Q(n1958) );
  DFFRX1 u_decode_u_regfile_reg_r11_q_reg_0_ ( .D(u_decode_u_regfile_N470), 
        .CK(n37851), .RN(n44131), .Q(n1959), .QN(n37300) );
  DFFRX1 u_decode_u_regfile_reg_r12_q_reg_0_ ( .D(u_decode_u_regfile_N507), 
        .CK(n37850), .RN(n44131), .Q(n1960) );
  DFFRX1 u_decode_u_regfile_reg_r13_q_reg_0_ ( .D(u_decode_u_regfile_N544), 
        .CK(n37849), .RN(n44131), .Q(n1961) );
  DFFRX1 u_decode_u_regfile_reg_r14_q_reg_0_ ( .D(u_decode_u_regfile_N581), 
        .CK(n37848), .RN(n44131), .Q(n1962) );
  DFFRX1 u_decode_u_regfile_reg_r15_q_reg_0_ ( .D(u_decode_u_regfile_N618), 
        .CK(n37847), .RN(n44131), .Q(n1963) );
  DFFRX1 u_decode_u_regfile_reg_r16_q_reg_0_ ( .D(u_decode_u_regfile_N655), 
        .CK(n37846), .RN(n44131), .Q(n1964), .QN(n42509) );
  DFFRX1 u_decode_u_regfile_reg_r17_q_reg_0_ ( .D(u_decode_u_regfile_N692), 
        .CK(n37845), .RN(n44131), .Q(n1965), .QN(n37302) );
  DFFRX1 u_decode_u_regfile_reg_r18_q_reg_0_ ( .D(u_decode_u_regfile_N729), 
        .CK(n37844), .RN(n44130), .QN(n36799) );
  DFFRX1 u_decode_u_regfile_reg_r19_q_reg_0_ ( .D(u_decode_u_regfile_N766), 
        .CK(n37843), .RN(n44131), .Q(n1967), .QN(n37298) );
  DFFRX1 u_decode_u_regfile_reg_r20_q_reg_0_ ( .D(u_decode_u_regfile_N803), 
        .CK(n37842), .RN(n44131), .Q(n1968), .QN(n37220) );
  DFFRX1 u_decode_u_regfile_reg_r22_q_reg_0_ ( .D(u_decode_u_regfile_N877), 
        .CK(n37841), .RN(n44131), .Q(n1970), .QN(n37217) );
  DFFRX1 u_decode_u_regfile_reg_r23_q_reg_0_ ( .D(u_decode_u_regfile_N914), 
        .CK(n37877), .RN(n44131), .Q(n1971) );
  DFFRX1 u_csr_branch_target_q_reg_1_ ( .D(u_csr_N3666), .CK(clk_i), .RN(
        n44145), .Q(n56772), .QN(n8836) );
  DFFRX1 u_fetch_branch_pc_q_reg_1_ ( .D(net2282), .CK(n37867), .RN(n44145), 
        .QN(n1972) );
  DFFRX1 u_csr_pc_m_q_reg_1_ ( .D(opcode_pc_w[1]), .CK(net1867), .RN(n44145), 
        .QN(n37746) );
  DFFRX1 u_csr_csr_stval_q_reg_1_ ( .D(u_csr_csr_stval_r[1]), .CK(clk_i), .RN(
        n44162), .Q(u_csr_csr_stval_q[1]) );
  DFFRX1 u_decode_u_regfile_reg_r1_q_reg_1_ ( .D(u_decode_u_regfile_N101), 
        .CK(n37865), .RN(n44121), .QN(n36820) );
  DFFRX1 u_decode_u_regfile_reg_r26_q_reg_1_ ( .D(u_decode_u_regfile_N1026), 
        .CK(n37864), .RN(n44120), .Q(n1976) );
  DFFRX1 u_decode_u_regfile_reg_r28_q_reg_1_ ( .D(u_decode_u_regfile_N1100), 
        .CK(n37862), .RN(n44120), .Q(n1978) );
  DFFRX1 u_decode_u_regfile_reg_r29_q_reg_1_ ( .D(u_decode_u_regfile_N1137), 
        .CK(n37861), .RN(n44119), .QN(n36815) );
  DFFRX1 u_decode_u_regfile_reg_r30_q_reg_1_ ( .D(u_decode_u_regfile_N1174), 
        .CK(n37860), .RN(n44120), .Q(n1980) );
  DFFRX1 u_decode_u_regfile_reg_r31_q_reg_1_ ( .D(u_decode_u_regfile_N1211), 
        .CK(n37859), .RN(n44119), .Q(n1981), .QN(n37196) );
  DFFRX1 u_decode_u_regfile_reg_r2_q_reg_1_ ( .D(u_decode_u_regfile_N138), 
        .CK(n37858), .RN(n44120), .Q(n1982) );
  DFFRX1 u_decode_u_regfile_reg_r4_q_reg_1_ ( .D(u_decode_u_regfile_N212), 
        .CK(n37856), .RN(n44120), .Q(n1984) );
  DFFRX1 u_decode_u_regfile_reg_r5_q_reg_1_ ( .D(u_decode_u_regfile_N249), 
        .CK(n37840), .RN(n44120), .Q(n1985), .QN(n36801) );
  DFFRX1 u_decode_u_regfile_reg_r6_q_reg_1_ ( .D(u_decode_u_regfile_N286), 
        .CK(n37855), .RN(n44120), .QN(n36810) );
  DFFRX1 u_decode_u_regfile_reg_r7_q_reg_1_ ( .D(u_decode_u_regfile_N323), 
        .CK(n37854), .RN(n44120), .QN(n36862) );
  DFFRX1 u_decode_u_regfile_reg_r8_q_reg_1_ ( .D(u_decode_u_regfile_N360), 
        .CK(n37839), .RN(n44121), .Q(n1988), .QN(n37294) );
  DFFRX1 u_decode_u_regfile_reg_r9_q_reg_1_ ( .D(u_decode_u_regfile_N397), 
        .CK(n37853), .RN(n44121), .Q(n1989), .QN(n37296) );
  DFFRX1 u_decode_u_regfile_reg_r10_q_reg_1_ ( .D(u_decode_u_regfile_N434), 
        .CK(n37852), .RN(n44120), .Q(n1990) );
  DFFRX1 u_decode_u_regfile_reg_r12_q_reg_1_ ( .D(u_decode_u_regfile_N508), 
        .CK(n37850), .RN(n44120), .Q(n1992) );
  DFFRX1 u_decode_u_regfile_reg_r13_q_reg_1_ ( .D(u_decode_u_regfile_N545), 
        .CK(n37849), .RN(n44120), .QN(n36814) );
  DFFRX1 u_decode_u_regfile_reg_r15_q_reg_1_ ( .D(u_decode_u_regfile_N619), 
        .CK(n37847), .RN(n44120), .Q(n1995), .QN(n37198) );
  DFFRX1 u_decode_u_regfile_reg_r16_q_reg_1_ ( .D(u_decode_u_regfile_N656), 
        .CK(n37846), .RN(n44121), .Q(n1996), .QN(n37295) );
  DFFRX1 u_decode_u_regfile_reg_r17_q_reg_1_ ( .D(u_decode_u_regfile_N693), 
        .CK(n37845), .RN(n44121), .Q(n1997), .QN(n37297) );
  DFFRX1 u_decode_u_regfile_reg_r20_q_reg_1_ ( .D(u_decode_u_regfile_N804), 
        .CK(n37842), .RN(n44120), .Q(n2000) );
  DFFRX1 u_decode_u_regfile_reg_r22_q_reg_1_ ( .D(u_decode_u_regfile_N878), 
        .CK(n37841), .RN(n44120), .Q(n2002), .QN(n37201) );
  DFFRX1 u_decode_u_regfile_reg_r23_q_reg_1_ ( .D(u_decode_u_regfile_N915), 
        .CK(n37877), .RN(n44120), .Q(n2003), .QN(n37211) );
  DFFRX1 u_csr_branch_target_q_reg_2_ ( .D(u_csr_N3667), .CK(clk_i), .RN(
        n44117), .Q(n54431), .QN(n8845) );
  DFFRX1 u_fetch_branch_pc_q_reg_2_ ( .D(net2283), .CK(n37867), .RN(n44117), 
        .QN(n2004) );
  DFFRX1 u_csr_csr_stval_q_reg_2_ ( .D(u_csr_csr_stval_r[2]), .CK(clk_i), .RN(
        n44162), .Q(u_csr_csr_stval_q[2]) );
  DFFRX1 u_decode_u_regfile_reg_r1_q_reg_2_ ( .D(u_decode_u_regfile_N102), 
        .CK(n37865), .RN(n44132), .Q(n2006), .QN(n37313) );
  DFFRX1 u_decode_u_regfile_reg_r26_q_reg_2_ ( .D(u_decode_u_regfile_N1027), 
        .CK(n37864), .RN(n44132), .Q(n2007) );
  DFFRX1 u_decode_u_regfile_reg_r27_q_reg_2_ ( .D(u_decode_u_regfile_N1064), 
        .CK(n37863), .RN(n44132), .Q(n2008) );
  DFFRX1 u_decode_u_regfile_reg_r28_q_reg_2_ ( .D(u_decode_u_regfile_N1101), 
        .CK(n37862), .RN(n44132), .Q(n2009), .QN(n37240) );
  DFFRX1 u_decode_u_regfile_reg_r29_q_reg_2_ ( .D(u_decode_u_regfile_N1138), 
        .CK(n37861), .RN(n44147), .Q(n2010) );
  DFFRX1 u_decode_u_regfile_reg_r30_q_reg_2_ ( .D(u_decode_u_regfile_N1175), 
        .CK(n37860), .RN(n44147), .Q(n2011), .QN(n37234) );
  DFFRX1 u_decode_u_regfile_reg_r31_q_reg_2_ ( .D(u_decode_u_regfile_N1212), 
        .CK(n37859), .RN(n44205), .Q(n2012), .QN(n37235) );
  DFFRX1 u_decode_u_regfile_reg_r2_q_reg_2_ ( .D(u_decode_u_regfile_N139), 
        .CK(n37858), .RN(n44148), .Q(n2013) );
  DFFRX1 u_decode_u_regfile_reg_r3_q_reg_2_ ( .D(u_decode_u_regfile_N176), 
        .CK(n37857), .RN(n44148), .Q(n2014), .QN(n37306) );
  DFFRX1 u_decode_u_regfile_reg_r4_q_reg_2_ ( .D(u_decode_u_regfile_N213), 
        .CK(n37856), .RN(n44148), .Q(n2015) );
  DFFRX1 u_decode_u_regfile_reg_r5_q_reg_2_ ( .D(u_decode_u_regfile_N250), 
        .CK(n37840), .RN(n44148), .Q(n2016) );
  DFFRX1 u_decode_u_regfile_reg_r6_q_reg_2_ ( .D(u_decode_u_regfile_N287), 
        .CK(n37855), .RN(n44136), .Q(n2017) );
  DFFRX1 u_decode_u_regfile_reg_r7_q_reg_2_ ( .D(u_decode_u_regfile_N324), 
        .CK(n37854), .RN(n44148), .Q(n2018), .QN(n37238) );
  DFFRX1 u_decode_u_regfile_reg_r8_q_reg_2_ ( .D(u_decode_u_regfile_N361), 
        .CK(n37839), .RN(n44132), .Q(n2019), .QN(n37307) );
  DFFRX1 u_decode_u_regfile_reg_r9_q_reg_2_ ( .D(u_decode_u_regfile_N398), 
        .CK(n37853), .RN(n44147), .Q(n2020), .QN(n42496) );
  DFFRX1 u_decode_u_regfile_reg_r10_q_reg_2_ ( .D(u_decode_u_regfile_N435), 
        .CK(n37852), .RN(n44132), .Q(n2021) );
  DFFRX1 u_decode_u_regfile_reg_r11_q_reg_2_ ( .D(u_decode_u_regfile_N472), 
        .CK(n37851), .RN(n44132), .Q(n2022), .QN(n37308) );
  DFFRX1 u_decode_u_regfile_reg_r12_q_reg_2_ ( .D(u_decode_u_regfile_N509), 
        .CK(n37850), .RN(n44132), .Q(n2023) );
  DFFRX1 u_decode_u_regfile_reg_r13_q_reg_2_ ( .D(u_decode_u_regfile_N546), 
        .CK(n37849), .RN(n44132), .Q(n2024) );
  DFFRX1 u_decode_u_regfile_reg_r14_q_reg_2_ ( .D(u_decode_u_regfile_N583), 
        .CK(n37848), .RN(n44132), .Q(n2025) );
  DFFRX1 u_decode_u_regfile_reg_r15_q_reg_2_ ( .D(u_decode_u_regfile_N620), 
        .CK(n37847), .RN(n44132), .Q(n2026) );
  DFFRX1 u_decode_u_regfile_reg_r16_q_reg_2_ ( .D(u_decode_u_regfile_N657), 
        .CK(n37846), .RN(n44132), .Q(n2027), .QN(n37309) );
  DFFRX1 u_decode_u_regfile_reg_r17_q_reg_2_ ( .D(u_decode_u_regfile_N694), 
        .CK(n37845), .RN(n44132), .Q(n2028), .QN(n37311) );
  DFFRX1 u_decode_u_regfile_reg_r18_q_reg_2_ ( .D(u_decode_u_regfile_N731), 
        .CK(n37844), .RN(n44147), .Q(n2029), .QN(n37239) );
  DFFRX1 u_decode_u_regfile_reg_r19_q_reg_2_ ( .D(u_decode_u_regfile_N768), 
        .CK(n37843), .RN(n44147), .Q(n2030), .QN(n37305) );
  DFFRX1 u_decode_u_regfile_reg_r20_q_reg_2_ ( .D(u_decode_u_regfile_N805), 
        .CK(n37842), .RN(n44148), .Q(n2031), .QN(n37236) );
  DFFRX1 u_decode_u_regfile_reg_r21_q_reg_2_ ( .D(u_decode_u_regfile_N842), 
        .CK(n37838), .RN(n44147), .Q(n2032), .QN(n37237) );
  DFFRX1 u_decode_u_regfile_reg_r22_q_reg_2_ ( .D(u_decode_u_regfile_N879), 
        .CK(n37841), .RN(n44148), .Q(n2033), .QN(n37233) );
  DFFRX1 u_decode_u_regfile_reg_r23_q_reg_2_ ( .D(u_decode_u_regfile_N916), 
        .CK(n37877), .RN(n44147), .Q(n2034) );
  DFFRX1 u_csr_branch_target_q_reg_3_ ( .D(u_csr_N3668), .CK(clk_i), .RN(
        n44117), .Q(n54564) );
  DFFRX1 u_fetch_branch_pc_q_reg_3_ ( .D(net2284), .CK(n37867), .RN(n44117), 
        .QN(n2035) );
  DFFRX1 u_csr_csr_stval_q_reg_3_ ( .D(u_csr_csr_stval_r[3]), .CK(clk_i), .RN(
        n44162), .Q(u_csr_csr_stval_q[3]) );
  DFFRX1 u_decode_u_regfile_reg_r26_q_reg_3_ ( .D(u_decode_u_regfile_N1028), 
        .CK(n37864), .RN(n44128), .Q(n2037) );
  DFFRX1 u_decode_u_regfile_reg_r1_q_reg_3_ ( .D(u_decode_u_regfile_N103), 
        .CK(n37865), .RN(n44130), .QN(n36902) );
  DFFRX1 u_decode_u_regfile_reg_r27_q_reg_3_ ( .D(u_decode_u_regfile_N1065), 
        .CK(n37863), .RN(n44130), .Q(n2039), .QN(n36907) );
  DFFRX1 u_decode_u_regfile_reg_r28_q_reg_3_ ( .D(u_decode_u_regfile_N1102), 
        .CK(n37862), .RN(n44129), .Q(n2040), .QN(n37147) );
  DFFRX1 u_decode_u_regfile_reg_r29_q_reg_3_ ( .D(u_decode_u_regfile_N1139), 
        .CK(n37861), .RN(n44129), .Q(n2041), .QN(n36901) );
  DFFRX1 u_decode_u_regfile_reg_r30_q_reg_3_ ( .D(u_decode_u_regfile_N1176), 
        .CK(n37860), .RN(n44129), .Q(n2042), .QN(n37140) );
  DFFRX1 u_decode_u_regfile_reg_r31_q_reg_3_ ( .D(u_decode_u_regfile_N1213), 
        .CK(n37859), .RN(n44128), .QN(n37032) );
  DFFRX1 u_decode_u_regfile_reg_r2_q_reg_3_ ( .D(u_decode_u_regfile_N140), 
        .CK(n37858), .RN(n44128), .Q(n2044), .QN(n40893) );
  DFFRX1 u_decode_u_regfile_reg_r3_q_reg_3_ ( .D(u_decode_u_regfile_N177), 
        .CK(n37857), .RN(n44130), .QN(n36900) );
  DFFRX1 u_decode_u_regfile_reg_r4_q_reg_3_ ( .D(u_decode_u_regfile_N214), 
        .CK(n37856), .RN(n44129), .Q(n2046), .QN(n40879) );
  DFFRX1 u_decode_u_regfile_reg_r5_q_reg_3_ ( .D(u_decode_u_regfile_N251), 
        .CK(n37840), .RN(n44129), .Q(n2047), .QN(n37047) );
  DFFRX1 u_decode_u_regfile_reg_r6_q_reg_3_ ( .D(u_decode_u_regfile_N288), 
        .CK(n37855), .RN(n44129), .Q(n2048), .QN(n36909) );
  DFFRX1 u_decode_u_regfile_reg_r7_q_reg_3_ ( .D(u_decode_u_regfile_N325), 
        .CK(n37854), .RN(n44128), .QN(n37093) );
  DFFRX1 u_decode_u_regfile_reg_r8_q_reg_3_ ( .D(u_decode_u_regfile_N362), 
        .CK(n37839), .RN(n44130), .QN(n37092) );
  DFFRX1 u_decode_u_regfile_reg_r9_q_reg_3_ ( .D(u_decode_u_regfile_N399), 
        .CK(n37853), .RN(n44129), .QN(n36898) );
  DFFRX1 u_decode_u_regfile_reg_r10_q_reg_3_ ( .D(u_decode_u_regfile_N436), 
        .CK(n37852), .RN(n44129), .Q(n2052), .QN(n40871) );
  DFFRX1 u_decode_u_regfile_reg_r11_q_reg_3_ ( .D(u_decode_u_regfile_N473), 
        .CK(n37851), .RN(n44130), .QN(n37024) );
  DFFRX1 u_decode_u_regfile_reg_r12_q_reg_3_ ( .D(u_decode_u_regfile_N510), 
        .CK(n37850), .RN(n44129), .Q(n2054), .QN(n40863) );
  DFFRX1 u_decode_u_regfile_reg_r13_q_reg_3_ ( .D(u_decode_u_regfile_N547), 
        .CK(n37849), .RN(n44129), .Q(n2055), .QN(n36904) );
  DFFRX1 u_decode_u_regfile_reg_r14_q_reg_3_ ( .D(u_decode_u_regfile_N584), 
        .CK(n37848), .RN(n44129), .Q(n2056), .QN(n36910) );
  DFFRX1 u_decode_u_regfile_reg_r15_q_reg_3_ ( .D(u_decode_u_regfile_N621), 
        .CK(n37847), .RN(n44129), .Q(n2057), .QN(n37040) );
  DFFRX1 u_decode_u_regfile_reg_r16_q_reg_3_ ( .D(u_decode_u_regfile_N658), 
        .CK(n37846), .RN(n44129), .QN(n37028) );
  DFFRX1 u_decode_u_regfile_reg_r17_q_reg_3_ ( .D(u_decode_u_regfile_N695), 
        .CK(n37845), .RN(n44130), .QN(n36913) );
  DFFRX1 u_decode_u_regfile_reg_r18_q_reg_3_ ( .D(u_decode_u_regfile_N732), 
        .CK(n37844), .RN(n44129), .QN(n36897) );
  DFFRX1 u_decode_u_regfile_reg_r19_q_reg_3_ ( .D(u_decode_u_regfile_N769), 
        .CK(n37843), .RN(n44130), .QN(n36899) );
  DFFRX1 u_decode_u_regfile_reg_r20_q_reg_3_ ( .D(u_decode_u_regfile_N806), 
        .CK(n37842), .RN(n44129), .QN(n36893) );
  DFFRX1 u_decode_u_regfile_reg_r21_q_reg_3_ ( .D(u_decode_u_regfile_N843), 
        .CK(n37838), .RN(n44129), .QN(n36903) );
  DFFRX1 u_decode_u_regfile_reg_r22_q_reg_3_ ( .D(u_decode_u_regfile_N880), 
        .CK(n37841), .RN(n44129), .QN(n36905) );
  DFFRX1 u_decode_u_regfile_reg_r23_q_reg_3_ ( .D(u_decode_u_regfile_N917), 
        .CK(n37877), .RN(n44129), .Q(n2065), .QN(n37039) );
  DFFRX1 u_csr_branch_target_q_reg_4_ ( .D(u_csr_N3669), .CK(clk_i), .RN(
        n44117), .Q(n54571) );
  DFFRX1 u_fetch_branch_pc_q_reg_4_ ( .D(net2285), .CK(n37867), .RN(n44117), 
        .QN(n2066) );
  DFFRX1 u_csr_pc_m_q_reg_4_ ( .D(opcode_pc_w[4]), .CK(net1867), .RN(n44117), 
        .QN(n37763) );
  DFFRX1 u_csr_csr_stval_q_reg_4_ ( .D(u_csr_csr_stval_r[4]), .CK(clk_i), .RN(
        n44162), .Q(u_csr_csr_stval_q[4]) );
  DFFRX1 u_decode_u_regfile_reg_r26_q_reg_4_ ( .D(u_decode_u_regfile_N1029), 
        .CK(n37864), .RN(n44146), .Q(n2069) );
  DFFRX1 u_decode_u_regfile_reg_r1_q_reg_4_ ( .D(u_decode_u_regfile_N104), 
        .CK(n37865), .RN(n44146), .QN(n36947) );
  DFFRX1 u_decode_u_regfile_reg_r27_q_reg_4_ ( .D(u_decode_u_regfile_N1066), 
        .CK(n37863), .RN(n44147), .Q(n2071), .QN(n40881) );
  DFFRX1 u_decode_u_regfile_reg_r28_q_reg_4_ ( .D(u_decode_u_regfile_N1103), 
        .CK(n37862), .RN(n44146), .Q(n2072), .QN(n37149) );
  DFFRX1 u_decode_u_regfile_reg_r29_q_reg_4_ ( .D(u_decode_u_regfile_N1140), 
        .CK(n37861), .RN(n44147), .Q(n2073), .QN(n36941) );
  DFFRX1 u_decode_u_regfile_reg_r30_q_reg_4_ ( .D(u_decode_u_regfile_N1177), 
        .CK(n37860), .RN(n44146), .Q(n2074), .QN(n37141) );
  DFFRX1 u_decode_u_regfile_reg_r31_q_reg_4_ ( .D(u_decode_u_regfile_N1214), 
        .CK(n37859), .RN(n44187), .QN(n36942) );
  DFFRX1 u_decode_u_regfile_reg_r2_q_reg_4_ ( .D(u_decode_u_regfile_N141), 
        .CK(n37858), .RN(n44146), .Q(n2076) );
  DFFRX1 u_decode_u_regfile_reg_r3_q_reg_4_ ( .D(u_decode_u_regfile_N178), 
        .CK(n37857), .RN(n44147), .QN(n36949) );
  DFFRX1 u_decode_u_regfile_reg_r4_q_reg_4_ ( .D(u_decode_u_regfile_N215), 
        .CK(n37856), .RN(n44146), .Q(n2078) );
  DFFRX1 u_decode_u_regfile_reg_r5_q_reg_4_ ( .D(u_decode_u_regfile_N252), 
        .CK(n37840), .RN(n44147), .Q(n2079), .QN(n36965) );
  DFFRX1 u_decode_u_regfile_reg_r6_q_reg_4_ ( .D(u_decode_u_regfile_N289), 
        .CK(n37855), .RN(n44146), .Q(n2080) );
  DFFRX1 u_decode_u_regfile_reg_r7_q_reg_4_ ( .D(u_decode_u_regfile_N326), 
        .CK(n37854), .RN(n44147), .Q(n2081), .QN(n37145) );
  DFFRX1 u_decode_u_regfile_reg_r8_q_reg_4_ ( .D(u_decode_u_regfile_N363), 
        .CK(n37839), .RN(n44146), .Q(n2082), .QN(n37291) );
  DFFRX1 u_decode_u_regfile_reg_r9_q_reg_4_ ( .D(u_decode_u_regfile_N400), 
        .CK(n37853), .RN(n44146), .QN(n36969) );
  DFFRX1 u_decode_u_regfile_reg_r10_q_reg_4_ ( .D(u_decode_u_regfile_N437), 
        .CK(n37852), .RN(n44146), .Q(n2084) );
  DFFRX1 u_decode_u_regfile_reg_r11_q_reg_4_ ( .D(u_decode_u_regfile_N474), 
        .CK(n37851), .RN(n44147), .QN(n36945) );
  DFFRX1 u_decode_u_regfile_reg_r12_q_reg_4_ ( .D(u_decode_u_regfile_N511), 
        .CK(n37850), .RN(n44146), .Q(n2086) );
  DFFRX1 u_decode_u_regfile_reg_r13_q_reg_4_ ( .D(u_decode_u_regfile_N548), 
        .CK(n37849), .RN(n44147), .Q(n2087), .QN(n40901) );
  DFFRX1 u_decode_u_regfile_reg_r14_q_reg_4_ ( .D(u_decode_u_regfile_N585), 
        .CK(n37848), .RN(n44146), .Q(n2088) );
  DFFRX1 u_decode_u_regfile_reg_r15_q_reg_4_ ( .D(u_decode_u_regfile_N622), 
        .CK(n37847), .RN(n44147), .Q(n2089), .QN(n36966) );
  DFFRX1 u_decode_u_regfile_reg_r16_q_reg_4_ ( .D(u_decode_u_regfile_N659), 
        .CK(n37846), .RN(n44145), .Q(n2090), .QN(n42501) );
  DFFRX1 u_decode_u_regfile_reg_r17_q_reg_4_ ( .D(u_decode_u_regfile_N696), 
        .CK(n37845), .RN(n44146), .QN(n36961) );
  DFFRX1 u_decode_u_regfile_reg_r18_q_reg_4_ ( .D(u_decode_u_regfile_N733), 
        .CK(n37844), .RN(n44146), .Q(n2092), .QN(n37146) );
  DFFRX1 u_decode_u_regfile_reg_r19_q_reg_4_ ( .D(u_decode_u_regfile_N770), 
        .CK(n37843), .RN(n44147), .QN(n36982) );
  DFFRX1 u_decode_u_regfile_reg_r20_q_reg_4_ ( .D(u_decode_u_regfile_N807), 
        .CK(n37842), .RN(n44146), .Q(n2094), .QN(n37143) );
  DFFRX1 u_decode_u_regfile_reg_r21_q_reg_4_ ( .D(u_decode_u_regfile_N844), 
        .CK(n37838), .RN(n44147), .QN(n36944) );
  DFFRX1 u_decode_u_regfile_reg_r22_q_reg_4_ ( .D(u_decode_u_regfile_N881), 
        .CK(n37841), .RN(n44146), .Q(n2096), .QN(n37138) );
  DFFRX1 u_decode_u_regfile_reg_r23_q_reg_4_ ( .D(u_decode_u_regfile_N918), 
        .CK(n37877), .RN(n44147), .Q(n2097), .QN(n36936) );
  DFFRX1 u_csr_branch_target_q_reg_5_ ( .D(u_csr_N3670), .CK(clk_i), .RN(
        n44118), .Q(n54642) );
  DFFRX1 u_fetch_branch_pc_q_reg_5_ ( .D(net2286), .CK(n37867), .RN(n44118), 
        .QN(n2098) );
  DFFRX1 u_csr_pc_m_q_reg_5_ ( .D(opcode_pc_w[5]), .CK(net1867), .RN(n44118), 
        .QN(n37765) );
  DFFRX1 u_decode_u_regfile_reg_r26_q_reg_5_ ( .D(u_decode_u_regfile_N1030), 
        .CK(n37864), .RN(n44143), .Q(n2101) );
  DFFRX1 u_decode_u_regfile_reg_r1_q_reg_5_ ( .D(u_decode_u_regfile_N105), 
        .CK(n37865), .RN(n44145), .Q(n2102), .QN(n37290) );
  DFFRX1 u_decode_u_regfile_reg_r27_q_reg_5_ ( .D(u_decode_u_regfile_N1067), 
        .CK(n37863), .RN(n44145), .Q(n2103) );
  DFFRX1 u_decode_u_regfile_reg_r28_q_reg_5_ ( .D(u_decode_u_regfile_N1104), 
        .CK(n37862), .RN(n44144), .Q(n2104), .QN(n37117) );
  DFFRX1 u_decode_u_regfile_reg_r29_q_reg_5_ ( .D(u_decode_u_regfile_N1141), 
        .CK(n37861), .RN(n44144), .Q(n2105) );
  DFFRX1 u_decode_u_regfile_reg_r30_q_reg_5_ ( .D(u_decode_u_regfile_N1178), 
        .CK(n37860), .RN(n44144), .Q(n2106), .QN(n37110) );
  DFFRX1 u_decode_u_regfile_reg_r31_q_reg_5_ ( .D(u_decode_u_regfile_N1215), 
        .CK(n37859), .RN(n44143), .QN(n37112) );
  DFFRX1 u_decode_u_regfile_reg_r2_q_reg_5_ ( .D(u_decode_u_regfile_N142), 
        .CK(n37858), .RN(n44143), .Q(n2108) );
  DFFRX1 u_decode_u_regfile_reg_r3_q_reg_5_ ( .D(u_decode_u_regfile_N179), 
        .CK(n37857), .RN(n44145), .Q(n2109), .QN(n37283) );
  DFFRX1 u_decode_u_regfile_reg_r4_q_reg_5_ ( .D(u_decode_u_regfile_N216), 
        .CK(n37856), .RN(n44143), .Q(n2110) );
  DFFRX1 u_decode_u_regfile_reg_r5_q_reg_5_ ( .D(u_decode_u_regfile_N253), 
        .CK(n37840), .RN(n44144), .Q(n2111) );
  DFFRX1 u_decode_u_regfile_reg_r6_q_reg_5_ ( .D(u_decode_u_regfile_N290), 
        .CK(n37855), .RN(n44144), .Q(n2112) );
  DFFRX1 u_decode_u_regfile_reg_r7_q_reg_5_ ( .D(u_decode_u_regfile_N327), 
        .CK(n37854), .RN(n44143), .Q(n2113), .QN(n37116) );
  DFFRX1 u_decode_u_regfile_reg_r8_q_reg_5_ ( .D(u_decode_u_regfile_N364), 
        .CK(n37839), .RN(n44145), .Q(n2114), .QN(n37282) );
  DFFRX1 u_decode_u_regfile_reg_r9_q_reg_5_ ( .D(u_decode_u_regfile_N401), 
        .CK(n37853), .RN(n44144), .Q(n2115), .QN(n37286) );
  DFFRX1 u_decode_u_regfile_reg_r10_q_reg_5_ ( .D(u_decode_u_regfile_N438), 
        .CK(n37852), .RN(n44144), .Q(n2116) );
  DFFRX1 u_decode_u_regfile_reg_r11_q_reg_5_ ( .D(u_decode_u_regfile_N475), 
        .CK(n37851), .RN(n44145), .Q(n2117), .QN(n37285) );
  DFFRX1 u_decode_u_regfile_reg_r12_q_reg_5_ ( .D(u_decode_u_regfile_N512), 
        .CK(n37850), .RN(n44144), .Q(n2118) );
  DFFRX1 u_decode_u_regfile_reg_r13_q_reg_5_ ( .D(u_decode_u_regfile_N549), 
        .CK(n37849), .RN(n44144), .Q(n2119) );
  DFFRX1 u_decode_u_regfile_reg_r14_q_reg_5_ ( .D(u_decode_u_regfile_N586), 
        .CK(n37848), .RN(n44144), .Q(n2120) );
  DFFRX1 u_decode_u_regfile_reg_r15_q_reg_5_ ( .D(u_decode_u_regfile_N623), 
        .CK(n37847), .RN(n44144), .Q(n2121) );
  DFFRX1 u_decode_u_regfile_reg_r16_q_reg_5_ ( .D(u_decode_u_regfile_N660), 
        .CK(n37846), .RN(n44144), .Q(n2122), .QN(n37284) );
  DFFRX1 u_decode_u_regfile_reg_r17_q_reg_5_ ( .D(u_decode_u_regfile_N697), 
        .CK(n37845), .RN(n44145), .Q(n2123), .QN(n37287) );
  DFFRX1 u_decode_u_regfile_reg_r18_q_reg_5_ ( .D(u_decode_u_regfile_N734), 
        .CK(n37844), .RN(n44144), .Q(n2124), .QN(n37097) );
  DFFRX1 u_decode_u_regfile_reg_r19_q_reg_5_ ( .D(u_decode_u_regfile_N771), 
        .CK(n37843), .RN(n44145), .Q(n2125), .QN(n37279) );
  DFFRX1 u_decode_u_regfile_reg_r20_q_reg_5_ ( .D(u_decode_u_regfile_N808), 
        .CK(n37842), .RN(n44144), .Q(n2126), .QN(n37113) );
  DFFRX1 u_decode_u_regfile_reg_r21_q_reg_5_ ( .D(u_decode_u_regfile_N845), 
        .CK(n37838), .RN(n44144), .Q(n2127), .QN(n37115) );
  DFFRX1 u_decode_u_regfile_reg_r22_q_reg_5_ ( .D(u_decode_u_regfile_N882), 
        .CK(n37841), .RN(n44144), .Q(n2128), .QN(n37109) );
  DFFRX1 u_decode_u_regfile_reg_r23_q_reg_5_ ( .D(u_decode_u_regfile_N919), 
        .CK(n37877), .RN(n44144), .Q(n2129) );
  DFFRX1 u_csr_branch_target_q_reg_6_ ( .D(u_csr_N3671), .CK(clk_i), .RN(
        n44118), .Q(n54703) );
  DFFRX1 u_fetch_branch_pc_q_reg_6_ ( .D(net2287), .CK(n37867), .RN(n44119), 
        .QN(n2130) );
  DFFRX1 u_csr_pc_m_q_reg_6_ ( .D(opcode_pc_w[6]), .CK(net1867), .RN(n44118), 
        .QN(n37766) );
  DFFRX1 u_csr_branch_target_q_reg_7_ ( .D(u_csr_N3672), .CK(clk_i), .RN(
        n44119), .Q(n54762) );
  DFFRX1 u_fetch_branch_pc_q_reg_7_ ( .D(net2288), .CK(n37867), .RN(n44119), 
        .QN(n2133) );
  DFFRX1 u_csr_pc_m_q_reg_7_ ( .D(opcode_pc_w[7]), .CK(net1867), .RN(n44119), 
        .QN(n37767) );
  DFFRX1 u_csr_branch_target_q_reg_8_ ( .D(u_csr_N3673), .CK(clk_i), .RN(
        n44103), .Q(n54875) );
  DFFRX1 u_fetch_branch_pc_q_reg_8_ ( .D(net2289), .CK(n37867), .RN(n44103), 
        .QN(n2136) );
  DFFRX1 u_csr_pc_m_q_reg_8_ ( .D(opcode_pc_w[8]), .CK(net1867), .RN(n44103), 
        .Q(n2138) );
  DFFRX1 u_csr_branch_target_q_reg_9_ ( .D(u_csr_N3674), .CK(clk_i), .RN(
        n44103), .Q(n54882) );
  DFFRX1 u_fetch_branch_pc_q_reg_9_ ( .D(net2290), .CK(n37867), .RN(n44103), 
        .QN(n2139) );
  DFFRX1 u_csr_pc_m_q_reg_9_ ( .D(opcode_pc_w[9]), .CK(net1867), .RN(n44103), 
        .QN(n37768) );
  DFFRX1 u_csr_branch_target_q_reg_10_ ( .D(u_csr_N3675), .CK(clk_i), .RN(
        n44104), .Q(n54951) );
  DFFRX1 u_fetch_branch_pc_q_reg_10_ ( .D(net2291), .CK(n37867), .RN(n44104), 
        .QN(n2142) );
  DFFRX1 u_csr_pc_m_q_reg_10_ ( .D(opcode_pc_w[10]), .CK(net1867), .RN(n44104), 
        .Q(n2144) );
  DFFRX1 u_csr_branch_target_q_reg_12_ ( .D(u_csr_N3677), .CK(clk_i), .RN(
        n44105), .Q(n55084) );
  DFFRX1 u_fetch_branch_pc_q_reg_12_ ( .D(net2293), .CK(n37867), .RN(n44105), 
        .QN(n2145) );
  DFFRX1 u_csr_pc_m_q_reg_12_ ( .D(opcode_pc_w[12]), .CK(net1872), .RN(n44105), 
        .Q(n2147) );
  DFFRX1 u_csr_branch_target_q_reg_13_ ( .D(u_csr_N3678), .CK(clk_i), .RN(
        n44106), .Q(n55133) );
  DFFRX1 u_fetch_branch_pc_q_reg_13_ ( .D(net2294), .CK(n37867), .RN(n44106), 
        .QN(n2148) );
  DFFRX1 u_csr_pc_m_q_reg_13_ ( .D(opcode_pc_w[13]), .CK(net1872), .RN(n44105), 
        .Q(n2150) );
  DFFRX1 u_csr_branch_target_q_reg_14_ ( .D(u_csr_N3679), .CK(clk_i), .RN(
        n44106), .Q(n55188) );
  DFFRX1 u_fetch_branch_pc_q_reg_14_ ( .D(net2295), .CK(n37867), .RN(n44106), 
        .QN(n2151) );
  DFFRX1 u_csr_pc_m_q_reg_14_ ( .D(opcode_pc_w[14]), .CK(net1872), .RN(n44106), 
        .Q(n2153) );
  DFFRX1 u_mmu_itlb_va_addr_q_reg_14_ ( .D(u_mmu_virt_addr_q[14]), .CK(n37871), 
        .RN(n44186), .QN(n17100) );
  DFFRX1 u_mmu_dtlb_va_addr_q_reg_14_ ( .D(u_mmu_virt_addr_q[14]), .CK(n37872), 
        .RN(n44206), .Q(u_mmu_dtlb_va_addr_q[14]) );
  DFFRX1 u_mmu_itlb_entry_q_reg_14_ ( .D(u_mmu_pte_entry_q[14]), .CK(net1792), 
        .RN(n44171), .Q(u_mmu_itlb_entry_q[14]) );
  DFFRX1 u_mmu_dtlb_entry_q_reg_14_ ( .D(u_mmu_pte_entry_q[14]), .CK(net1782), 
        .RN(n44211), .QN(n2154) );
  DFFRX1 u_csr_branch_target_q_reg_15_ ( .D(u_csr_N3680), .CK(clk_i), .RN(
        n44107), .Q(n55248) );
  DFFRX1 u_fetch_branch_pc_q_reg_15_ ( .D(net2296), .CK(n37867), .RN(n44107), 
        .QN(n2155) );
  DFFRX1 u_mmu_itlb_va_addr_q_reg_15_ ( .D(u_mmu_virt_addr_q[15]), .CK(n37871), 
        .RN(n44186), .Q(n2157) );
  DFFRX1 u_mmu_dtlb_va_addr_q_reg_15_ ( .D(u_mmu_virt_addr_q[15]), .CK(n37872), 
        .RN(n44206), .Q(u_mmu_dtlb_va_addr_q[15]) );
  DFFRX1 u_mmu_itlb_entry_q_reg_15_ ( .D(u_mmu_pte_entry_q[15]), .CK(net1792), 
        .RN(n44171), .Q(u_mmu_itlb_entry_q[15]) );
  DFFRX1 u_mmu_dtlb_entry_q_reg_15_ ( .D(u_mmu_pte_entry_q[15]), .CK(net1782), 
        .RN(n44211), .QN(n2158) );
  DFFRX1 u_csr_branch_target_q_reg_16_ ( .D(u_csr_N3681), .CK(clk_i), .RN(
        n44107), .Q(n55301) );
  DFFRX1 u_fetch_branch_pc_q_reg_16_ ( .D(net2302), .CK(n37866), .RN(n44107), 
        .QN(n2159) );
  DFFRX1 u_csr_pc_m_q_reg_16_ ( .D(opcode_pc_w[16]), .CK(net1872), .RN(n44107), 
        .Q(n2161) );
  DFFRX1 u_csr_branch_target_q_reg_17_ ( .D(u_csr_N3682), .CK(clk_i), .RN(
        n44108), .Q(n55361) );
  DFFRX1 u_fetch_branch_pc_q_reg_17_ ( .D(net2303), .CK(n37866), .RN(n44108), 
        .QN(n2162) );
  DFFRX1 u_csr_pc_m_q_reg_17_ ( .D(opcode_pc_w[17]), .CK(net1872), .RN(n44108), 
        .Q(n2164) );
  DFFRX1 u_csr_branch_target_q_reg_18_ ( .D(u_csr_N3683), .CK(clk_i), .RN(
        n44108), .Q(n55413) );
  DFFRX1 u_fetch_branch_pc_q_reg_18_ ( .D(net2304), .CK(n37866), .RN(n44108), 
        .QN(n2165) );
  DFFRX1 u_csr_pc_m_q_reg_18_ ( .D(opcode_pc_w[18]), .CK(net1872), .RN(n44108), 
        .Q(n2167) );
  DFFRX1 u_csr_branch_target_q_reg_19_ ( .D(u_csr_N3684), .CK(clk_i), .RN(
        n44109), .Q(n55464) );
  DFFRX1 u_fetch_branch_pc_q_reg_19_ ( .D(net2305), .CK(n37866), .RN(n44109), 
        .QN(n2168) );
  DFFRX1 u_csr_pc_m_q_reg_19_ ( .D(opcode_pc_w[19]), .CK(net1872), .RN(n44109), 
        .Q(n2170) );
  DFFRX1 u_csr_branch_target_q_reg_20_ ( .D(u_csr_N3685), .CK(clk_i), .RN(
        n44109), .Q(n55519) );
  DFFRX1 u_fetch_branch_pc_q_reg_20_ ( .D(net2306), .CK(n37866), .RN(n44109), 
        .QN(n2171) );
  DFFRX1 u_csr_pc_m_q_reg_20_ ( .D(opcode_pc_w[20]), .CK(net1872), .RN(n44109), 
        .Q(n2173) );
  DFFRX1 u_csr_branch_target_q_reg_21_ ( .D(u_csr_N3686), .CK(clk_i), .RN(
        n44110), .Q(n55572) );
  DFFRX1 u_fetch_branch_pc_q_reg_21_ ( .D(net2307), .CK(n37866), .RN(n44110), 
        .QN(n2174) );
  DFFRX1 u_csr_pc_m_q_reg_21_ ( .D(opcode_pc_w[21]), .CK(net1872), .RN(n44110), 
        .Q(n2176) );
  DFFRX1 u_csr_branch_target_q_reg_22_ ( .D(u_csr_N3687), .CK(clk_i), .RN(
        n44110), .Q(n55620) );
  DFFRX1 u_fetch_branch_pc_q_reg_22_ ( .D(net2308), .CK(n37866), .RN(n44110), 
        .QN(n2177) );
  DFFRX1 u_csr_pc_m_q_reg_22_ ( .D(opcode_pc_w[22]), .CK(net1872), .RN(n44110), 
        .QN(n37770) );
  DFFRX1 u_csr_branch_target_q_reg_23_ ( .D(u_csr_N3688), .CK(clk_i), .RN(
        n44111), .Q(n55667) );
  DFFRX1 u_fetch_branch_pc_q_reg_23_ ( .D(net2309), .CK(n37866), .RN(n44111), 
        .QN(n2180) );
  DFFRX1 u_csr_pc_m_q_reg_23_ ( .D(opcode_pc_w[23]), .CK(net1872), .RN(n44111), 
        .QN(n37771) );
  DFFRX1 u_csr_branch_target_q_reg_24_ ( .D(u_csr_N3689), .CK(clk_i), .RN(
        n44192), .Q(n55718) );
  DFFRX1 u_fetch_branch_pc_q_reg_24_ ( .D(net2310), .CK(n37866), .RN(n44188), 
        .QN(n2183) );
  DFFRX1 u_csr_pc_m_q_reg_24_ ( .D(opcode_pc_w[24]), .CK(net1872), .RN(n44111), 
        .QN(n37772) );
  DFFRX1 u_csr_branch_target_q_reg_25_ ( .D(u_csr_N3690), .CK(clk_i), .RN(
        n44188), .Q(n55766) );
  DFFRX1 u_csr_pc_m_q_reg_25_ ( .D(opcode_pc_w[25]), .CK(net1872), .RN(n44188), 
        .QN(n37773) );
  DFFRX1 u_csr_branch_target_q_reg_26_ ( .D(u_csr_N3691), .CK(clk_i), .RN(
        n44189), .Q(n55812) );
  DFFRX1 u_csr_pc_m_q_reg_26_ ( .D(opcode_pc_w[26]), .CK(net1872), .RN(n44188), 
        .QN(n37774) );
  DFFRX1 u_csr_pc_m_q_reg_27_ ( .D(n8502), .CK(clk_i), .RN(n44191), .Q(
        u_csr_pc_m_q[27]), .QN(n37757) );
  DFFRX1 u_csr_pc_m_q_reg_28_ ( .D(n8501), .CK(clk_i), .RN(n44193), .Q(
        u_csr_pc_m_q[28]), .QN(n37758) );
  DFFRX1 u_mmu_itlb_va_addr_q_reg_28_ ( .D(n8440), .CK(clk_i), .RN(n44185), 
        .Q(u_mmu_itlb_va_addr_q[28]) );
  DFFRX1 u_mmu_dtlb_va_addr_q_reg_28_ ( .D(n8439), .CK(clk_i), .RN(n44206), 
        .Q(u_mmu_dtlb_va_addr_q[28]) );
  DFFRX1 u_decode_u_regfile_reg_r25_q_reg_28_ ( .D(u_decode_u_regfile_N1016), 
        .CK(n37837), .RN(n44192), .Q(n2192), .QN(n37054) );
  DFFRX1 u_decode_u_regfile_reg_r26_q_reg_28_ ( .D(u_decode_u_regfile_N1053), 
        .CK(n37836), .RN(n44192), .Q(n2193), .QN(n36811) );
  DFFRX1 u_decode_u_regfile_reg_r27_q_reg_28_ ( .D(u_decode_u_regfile_N1090), 
        .CK(n37835), .RN(n44192), .Q(n2194), .QN(n37035) );
  DFFRX1 u_decode_u_regfile_reg_r28_q_reg_28_ ( .D(u_decode_u_regfile_N1127), 
        .CK(n37834), .RN(n44192), .Q(n2195), .QN(n36807) );
  DFFRX1 u_decode_u_regfile_reg_r29_q_reg_28_ ( .D(u_decode_u_regfile_N1164), 
        .CK(n37833), .RN(n44193), .Q(n2196), .QN(n36870) );
  DFFRX1 u_decode_u_regfile_reg_r30_q_reg_28_ ( .D(u_decode_u_regfile_N1201), 
        .CK(n37832), .RN(n44192), .Q(n2197) );
  DFFRX1 u_decode_u_regfile_reg_r31_q_reg_28_ ( .D(u_decode_u_regfile_N1238), 
        .CK(n37831), .RN(n44193), .Q(n2198), .QN(n36808) );
  DFFRX1 u_decode_u_regfile_reg_r1_q_reg_28_ ( .D(u_decode_u_regfile_N128), 
        .CK(n37830), .RN(n44192), .Q(n2199), .QN(n37053) );
  DFFRX1 u_decode_u_regfile_reg_r2_q_reg_28_ ( .D(u_decode_u_regfile_N165), 
        .CK(n37829), .RN(n44191), .Q(n2200), .QN(n36806) );
  DFFRX1 u_decode_u_regfile_reg_r3_q_reg_28_ ( .D(u_decode_u_regfile_N202), 
        .CK(n37828), .RN(n44192), .Q(n2201), .QN(n37044) );
  DFFRX1 u_decode_u_regfile_reg_r4_q_reg_28_ ( .D(u_decode_u_regfile_N239), 
        .CK(n37827), .RN(n44192), .Q(n2202), .QN(n36804) );
  DFFRX1 u_decode_u_regfile_reg_r5_q_reg_28_ ( .D(u_decode_u_regfile_N276), 
        .CK(n37826), .RN(n44193), .Q(n2203), .QN(n40883) );
  DFFRX1 u_decode_u_regfile_reg_r6_q_reg_28_ ( .D(u_decode_u_regfile_N313), 
        .CK(n37825), .RN(n44192), .Q(n2204) );
  DFFRX1 u_decode_u_regfile_reg_r7_q_reg_28_ ( .D(u_decode_u_regfile_N350), 
        .CK(n37824), .RN(n44193), .QN(n36805) );
  DFFRX1 u_decode_u_regfile_reg_r8_q_reg_28_ ( .D(u_decode_u_regfile_N387), 
        .CK(n37823), .RN(n44191), .Q(n2206), .QN(n37042) );
  DFFRX1 u_decode_u_regfile_reg_r9_q_reg_28_ ( .D(u_decode_u_regfile_N424), 
        .CK(n37822), .RN(n44192), .Q(n2207), .QN(n37046) );
  DFFRX1 u_decode_u_regfile_reg_r10_q_reg_28_ ( .D(u_decode_u_regfile_N461), 
        .CK(n37821), .RN(n44191), .Q(n2208), .QN(n36809) );
  DFFRX1 u_decode_u_regfile_reg_r11_q_reg_28_ ( .D(u_decode_u_regfile_N498), 
        .CK(n37820), .RN(n44192), .Q(n2209), .QN(n37043) );
  DFFRX1 u_decode_u_regfile_reg_r12_q_reg_28_ ( .D(u_decode_u_regfile_N535), 
        .CK(n37819), .RN(n44192), .Q(n2210), .QN(n36803) );
  DFFRX1 u_decode_u_regfile_reg_r13_q_reg_28_ ( .D(u_decode_u_regfile_N572), 
        .CK(n37818), .RN(n44193), .Q(n2211), .QN(n36866) );
  DFFRX1 u_decode_u_regfile_reg_r14_q_reg_28_ ( .D(u_decode_u_regfile_N609), 
        .CK(n37817), .RN(n44192), .Q(n2212) );
  DFFRX1 u_decode_u_regfile_reg_r15_q_reg_28_ ( .D(u_decode_u_regfile_N646), 
        .CK(n37816), .RN(n44193), .Q(n2213) );
  DFFRX1 u_decode_u_regfile_reg_r16_q_reg_28_ ( .D(u_decode_u_regfile_N683), 
        .CK(n37815), .RN(n44191), .Q(n2214) );
  DFFRX1 u_decode_u_regfile_reg_r17_q_reg_28_ ( .D(u_decode_u_regfile_N720), 
        .CK(n37814), .RN(n44192), .Q(n2215), .QN(n37057) );
  DFFRX1 u_decode_u_regfile_reg_r18_q_reg_28_ ( .D(u_decode_u_regfile_N757), 
        .CK(n37813), .RN(n44191), .Q(n2216) );
  DFFRX1 u_decode_u_regfile_reg_r19_q_reg_28_ ( .D(u_decode_u_regfile_N794), 
        .CK(n37812), .RN(n44192), .Q(n2217) );
  DFFRX1 u_decode_u_regfile_reg_r20_q_reg_28_ ( .D(u_decode_u_regfile_N831), 
        .CK(n37811), .RN(n44192), .Q(n2218), .QN(n36813) );
  DFFRX1 u_decode_u_regfile_reg_r21_q_reg_28_ ( .D(u_decode_u_regfile_N868), 
        .CK(n37810), .RN(n44193), .Q(n2219) );
  DFFRX1 u_decode_u_regfile_reg_r22_q_reg_28_ ( .D(u_decode_u_regfile_N905), 
        .CK(n37809), .RN(n44192), .Q(n2220) );
  DFFRX1 u_csr_pc_m_q_reg_29_ ( .D(n8500), .CK(clk_i), .RN(n44195), .Q(
        u_csr_pc_m_q[29]), .QN(n37759) );
  DFFRX1 u_csr_branch_target_q_reg_30_ ( .D(u_csr_N3695), .CK(clk_i), .RN(
        n44182), .Q(n56542) );
  DFFRX1 u_decode_u_regfile_reg_r25_q_reg_15_ ( .D(u_decode_u_regfile_N1003), 
        .CK(n37879), .RN(n44124), .Q(n2222), .QN(n37162) );
  DFFRX1 u_decode_u_regfile_reg_r26_q_reg_15_ ( .D(u_decode_u_regfile_N1040), 
        .CK(n37864), .RN(n44124), .Q(n2223) );
  DFFRX1 u_decode_u_regfile_reg_r27_q_reg_15_ ( .D(u_decode_u_regfile_N1077), 
        .CK(n37863), .RN(n44125), .Q(n2224) );
  DFFRX1 u_decode_u_regfile_reg_r28_q_reg_15_ ( .D(u_decode_u_regfile_N1114), 
        .CK(n37862), .RN(n44124), .Q(n2225), .QN(n36895) );
  DFFRX1 u_decode_u_regfile_reg_r1_q_reg_15_ ( .D(u_decode_u_regfile_N115), 
        .CK(n37865), .RN(n44124), .Q(n2226), .QN(n37167) );
  DFFRX1 u_decode_u_regfile_reg_r29_q_reg_15_ ( .D(u_decode_u_regfile_N1151), 
        .CK(n37861), .RN(n44125), .Q(n2227) );
  DFFRX1 u_decode_u_regfile_reg_r30_q_reg_15_ ( .D(u_decode_u_regfile_N1188), 
        .CK(n37860), .RN(n44124), .Q(n2228), .QN(n36882) );
  DFFRX1 u_decode_u_regfile_reg_r31_q_reg_15_ ( .D(u_decode_u_regfile_N1225), 
        .CK(n37859), .RN(n44125), .Q(n2229), .QN(n36883) );
  DFFRX1 u_decode_u_regfile_reg_r2_q_reg_15_ ( .D(u_decode_u_regfile_N152), 
        .CK(n37858), .RN(n44124), .Q(n2230), .QN(n42471) );
  DFFRX1 u_decode_u_regfile_reg_r3_q_reg_15_ ( .D(u_decode_u_regfile_N189), 
        .CK(n37857), .RN(n44125), .Q(n2231), .QN(n37127) );
  DFFRX1 u_decode_u_regfile_reg_r4_q_reg_15_ ( .D(u_decode_u_regfile_N226), 
        .CK(n37856), .RN(n44124), .Q(n2232) );
  DFFRX1 u_decode_u_regfile_reg_r5_q_reg_15_ ( .D(u_decode_u_regfile_N263), 
        .CK(n37840), .RN(n44125), .Q(n2233) );
  DFFRX1 u_decode_u_regfile_reg_r6_q_reg_15_ ( .D(u_decode_u_regfile_N300), 
        .CK(n37855), .RN(n44124), .Q(n2234) );
  DFFRX1 u_decode_u_regfile_reg_r7_q_reg_15_ ( .D(u_decode_u_regfile_N337), 
        .CK(n37854), .RN(n44125), .QN(n36890) );
  DFFRX1 u_decode_u_regfile_reg_r8_q_reg_15_ ( .D(u_decode_u_regfile_N374), 
        .CK(n37839), .RN(n44124), .Q(n2236), .QN(n37153) );
  DFFRX1 u_decode_u_regfile_reg_r9_q_reg_15_ ( .D(u_decode_u_regfile_N411), 
        .CK(n37853), .RN(n44124), .Q(n2237), .QN(n37188) );
  DFFRX1 u_decode_u_regfile_reg_r10_q_reg_15_ ( .D(u_decode_u_regfile_N448), 
        .CK(n37852), .RN(n44124), .Q(n2238) );
  DFFRX1 u_decode_u_regfile_reg_r11_q_reg_15_ ( .D(u_decode_u_regfile_N485), 
        .CK(n37851), .RN(n44125), .Q(n2239), .QN(n37158) );
  DFFRX1 u_decode_u_regfile_reg_r12_q_reg_15_ ( .D(u_decode_u_regfile_N522), 
        .CK(n37850), .RN(n44124), .Q(n2240) );
  DFFRX1 u_decode_u_regfile_reg_r13_q_reg_15_ ( .D(u_decode_u_regfile_N559), 
        .CK(n37849), .RN(n44125), .Q(n2241) );
  DFFRX1 u_decode_u_regfile_reg_r14_q_reg_15_ ( .D(u_decode_u_regfile_N596), 
        .CK(n37848), .RN(n44124), .Q(n2242) );
  DFFRX1 u_decode_u_regfile_reg_r15_q_reg_15_ ( .D(u_decode_u_regfile_N633), 
        .CK(n37847), .RN(n44125), .Q(n2243) );
  DFFRX1 u_decode_u_regfile_reg_r16_q_reg_15_ ( .D(u_decode_u_regfile_N670), 
        .CK(n37846), .RN(n44123), .Q(n2244), .QN(n37157) );
  DFFRX1 u_decode_u_regfile_reg_r17_q_reg_15_ ( .D(u_decode_u_regfile_N707), 
        .CK(n37845), .RN(n44124), .Q(n2245), .QN(n37161) );
  DFFRX1 u_decode_u_regfile_reg_r18_q_reg_15_ ( .D(u_decode_u_regfile_N744), 
        .CK(n37844), .RN(n44124), .Q(n2246), .QN(n36889) );
  DFFRX1 u_decode_u_regfile_reg_r19_q_reg_15_ ( .D(u_decode_u_regfile_N781), 
        .CK(n37843), .RN(n44125), .Q(n2247), .QN(n37122) );
  DFFRX1 u_decode_u_regfile_reg_r20_q_reg_15_ ( .D(u_decode_u_regfile_N818), 
        .CK(n37842), .RN(n44124), .Q(n2248), .QN(n36885) );
  DFFRX1 u_decode_u_regfile_reg_r21_q_reg_15_ ( .D(u_decode_u_regfile_N855), 
        .CK(n37838), .RN(n44125), .Q(n2249), .QN(n36888) );
  DFFRX1 u_decode_u_regfile_reg_r22_q_reg_15_ ( .D(u_decode_u_regfile_N892), 
        .CK(n37841), .RN(n44124), .Q(n2250), .QN(n36878) );
  DFFRX1 u_lsu_mem_addr_q_reg_11_ ( .D(u_lsu_mem_addr_r[11]), .CK(n37869), 
        .RN(n44210), .Q(mmu_lsu_addr_w[11]), .QN(n2251) );
  DFFRX1 u_mmu_lsu_in_addr_q_reg_11_ ( .D(mmu_lsu_addr_w[11]), .CK(n37875), 
        .RN(n44210), .QN(n2252) );
  DFFRX1 u_muldiv_dividend_q_reg_11_ ( .D(u_muldiv_N243), .CK(net1908), .RN(
        n44161), .Q(u_muldiv_dividend_q[11]), .QN(n37439) );
  DFFRX1 u_decode_u_regfile_reg_r26_q_reg_11_ ( .D(u_decode_u_regfile_N1036), 
        .CK(n37864), .RN(n44136), .Q(n2253) );
  DFFRX1 u_decode_u_regfile_reg_r27_q_reg_11_ ( .D(u_decode_u_regfile_N1073), 
        .CK(n37863), .RN(n44137), .Q(n2254) );
  DFFRX1 u_decode_u_regfile_reg_r1_q_reg_11_ ( .D(u_decode_u_regfile_N111), 
        .CK(n37865), .RN(n44137), .Q(n2255), .QN(n37231) );
  DFFRX1 u_decode_u_regfile_reg_r28_q_reg_11_ ( .D(u_decode_u_regfile_N1110), 
        .CK(n37862), .RN(n44137), .Q(n2256), .QN(n36994) );
  DFFRX1 u_decode_u_regfile_reg_r29_q_reg_11_ ( .D(u_decode_u_regfile_N1147), 
        .CK(n37861), .RN(n44137), .Q(n2257) );
  DFFRX1 u_decode_u_regfile_reg_r30_q_reg_11_ ( .D(u_decode_u_regfile_N1184), 
        .CK(n37860), .RN(n44137), .Q(n2258), .QN(n36963) );
  DFFRX1 u_decode_u_regfile_reg_r31_q_reg_11_ ( .D(u_decode_u_regfile_N1221), 
        .CK(n37859), .RN(n44138), .Q(n2259), .QN(n36956) );
  DFFRX1 u_decode_u_regfile_reg_r2_q_reg_11_ ( .D(u_decode_u_regfile_N148), 
        .CK(n37858), .RN(n44136), .Q(n2260) );
  DFFRX1 u_decode_u_regfile_reg_r3_q_reg_11_ ( .D(u_decode_u_regfile_N185), 
        .CK(n37857), .RN(n44137), .Q(n2261), .QN(n37221) );
  DFFRX1 u_decode_u_regfile_reg_r4_q_reg_11_ ( .D(u_decode_u_regfile_N222), 
        .CK(n37856), .RN(n44137), .Q(n2262) );
  DFFRX1 u_decode_u_regfile_reg_r5_q_reg_11_ ( .D(u_decode_u_regfile_N259), 
        .CK(n37840), .RN(n44137), .Q(n2263) );
  DFFRX1 u_decode_u_regfile_reg_r6_q_reg_11_ ( .D(u_decode_u_regfile_N296), 
        .CK(n37855), .RN(n44137), .Q(n2264) );
  DFFRX1 u_decode_u_regfile_reg_r7_q_reg_11_ ( .D(u_decode_u_regfile_N333), 
        .CK(n37854), .RN(n44138), .QN(n36977) );
  DFFRX1 u_decode_u_regfile_reg_r8_q_reg_11_ ( .D(u_decode_u_regfile_N370), 
        .CK(n37839), .RN(n44136), .Q(n2266), .QN(n37223) );
  DFFRX1 u_decode_u_regfile_reg_r9_q_reg_11_ ( .D(u_decode_u_regfile_N407), 
        .CK(n37853), .RN(n44137), .Q(n2267), .QN(n37229) );
  DFFRX1 u_decode_u_regfile_reg_r10_q_reg_11_ ( .D(u_decode_u_regfile_N444), 
        .CK(n37852), .RN(n44136), .Q(n2268) );
  DFFRX1 u_decode_u_regfile_reg_r11_q_reg_11_ ( .D(u_decode_u_regfile_N481), 
        .CK(n37851), .RN(n44137), .Q(n2269), .QN(n37225) );
  DFFRX1 u_decode_u_regfile_reg_r12_q_reg_11_ ( .D(u_decode_u_regfile_N518), 
        .CK(n37850), .RN(n44137), .Q(n2270) );
  DFFRX1 u_decode_u_regfile_reg_r13_q_reg_11_ ( .D(u_decode_u_regfile_N555), 
        .CK(n37849), .RN(n44138), .Q(n2271) );
  DFFRX1 u_decode_u_regfile_reg_r14_q_reg_11_ ( .D(u_decode_u_regfile_N592), 
        .CK(n37848), .RN(n44137), .Q(n2272) );
  DFFRX1 u_decode_u_regfile_reg_r15_q_reg_11_ ( .D(u_decode_u_regfile_N629), 
        .CK(n37847), .RN(n44138), .Q(n2273) );
  DFFRX1 u_decode_u_regfile_reg_r16_q_reg_11_ ( .D(u_decode_u_regfile_N666), 
        .CK(n37846), .RN(n44136), .Q(n2274), .QN(n37230) );
  DFFRX1 u_decode_u_regfile_reg_r17_q_reg_11_ ( .D(u_decode_u_regfile_N703), 
        .CK(n37845), .RN(n44137), .Q(n2275), .QN(n37232) );
  DFFRX1 u_decode_u_regfile_reg_r18_q_reg_11_ ( .D(u_decode_u_regfile_N740), 
        .CK(n37844), .RN(n44136), .Q(n2276), .QN(n36976) );
  DFFRX1 u_decode_u_regfile_reg_r19_q_reg_11_ ( .D(u_decode_u_regfile_N777), 
        .CK(n37843), .RN(n44137), .Q(n2277), .QN(n37224) );
  DFFRX1 u_decode_u_regfile_reg_r20_q_reg_11_ ( .D(u_decode_u_regfile_N814), 
        .CK(n37842), .RN(n44137), .Q(n2278), .QN(n36967) );
  DFFRX1 u_decode_u_regfile_reg_r21_q_reg_11_ ( .D(u_decode_u_regfile_N851), 
        .CK(n37838), .RN(n44138), .Q(n2279), .QN(n36974) );
  DFFRX1 u_decode_u_regfile_reg_r22_q_reg_11_ ( .D(u_decode_u_regfile_N888), 
        .CK(n37841), .RN(n44137), .Q(n2280), .QN(n36943) );
  DFFRX1 u_decode_u_regfile_reg_r23_q_reg_11_ ( .D(u_decode_u_regfile_N925), 
        .CK(n37877), .RN(n44138), .Q(n2281) );
  DFFRX1 u_decode_u_regfile_reg_r24_q_reg_11_ ( .D(u_decode_u_regfile_N962), 
        .CK(n37878), .RN(n44136), .Q(n2282), .QN(n37228) );
  DFFRX1 u_lsu_mem_addr_q_reg_19_ ( .D(u_lsu_mem_addr_r[19]), .CK(n37876), 
        .RN(n44185), .Q(mmu_lsu_addr_w[19]), .QN(n8310) );
  DFFRX1 u_mmu_lsu_in_addr_q_reg_19_ ( .D(mmu_lsu_addr_w[19]), .CK(n37873), 
        .RN(n44185), .QN(n2283) );
  DFFRX1 u_mmu_itlb_va_addr_q_reg_19_ ( .D(u_mmu_virt_addr_q[19]), .CK(n37871), 
        .RN(n44185), .Q(n2284) );
  DFFRX1 u_mmu_dtlb_va_addr_q_reg_19_ ( .D(u_mmu_virt_addr_q[19]), .CK(n37872), 
        .RN(n44207), .Q(u_mmu_dtlb_va_addr_q[19]) );
  DFFRX1 u_mmu_itlb_entry_q_reg_19_ ( .D(u_mmu_pte_entry_q[19]), .CK(net1792), 
        .RN(n44171), .Q(u_mmu_itlb_entry_q[19]) );
  DFFRX1 u_mmu_dtlb_entry_q_reg_19_ ( .D(u_mmu_pte_entry_q[19]), .CK(net1782), 
        .RN(n44196), .QN(n2285) );
  DFFRX1 u_decode_u_regfile_reg_r25_q_reg_19_ ( .D(u_decode_u_regfile_N1007), 
        .CK(n37837), .RN(n44103), .Q(n2286) );
  DFFRX1 u_decode_u_regfile_reg_r26_q_reg_19_ ( .D(u_decode_u_regfile_N1044), 
        .CK(n37836), .RN(n44102), .Q(n2287) );
  DFFRX1 u_decode_u_regfile_reg_r27_q_reg_19_ ( .D(u_decode_u_regfile_N1081), 
        .CK(n37835), .RN(n44087), .Q(n2288) );
  DFFRX1 u_decode_u_regfile_reg_r28_q_reg_19_ ( .D(u_decode_u_regfile_N1118), 
        .CK(n37834), .RN(n44102), .Q(n2289), .QN(n36892) );
  DFFRX1 u_decode_u_regfile_reg_r29_q_reg_19_ ( .D(u_decode_u_regfile_N1155), 
        .CK(n37833), .RN(n44087), .Q(n2290) );
  DFFRX1 u_decode_u_regfile_reg_r1_q_reg_19_ ( .D(u_decode_u_regfile_N119), 
        .CK(n37830), .RN(n44103), .Q(n2291) );
  DFFRX1 u_decode_u_regfile_reg_r30_q_reg_19_ ( .D(u_decode_u_regfile_N1192), 
        .CK(n37832), .RN(n44103), .Q(n2292), .QN(n36894) );
  DFFRX1 u_decode_u_regfile_reg_r31_q_reg_19_ ( .D(u_decode_u_regfile_N1229), 
        .CK(n37831), .RN(n44087), .Q(n2293), .QN(n36881) );
  DFFRX1 u_decode_u_regfile_reg_r2_q_reg_19_ ( .D(u_decode_u_regfile_N156), 
        .CK(n37829), .RN(n44102), .Q(n2294) );
  DFFRX1 u_decode_u_regfile_reg_r3_q_reg_19_ ( .D(u_decode_u_regfile_N193), 
        .CK(n37828), .RN(n44087), .Q(n2295) );
  DFFRX1 u_decode_u_regfile_reg_r4_q_reg_19_ ( .D(u_decode_u_regfile_N230), 
        .CK(n37827), .RN(n44102), .Q(n2296) );
  DFFRX1 u_decode_u_regfile_reg_r5_q_reg_19_ ( .D(u_decode_u_regfile_N267), 
        .CK(n37826), .RN(n44087), .Q(n2297), .QN(n42527) );
  DFFRX1 u_decode_u_regfile_reg_r6_q_reg_19_ ( .D(u_decode_u_regfile_N304), 
        .CK(n37825), .RN(n44103), .Q(n2298), .QN(n42526) );
  DFFRX1 u_decode_u_regfile_reg_r7_q_reg_19_ ( .D(u_decode_u_regfile_N341), 
        .CK(n37824), .RN(n44087), .QN(n36887) );
  DFFRX1 u_decode_u_regfile_reg_r8_q_reg_19_ ( .D(u_decode_u_regfile_N378), 
        .CK(n37823), .RN(n44102), .Q(n2300) );
  DFFRX1 u_decode_u_regfile_reg_r9_q_reg_19_ ( .D(u_decode_u_regfile_N415), 
        .CK(n37822), .RN(n44103), .Q(n2301) );
  DFFRX1 u_decode_u_regfile_reg_r10_q_reg_19_ ( .D(u_decode_u_regfile_N452), 
        .CK(n37821), .RN(n44102), .Q(n2302) );
  DFFRX1 u_decode_u_regfile_reg_r11_q_reg_19_ ( .D(u_decode_u_regfile_N489), 
        .CK(n37820), .RN(n44087), .Q(n2303), .QN(n42474) );
  DFFRX1 u_decode_u_regfile_reg_r12_q_reg_19_ ( .D(u_decode_u_regfile_N526), 
        .CK(n37819), .RN(n44102), .Q(n2304) );
  DFFRX1 u_decode_u_regfile_reg_r13_q_reg_19_ ( .D(u_decode_u_regfile_N563), 
        .CK(n37818), .RN(n44087), .Q(n2305) );
  DFFRX1 u_decode_u_regfile_reg_r14_q_reg_19_ ( .D(u_decode_u_regfile_N600), 
        .CK(n37817), .RN(n44103), .Q(n2306) );
  DFFRX1 u_decode_u_regfile_reg_r15_q_reg_19_ ( .D(u_decode_u_regfile_N637), 
        .CK(n37816), .RN(n44088), .Q(n2307) );
  DFFRX1 u_decode_u_regfile_reg_r16_q_reg_19_ ( .D(u_decode_u_regfile_N674), 
        .CK(n37815), .RN(n44102), .Q(n2308) );
  DFFRX1 u_decode_u_regfile_reg_r17_q_reg_19_ ( .D(u_decode_u_regfile_N711), 
        .CK(n37814), .RN(n44103), .Q(n2309) );
  DFFRX1 u_decode_u_regfile_reg_r18_q_reg_19_ ( .D(u_decode_u_regfile_N748), 
        .CK(n37813), .RN(n44102), .Q(n2310), .QN(n36884) );
  DFFRX1 u_decode_u_regfile_reg_r19_q_reg_19_ ( .D(u_decode_u_regfile_N785), 
        .CK(n37812), .RN(n44091), .Q(n2311) );
  DFFRX1 u_decode_u_regfile_reg_r20_q_reg_19_ ( .D(u_decode_u_regfile_N822), 
        .CK(n37811), .RN(n44102), .Q(n2312), .QN(n36891) );
  DFFRX1 u_decode_u_regfile_reg_r21_q_reg_19_ ( .D(u_decode_u_regfile_N859), 
        .CK(n37810), .RN(n44087), .Q(n2313), .QN(n36896) );
  DFFRX1 u_decode_u_regfile_reg_r22_q_reg_19_ ( .D(u_decode_u_regfile_N896), 
        .CK(n37809), .RN(n44102), .Q(n2314), .QN(n36886) );
  DFFRX1 u_decode_u_regfile_reg_r23_q_reg_19_ ( .D(u_decode_u_regfile_N933), 
        .CK(n37880), .RN(n44087), .Q(n2315) );
  DFFRX1 u_lsu_mem_addr_q_reg_6_ ( .D(u_lsu_mem_addr_r[6]), .CK(n37869), .RN(
        n44199), .Q(mmu_lsu_addr_w[6]), .QN(n2316) );
  DFFRX1 u_mmu_lsu_in_addr_q_reg_6_ ( .D(mmu_lsu_addr_w[6]), .CK(n37875), .RN(
        n44199), .QN(n2317) );
  DFFRX1 u_muldiv_dividend_q_reg_6_ ( .D(u_muldiv_N238), .CK(net1908), .RN(
        n44161), .Q(u_muldiv_dividend_q[6]), .QN(n37423) );
  DFFRX1 u_decode_u_regfile_reg_r26_q_reg_6_ ( .D(u_decode_u_regfile_N1031), 
        .CK(n37864), .RN(n44142), .Q(n2318) );
  DFFRX1 u_decode_u_regfile_reg_r1_q_reg_6_ ( .D(u_decode_u_regfile_N106), 
        .CK(n37865), .RN(n44143), .Q(n2319), .QN(n37281) );
  DFFRX1 u_decode_u_regfile_reg_r27_q_reg_6_ ( .D(u_decode_u_regfile_N1068), 
        .CK(n37863), .RN(n44143), .Q(n2320) );
  DFFRX1 u_decode_u_regfile_reg_r28_q_reg_6_ ( .D(u_decode_u_regfile_N1105), 
        .CK(n37862), .RN(n44142), .Q(n2321), .QN(n37106) );
  DFFRX1 u_decode_u_regfile_reg_r29_q_reg_6_ ( .D(u_decode_u_regfile_N1142), 
        .CK(n37861), .RN(n44142), .Q(n2322) );
  DFFRX1 u_decode_u_regfile_reg_r30_q_reg_6_ ( .D(u_decode_u_regfile_N1179), 
        .CK(n37860), .RN(n44142), .Q(n2323), .QN(n37101) );
  DFFRX1 u_decode_u_regfile_reg_r31_q_reg_6_ ( .D(u_decode_u_regfile_N1216), 
        .CK(n37859), .RN(n44141), .Q(n2324), .QN(n37100) );
  DFFRX1 u_decode_u_regfile_reg_r2_q_reg_6_ ( .D(u_decode_u_regfile_N143), 
        .CK(n37858), .RN(n44142), .Q(n2325) );
  DFFRX1 u_decode_u_regfile_reg_r3_q_reg_6_ ( .D(u_decode_u_regfile_N180), 
        .CK(n37857), .RN(n44143), .Q(n2326), .QN(n37272) );
  DFFRX1 u_decode_u_regfile_reg_r4_q_reg_6_ ( .D(u_decode_u_regfile_N217), 
        .CK(n37856), .RN(n44142), .Q(n2327) );
  DFFRX1 u_decode_u_regfile_reg_r5_q_reg_6_ ( .D(u_decode_u_regfile_N254), 
        .CK(n37840), .RN(n44142), .Q(n2328) );
  DFFRX1 u_decode_u_regfile_reg_r6_q_reg_6_ ( .D(u_decode_u_regfile_N291), 
        .CK(n37855), .RN(n44142), .Q(n2329) );
  DFFRX1 u_decode_u_regfile_reg_r7_q_reg_6_ ( .D(u_decode_u_regfile_N328), 
        .CK(n37854), .RN(n44142), .QN(n37104) );
  DFFRX1 u_decode_u_regfile_reg_r8_q_reg_6_ ( .D(u_decode_u_regfile_N365), 
        .CK(n37839), .RN(n44143), .Q(n2331), .QN(n37273) );
  DFFRX1 u_decode_u_regfile_reg_r9_q_reg_6_ ( .D(u_decode_u_regfile_N402), 
        .CK(n37853), .RN(n44143), .Q(n2332), .QN(n37275) );
  DFFRX1 u_decode_u_regfile_reg_r10_q_reg_6_ ( .D(u_decode_u_regfile_N439), 
        .CK(n37852), .RN(n44142), .Q(n2333) );
  DFFRX1 u_decode_u_regfile_reg_r11_q_reg_6_ ( .D(u_decode_u_regfile_N476), 
        .CK(n37851), .RN(n44143), .Q(n2334), .QN(n37276) );
  DFFRX1 u_decode_u_regfile_reg_r12_q_reg_6_ ( .D(u_decode_u_regfile_N513), 
        .CK(n37850), .RN(n44143), .Q(n2335) );
  DFFRX1 u_decode_u_regfile_reg_r13_q_reg_6_ ( .D(u_decode_u_regfile_N550), 
        .CK(n37849), .RN(n44142), .Q(n2336) );
  DFFRX1 u_decode_u_regfile_reg_r14_q_reg_6_ ( .D(u_decode_u_regfile_N587), 
        .CK(n37848), .RN(n44142), .Q(n2337) );
  DFFRX1 u_decode_u_regfile_reg_r15_q_reg_6_ ( .D(u_decode_u_regfile_N624), 
        .CK(n37847), .RN(n44142), .Q(n2338) );
  DFFRX1 u_decode_u_regfile_reg_r16_q_reg_6_ ( .D(u_decode_u_regfile_N661), 
        .CK(n37846), .RN(n44143), .Q(n2339), .QN(n37274) );
  DFFRX1 u_decode_u_regfile_reg_r17_q_reg_6_ ( .D(u_decode_u_regfile_N698), 
        .CK(n37845), .RN(n44143), .Q(n2340), .QN(n37277) );
  DFFRX1 u_decode_u_regfile_reg_r18_q_reg_6_ ( .D(u_decode_u_regfile_N735), 
        .CK(n37844), .RN(n44142), .Q(n2341), .QN(n37105) );
  DFFRX1 u_decode_u_regfile_reg_r19_q_reg_6_ ( .D(u_decode_u_regfile_N772), 
        .CK(n37843), .RN(n44143), .Q(n2342), .QN(n37271) );
  DFFRX1 u_decode_u_regfile_reg_r20_q_reg_6_ ( .D(u_decode_u_regfile_N809), 
        .CK(n37842), .RN(n44142), .Q(n2343), .QN(n37102) );
  DFFRX1 u_decode_u_regfile_reg_r21_q_reg_6_ ( .D(u_decode_u_regfile_N846), 
        .CK(n37838), .RN(n44142), .Q(n2344), .QN(n37103) );
  DFFRX1 u_decode_u_regfile_reg_r22_q_reg_6_ ( .D(u_decode_u_regfile_N883), 
        .CK(n37841), .RN(n44142), .Q(n2345), .QN(n37099) );
  DFFRX1 u_decode_u_regfile_reg_r23_q_reg_6_ ( .D(u_decode_u_regfile_N920), 
        .CK(n37877), .RN(n44142), .Q(n2346) );
  DFFRX1 u_decode_u_regfile_reg_r24_q_reg_6_ ( .D(u_decode_u_regfile_N957), 
        .CK(n37878), .RN(n44143), .Q(n2347), .QN(n37280) );
  DFFRX1 u_lsu_mem_data_wr_q_reg_6_ ( .D(u_lsu_N200), .CK(n37874), .RN(n44200), 
        .QN(n2348) );
  DFFRX1 u_lsu_mem_data_wr_q_reg_2_ ( .D(u_lsu_N196), .CK(n37874), .RN(n44200), 
        .QN(n2349) );
  DFFRX1 u_lsu_mem_addr_q_reg_10_ ( .D(u_lsu_mem_addr_r[10]), .CK(n37869), 
        .RN(n44210), .Q(mmu_lsu_addr_w[10]), .QN(n2350) );
  DFFRX1 u_mmu_lsu_in_addr_q_reg_10_ ( .D(mmu_lsu_addr_w[10]), .CK(n37875), 
        .RN(n44210), .QN(n2351) );
  DFFRX1 u_muldiv_dividend_q_reg_10_ ( .D(u_muldiv_N242), .CK(net1908), .RN(
        n44161), .Q(u_muldiv_dividend_q[10]), .QN(n37437) );
  DFFRX1 u_decode_u_regfile_reg_r26_q_reg_10_ ( .D(u_decode_u_regfile_N1035), 
        .CK(n37864), .RN(n44135), .Q(n2352), .QN(n42512) );
  DFFRX1 u_decode_u_regfile_reg_r27_q_reg_10_ ( .D(u_decode_u_regfile_N1072), 
        .CK(n37863), .RN(n44135), .Q(n2353) );
  DFFRX1 u_decode_u_regfile_reg_r1_q_reg_10_ ( .D(u_decode_u_regfile_N110), 
        .CK(n37865), .RN(n44135), .Q(n2354), .QN(n37265) );
  DFFRX1 u_decode_u_regfile_reg_r28_q_reg_10_ ( .D(u_decode_u_regfile_N1109), 
        .CK(n37862), .RN(n44135), .Q(n2355), .QN(n37089) );
  DFFRX1 u_decode_u_regfile_reg_r29_q_reg_10_ ( .D(u_decode_u_regfile_N1146), 
        .CK(n37861), .RN(n44136), .Q(n2356) );
  DFFRX1 u_decode_u_regfile_reg_r30_q_reg_10_ ( .D(u_decode_u_regfile_N1183), 
        .CK(n37860), .RN(n44135), .Q(n2357), .QN(n37077) );
  DFFRX1 u_decode_u_regfile_reg_r31_q_reg_10_ ( .D(u_decode_u_regfile_N1220), 
        .CK(n37859), .RN(n44136), .Q(n2358), .QN(n37078) );
  DFFRX1 u_decode_u_regfile_reg_r2_q_reg_10_ ( .D(u_decode_u_regfile_N147), 
        .CK(n37858), .RN(n44135), .Q(n2359) );
  DFFRX1 u_decode_u_regfile_reg_r3_q_reg_10_ ( .D(u_decode_u_regfile_N184), 
        .CK(n37857), .RN(n44135), .Q(n2360), .QN(n37253) );
  DFFRX1 u_decode_u_regfile_reg_r4_q_reg_10_ ( .D(u_decode_u_regfile_N221), 
        .CK(n37856), .RN(n44135), .Q(n2361) );
  DFFRX1 u_decode_u_regfile_reg_r5_q_reg_10_ ( .D(u_decode_u_regfile_N258), 
        .CK(n37840), .RN(n44136), .Q(n2362) );
  DFFRX1 u_decode_u_regfile_reg_r6_q_reg_10_ ( .D(u_decode_u_regfile_N295), 
        .CK(n37855), .RN(n44135), .Q(n2363) );
  DFFRX1 u_decode_u_regfile_reg_r7_q_reg_10_ ( .D(u_decode_u_regfile_N332), 
        .CK(n37854), .RN(n44136), .QN(n37085) );
  DFFRX1 u_decode_u_regfile_reg_r8_q_reg_10_ ( .D(u_decode_u_regfile_N369), 
        .CK(n37839), .RN(n44134), .Q(n2365), .QN(n37254) );
  DFFRX1 u_decode_u_regfile_reg_r9_q_reg_10_ ( .D(u_decode_u_regfile_N406), 
        .CK(n37853), .RN(n44135), .Q(n2366), .QN(n37256) );
  DFFRX1 u_decode_u_regfile_reg_r10_q_reg_10_ ( .D(u_decode_u_regfile_N443), 
        .CK(n37852), .RN(n44134), .Q(n2367) );
  DFFRX1 u_decode_u_regfile_reg_r11_q_reg_10_ ( .D(u_decode_u_regfile_N480), 
        .CK(n37851), .RN(n44136), .Q(n2368), .QN(n37255) );
  DFFRX1 u_decode_u_regfile_reg_r12_q_reg_10_ ( .D(u_decode_u_regfile_N517), 
        .CK(n37850), .RN(n44135), .Q(n2369) );
  DFFRX1 u_decode_u_regfile_reg_r13_q_reg_10_ ( .D(u_decode_u_regfile_N554), 
        .CK(n37849), .RN(n44136), .Q(n2370) );
  DFFRX1 u_decode_u_regfile_reg_r14_q_reg_10_ ( .D(u_decode_u_regfile_N591), 
        .CK(n37848), .RN(n44135), .Q(n2371) );
  DFFRX1 u_decode_u_regfile_reg_r15_q_reg_10_ ( .D(u_decode_u_regfile_N628), 
        .CK(n37847), .RN(n44136), .Q(n2372) );
  DFFRX1 u_decode_u_regfile_reg_r16_q_reg_10_ ( .D(u_decode_u_regfile_N665), 
        .CK(n37846), .RN(n44134), .Q(n2373), .QN(n37257) );
  DFFRX1 u_decode_u_regfile_reg_r17_q_reg_10_ ( .D(u_decode_u_regfile_N702), 
        .CK(n37845), .RN(n44135), .Q(n2374), .QN(n37261) );
  DFFRX1 u_decode_u_regfile_reg_r18_q_reg_10_ ( .D(u_decode_u_regfile_N739), 
        .CK(n37844), .RN(n44135), .Q(n2375), .QN(n37084) );
  DFFRX1 u_decode_u_regfile_reg_r19_q_reg_10_ ( .D(u_decode_u_regfile_N776), 
        .CK(n37843), .RN(n44135), .Q(n2376), .QN(n37251) );
  DFFRX1 u_decode_u_regfile_reg_r20_q_reg_10_ ( .D(u_decode_u_regfile_N813), 
        .CK(n37842), .RN(n44135), .Q(n2377), .QN(n37079) );
  DFFRX1 u_decode_u_regfile_reg_r21_q_reg_10_ ( .D(u_decode_u_regfile_N850), 
        .CK(n37838), .RN(n44136), .Q(n2378), .QN(n37081) );
  DFFRX1 u_decode_u_regfile_reg_r22_q_reg_10_ ( .D(u_decode_u_regfile_N887), 
        .CK(n37841), .RN(n44135), .Q(n2379), .QN(n37075) );
  DFFRX1 u_decode_u_regfile_reg_r23_q_reg_10_ ( .D(u_decode_u_regfile_N924), 
        .CK(n37877), .RN(n44136), .Q(n2380) );
  DFFRX1 u_decode_u_regfile_reg_r24_q_reg_10_ ( .D(u_decode_u_regfile_N961), 
        .CK(n37878), .RN(n44134), .Q(n2381), .QN(n37262) );
  DFFRX1 u_lsu_mem_data_wr_q_reg_10_ ( .D(u_lsu_N204), .CK(n37874), .RN(n44161), .QN(n2382) );
  DFFRX1 u_lsu_mem_addr_q_reg_20_ ( .D(u_lsu_mem_addr_r[20]), .CK(n37876), 
        .RN(n44184), .Q(mmu_lsu_addr_w[20]), .QN(n8314) );
  DFFRX1 u_mmu_lsu_in_addr_q_reg_20_ ( .D(mmu_lsu_addr_w[20]), .CK(n37873), 
        .RN(n44184), .QN(n2383) );
  DFFRX1 u_mmu_itlb_va_addr_q_reg_20_ ( .D(u_mmu_virt_addr_q[20]), .CK(n37871), 
        .RN(n44184), .Q(n2384) );
  DFFRX1 u_mmu_dtlb_va_addr_q_reg_20_ ( .D(u_mmu_virt_addr_q[20]), .CK(n37872), 
        .RN(n44207), .Q(u_mmu_dtlb_va_addr_q[20]) );
  DFFRX1 u_mmu_itlb_entry_q_reg_20_ ( .D(u_mmu_pte_entry_q[20]), .CK(net1792), 
        .RN(n44171), .Q(u_mmu_itlb_entry_q[20]) );
  DFFRX1 u_mmu_dtlb_entry_q_reg_20_ ( .D(u_mmu_pte_entry_q[20]), .CK(net1782), 
        .RN(n44197), .QN(n2385) );
  DFFRX1 u_decode_u_regfile_reg_r25_q_reg_20_ ( .D(u_decode_u_regfile_N1008), 
        .CK(n37837), .RN(n44088), .Q(n2386) );
  DFFRX1 u_decode_u_regfile_reg_r26_q_reg_20_ ( .D(u_decode_u_regfile_N1045), 
        .CK(n37836), .RN(n44088), .Q(n2387), .QN(n37061) );
  DFFRX1 u_decode_u_regfile_reg_r27_q_reg_20_ ( .D(u_decode_u_regfile_N1082), 
        .CK(n37835), .RN(n44089), .Q(n2388), .QN(n37118) );
  DFFRX1 u_decode_u_regfile_reg_r28_q_reg_20_ ( .D(u_decode_u_regfile_N1119), 
        .CK(n37834), .RN(n44088), .Q(n2389), .QN(n37041) );
  DFFRX1 u_decode_u_regfile_reg_r29_q_reg_20_ ( .D(u_decode_u_regfile_N1156), 
        .CK(n37833), .RN(n44089), .Q(n2390), .QN(n37073) );
  DFFRX1 u_decode_u_regfile_reg_r30_q_reg_20_ ( .D(u_decode_u_regfile_N1193), 
        .CK(n37832), .RN(n44088), .Q(n2391) );
  DFFRX1 u_decode_u_regfile_reg_r1_q_reg_20_ ( .D(u_decode_u_regfile_N120), 
        .CK(n37830), .RN(n44088), .Q(n2392) );
  DFFRX1 u_decode_u_regfile_reg_r31_q_reg_20_ ( .D(u_decode_u_regfile_N1230), 
        .CK(n37831), .RN(n44089), .Q(n2393) );
  DFFRX1 u_decode_u_regfile_reg_r2_q_reg_20_ ( .D(u_decode_u_regfile_N157), 
        .CK(n37829), .RN(n44088), .Q(n2394), .QN(n37052) );
  DFFRX1 u_decode_u_regfile_reg_r3_q_reg_20_ ( .D(u_decode_u_regfile_N194), 
        .CK(n37828), .RN(n44089), .Q(n2395), .QN(n37114) );
  DFFRX1 u_decode_u_regfile_reg_r4_q_reg_20_ ( .D(u_decode_u_regfile_N231), 
        .CK(n37827), .RN(n44088), .Q(n2396), .QN(n37070) );
  DFFRX1 u_decode_u_regfile_reg_r5_q_reg_20_ ( .D(u_decode_u_regfile_N268), 
        .CK(n37826), .RN(n44089), .Q(n2397), .QN(n37050) );
  DFFRX1 u_decode_u_regfile_reg_r6_q_reg_20_ ( .D(u_decode_u_regfile_N305), 
        .CK(n37825), .RN(n44088), .Q(n2398) );
  DFFRX1 u_decode_u_regfile_reg_r7_q_reg_20_ ( .D(u_decode_u_regfile_N342), 
        .CK(n37824), .RN(n44089), .Q(n2399), .QN(n37316) );
  DFFRX1 u_decode_u_regfile_reg_r8_q_reg_20_ ( .D(u_decode_u_regfile_N379), 
        .CK(n37823), .RN(n44087), .Q(n2400) );
  DFFRX1 u_decode_u_regfile_reg_r9_q_reg_20_ ( .D(u_decode_u_regfile_N416), 
        .CK(n37822), .RN(n44088), .Q(n2401) );
  DFFRX1 u_decode_u_regfile_reg_r10_q_reg_20_ ( .D(u_decode_u_regfile_N453), 
        .CK(n37821), .RN(n44088), .Q(n2402), .QN(n37062) );
  DFFRX1 u_decode_u_regfile_reg_r11_q_reg_20_ ( .D(u_decode_u_regfile_N490), 
        .CK(n37820), .RN(n44089), .Q(n2403), .QN(n37180) );
  DFFRX1 u_decode_u_regfile_reg_r12_q_reg_20_ ( .D(u_decode_u_regfile_N527), 
        .CK(n37819), .RN(n44088), .Q(n2404), .QN(n37068) );
  DFFRX1 u_decode_u_regfile_reg_r13_q_reg_20_ ( .D(u_decode_u_regfile_N564), 
        .CK(n37818), .RN(n44089), .Q(n2405), .QN(n37069) );
  DFFRX1 u_decode_u_regfile_reg_r14_q_reg_20_ ( .D(u_decode_u_regfile_N601), 
        .CK(n37817), .RN(n44088), .Q(n2406), .QN(n37055) );
  DFFRX1 u_decode_u_regfile_reg_r15_q_reg_20_ ( .D(u_decode_u_regfile_N638), 
        .CK(n37816), .RN(n44089), .Q(n2407), .QN(n37051) );
  DFFRX1 u_decode_u_regfile_reg_r17_q_reg_20_ ( .D(u_decode_u_regfile_N712), 
        .CK(n37814), .RN(n44089), .Q(n2409) );
  DFFRX1 u_decode_u_regfile_reg_r18_q_reg_20_ ( .D(u_decode_u_regfile_N749), 
        .CK(n37813), .RN(n44088), .Q(n2410) );
  DFFRX1 u_decode_u_regfile_reg_r20_q_reg_20_ ( .D(u_decode_u_regfile_N823), 
        .CK(n37811), .RN(n44088), .Q(n2412), .QN(n37060) );
  DFFRX1 u_decode_u_regfile_reg_r21_q_reg_20_ ( .D(u_decode_u_regfile_N860), 
        .CK(n37810), .RN(n44089), .Q(n2413) );
  DFFRX1 u_decode_u_regfile_reg_r22_q_reg_20_ ( .D(u_decode_u_regfile_N897), 
        .CK(n37809), .RN(n44088), .Q(n2414) );
  DFFRX1 u_decode_u_regfile_reg_r23_q_reg_20_ ( .D(u_decode_u_regfile_N934), 
        .CK(n37880), .RN(n44089), .Q(n2415) );
  DFFRX1 u_lsu_mem_data_wr_q_reg_3_ ( .D(u_lsu_N197), .CK(n37874), .RN(n44200), 
        .QN(n2416) );
  DFFRX1 u_lsu_mem_data_wr_q_reg_11_ ( .D(u_lsu_N205), .CK(n37874), .RN(n44161), .QN(n2417) );
  DFFRX1 u_lsu_mem_data_wr_q_reg_19_ ( .D(u_lsu_N213), .CK(net1847), .RN(
        n44161), .QN(n2418) );
  DFFRX1 u_lsu_mem_addr_q_reg_9_ ( .D(u_lsu_mem_addr_r[9]), .CK(n37869), .RN(
        n44199), .Q(mmu_lsu_addr_w[9]), .QN(n2419) );
  DFFRX1 u_mmu_lsu_in_addr_q_reg_9_ ( .D(mmu_lsu_addr_w[9]), .CK(n37875), .RN(
        n44199), .QN(n2420) );
  DFFRX1 u_muldiv_dividend_q_reg_9_ ( .D(u_muldiv_N241), .CK(net1908), .RN(
        n44161), .Q(u_muldiv_dividend_q[9]) );
  DFFRX1 u_decode_u_regfile_reg_r26_q_reg_9_ ( .D(u_decode_u_regfile_N1034), 
        .CK(n37864), .RN(n44133), .Q(n2421), .QN(n42513) );
  DFFRX1 u_decode_u_regfile_reg_r27_q_reg_9_ ( .D(u_decode_u_regfile_N1071), 
        .CK(n37863), .RN(n44134), .Q(n2422) );
  DFFRX1 u_decode_u_regfile_reg_r1_q_reg_9_ ( .D(u_decode_u_regfile_N109), 
        .CK(n37865), .RN(n44133), .Q(n2423), .QN(n37270) );
  DFFRX1 u_decode_u_regfile_reg_r28_q_reg_9_ ( .D(u_decode_u_regfile_N1108), 
        .CK(n37862), .RN(n44133), .Q(n2424), .QN(n37090) );
  DFFRX1 u_decode_u_regfile_reg_r29_q_reg_9_ ( .D(u_decode_u_regfile_N1145), 
        .CK(n37861), .RN(n44134), .Q(n2425) );
  DFFRX1 u_decode_u_regfile_reg_r30_q_reg_9_ ( .D(u_decode_u_regfile_N1182), 
        .CK(n37860), .RN(n44133), .Q(n2426), .QN(n37080) );
  DFFRX1 u_decode_u_regfile_reg_r31_q_reg_9_ ( .D(u_decode_u_regfile_N1219), 
        .CK(n37859), .RN(n44134), .Q(n2427), .QN(n37082) );
  DFFRX1 u_decode_u_regfile_reg_r2_q_reg_9_ ( .D(u_decode_u_regfile_N146), 
        .CK(n37858), .RN(n44133), .Q(n2428) );
  DFFRX1 u_decode_u_regfile_reg_r3_q_reg_9_ ( .D(u_decode_u_regfile_N183), 
        .CK(n37857), .RN(n44134), .Q(n2429), .QN(n37258) );
  DFFRX1 u_decode_u_regfile_reg_r4_q_reg_9_ ( .D(u_decode_u_regfile_N220), 
        .CK(n37856), .RN(n44133), .Q(n2430) );
  DFFRX1 u_decode_u_regfile_reg_r5_q_reg_9_ ( .D(u_decode_u_regfile_N257), 
        .CK(n37840), .RN(n44134), .Q(n2431) );
  DFFRX1 u_decode_u_regfile_reg_r6_q_reg_9_ ( .D(u_decode_u_regfile_N294), 
        .CK(n37855), .RN(n44133), .Q(n2432) );
  DFFRX1 u_decode_u_regfile_reg_r7_q_reg_9_ ( .D(u_decode_u_regfile_N331), 
        .CK(n37854), .RN(n44134), .QN(n37087) );
  DFFRX1 u_decode_u_regfile_reg_r8_q_reg_9_ ( .D(u_decode_u_regfile_N368), 
        .CK(n37839), .RN(n44133), .Q(n2434), .QN(n37259) );
  DFFRX1 u_decode_u_regfile_reg_r9_q_reg_9_ ( .D(u_decode_u_regfile_N405), 
        .CK(n37853), .RN(n44133), .Q(n2435), .QN(n37266) );
  DFFRX1 u_decode_u_regfile_reg_r10_q_reg_9_ ( .D(u_decode_u_regfile_N442), 
        .CK(n37852), .RN(n44133), .Q(n2436) );
  DFFRX1 u_decode_u_regfile_reg_r11_q_reg_9_ ( .D(u_decode_u_regfile_N479), 
        .CK(n37851), .RN(n44134), .Q(n2437), .QN(n37264) );
  DFFRX1 u_decode_u_regfile_reg_r12_q_reg_9_ ( .D(u_decode_u_regfile_N516), 
        .CK(n37850), .RN(n44133), .Q(n2438) );
  DFFRX1 u_decode_u_regfile_reg_r13_q_reg_9_ ( .D(u_decode_u_regfile_N553), 
        .CK(n37849), .RN(n44134), .Q(n2439) );
  DFFRX1 u_decode_u_regfile_reg_r14_q_reg_9_ ( .D(u_decode_u_regfile_N590), 
        .CK(n37848), .RN(n44133), .Q(n2440) );
  DFFRX1 u_decode_u_regfile_reg_r15_q_reg_9_ ( .D(u_decode_u_regfile_N627), 
        .CK(n37847), .RN(n44134), .Q(n2441) );
  DFFRX1 u_decode_u_regfile_reg_r16_q_reg_9_ ( .D(u_decode_u_regfile_N664), 
        .CK(n37846), .RN(n44133), .Q(n2442), .QN(n37263) );
  DFFRX1 u_decode_u_regfile_reg_r17_q_reg_9_ ( .D(u_decode_u_regfile_N701), 
        .CK(n37845), .RN(n44134), .Q(n2443), .QN(n37268) );
  DFFRX1 u_decode_u_regfile_reg_r18_q_reg_9_ ( .D(u_decode_u_regfile_N738), 
        .CK(n37844), .RN(n44133), .Q(n2444), .QN(n37088) );
  DFFRX1 u_decode_u_regfile_reg_r19_q_reg_9_ ( .D(u_decode_u_regfile_N775), 
        .CK(n37843), .RN(n44134), .Q(n2445), .QN(n37252) );
  DFFRX1 u_decode_u_regfile_reg_r20_q_reg_9_ ( .D(u_decode_u_regfile_N812), 
        .CK(n37842), .RN(n44133), .Q(n2446), .QN(n37083) );
  DFFRX1 u_decode_u_regfile_reg_r21_q_reg_9_ ( .D(u_decode_u_regfile_N849), 
        .CK(n37838), .RN(n44134), .Q(n2447), .QN(n37086) );
  DFFRX1 u_decode_u_regfile_reg_r22_q_reg_9_ ( .D(u_decode_u_regfile_N886), 
        .CK(n37841), .RN(n44133), .Q(n2448), .QN(n37076) );
  DFFRX1 u_decode_u_regfile_reg_r23_q_reg_9_ ( .D(u_decode_u_regfile_N923), 
        .CK(n37877), .RN(n44134), .Q(n2449) );
  DFFRX1 u_decode_u_regfile_reg_r24_q_reg_9_ ( .D(u_decode_u_regfile_N960), 
        .CK(n37878), .RN(n44133), .Q(n2450), .QN(n37269) );
  DFFRX1 u_lsu_mem_addr_q_reg_23_ ( .D(u_lsu_mem_addr_r[23]), .CK(n37876), 
        .RN(n44185), .Q(mmu_lsu_addr_w[23]), .QN(n8320) );
  DFFRX1 u_mmu_lsu_in_addr_q_reg_23_ ( .D(mmu_lsu_addr_w[23]), .CK(n37873), 
        .RN(n44185), .QN(n2451) );
  DFFRX1 u_mmu_itlb_va_addr_q_reg_23_ ( .D(n8438), .CK(clk_i), .RN(n44185), 
        .Q(u_mmu_itlb_va_addr_q[23]) );
  DFFRX1 u_mmu_dtlb_va_addr_q_reg_23_ ( .D(n8437), .CK(clk_i), .RN(n44206), 
        .Q(u_mmu_dtlb_va_addr_q[23]) );
  DFFRX1 u_decode_u_regfile_reg_r25_q_reg_23_ ( .D(u_decode_u_regfile_N1011), 
        .CK(n37837), .RN(n44094), .Q(n2453), .QN(n40858) );
  DFFRX1 u_decode_u_regfile_reg_r26_q_reg_23_ ( .D(u_decode_u_regfile_N1048), 
        .CK(n37836), .RN(n44093), .Q(n2454), .QN(n36970) );
  DFFRX1 u_decode_u_regfile_reg_r27_q_reg_23_ ( .D(u_decode_u_regfile_N1085), 
        .CK(n37835), .RN(n44094), .Q(n2455), .QN(n42466) );
  DFFRX1 u_decode_u_regfile_reg_r28_q_reg_23_ ( .D(u_decode_u_regfile_N1122), 
        .CK(n37834), .RN(n44093), .Q(n2456) );
  DFFRX1 u_decode_u_regfile_reg_r29_q_reg_23_ ( .D(u_decode_u_regfile_N1159), 
        .CK(n37833), .RN(n44094), .Q(n2457) );
  DFFRX1 u_decode_u_regfile_reg_r30_q_reg_23_ ( .D(u_decode_u_regfile_N1196), 
        .CK(n37832), .RN(n44094), .Q(n2458) );
  DFFRX1 u_decode_u_regfile_reg_r1_q_reg_23_ ( .D(u_decode_u_regfile_N123), 
        .CK(n37830), .RN(n44094), .Q(n2459) );
  DFFRX1 u_decode_u_regfile_reg_r31_q_reg_23_ ( .D(u_decode_u_regfile_N1233), 
        .CK(n37831), .RN(n44095), .Q(n2460) );
  DFFRX1 u_decode_u_regfile_reg_r2_q_reg_23_ ( .D(u_decode_u_regfile_N160), 
        .CK(n37829), .RN(n44093), .Q(n2461), .QN(n36955) );
  DFFRX1 u_decode_u_regfile_reg_r3_q_reg_23_ ( .D(u_decode_u_regfile_N197), 
        .CK(n37828), .RN(n44094), .Q(n2462) );
  DFFRX1 u_decode_u_regfile_reg_r4_q_reg_23_ ( .D(u_decode_u_regfile_N234), 
        .CK(n37827), .RN(n44093), .Q(n2463), .QN(n36984) );
  DFFRX1 u_decode_u_regfile_reg_r5_q_reg_23_ ( .D(u_decode_u_regfile_N271), 
        .CK(n37826), .RN(n44094), .Q(n2464), .QN(n36952) );
  DFFRX1 u_decode_u_regfile_reg_r6_q_reg_23_ ( .D(u_decode_u_regfile_N308), 
        .CK(n37825), .RN(n44094), .Q(n2465), .QN(n36938) );
  DFFRX1 u_decode_u_regfile_reg_r8_q_reg_23_ ( .D(u_decode_u_regfile_N382), 
        .CK(n37823), .RN(n44093), .Q(n2467) );
  DFFRX1 u_decode_u_regfile_reg_r9_q_reg_23_ ( .D(u_decode_u_regfile_N419), 
        .CK(n37822), .RN(n44094), .Q(n2468) );
  DFFRX1 u_decode_u_regfile_reg_r10_q_reg_23_ ( .D(u_decode_u_regfile_N456), 
        .CK(n37821), .RN(n44093), .Q(n2469), .QN(n36968) );
  DFFRX1 u_decode_u_regfile_reg_r11_q_reg_23_ ( .D(u_decode_u_regfile_N493), 
        .CK(n37820), .RN(n44094), .Q(n2470), .QN(n38678) );
  DFFRX1 u_decode_u_regfile_reg_r12_q_reg_23_ ( .D(u_decode_u_regfile_N530), 
        .CK(n37819), .RN(n44093), .Q(n2471), .QN(n36978) );
  DFFRX1 u_decode_u_regfile_reg_r13_q_reg_23_ ( .D(u_decode_u_regfile_N567), 
        .CK(n37818), .RN(n44094), .Q(n2472) );
  DFFRX1 u_decode_u_regfile_reg_r14_q_reg_23_ ( .D(u_decode_u_regfile_N604), 
        .CK(n37817), .RN(n44094), .Q(n2473), .QN(n36958) );
  DFFRX1 u_decode_u_regfile_reg_r15_q_reg_23_ ( .D(u_decode_u_regfile_N641), 
        .CK(n37816), .RN(n44094), .Q(n2474) );
  DFFRX1 u_decode_u_regfile_reg_r16_q_reg_23_ ( .D(u_decode_u_regfile_N678), 
        .CK(n37815), .RN(n44093), .Q(n2475), .QN(n37096) );
  DFFRX1 u_decode_u_regfile_reg_r17_q_reg_23_ ( .D(u_decode_u_regfile_N715), 
        .CK(n37814), .RN(n44094), .Q(n2476), .QN(n37107) );
  DFFRX1 u_decode_u_regfile_reg_r18_q_reg_23_ ( .D(u_decode_u_regfile_N752), 
        .CK(n37813), .RN(n44093), .Q(n2477) );
  DFFRX1 u_decode_u_regfile_reg_r19_q_reg_23_ ( .D(u_decode_u_regfile_N789), 
        .CK(n37812), .RN(n44094), .Q(n2478), .QN(n37111) );
  DFFRX1 u_decode_u_regfile_reg_r20_q_reg_23_ ( .D(u_decode_u_regfile_N826), 
        .CK(n37811), .RN(n44093), .Q(n2479), .QN(n36946) );
  DFFRX1 u_decode_u_regfile_reg_r21_q_reg_23_ ( .D(u_decode_u_regfile_N863), 
        .CK(n37810), .RN(n44094), .Q(n2480), .QN(n36950) );
  DFFRX1 u_decode_u_regfile_reg_r22_q_reg_23_ ( .D(u_decode_u_regfile_N900), 
        .CK(n37809), .RN(n44094), .Q(n2481), .QN(n36951) );
  DFFRX1 u_decode_u_regfile_reg_r23_q_reg_23_ ( .D(u_decode_u_regfile_N937), 
        .CK(n37880), .RN(n44094), .Q(n2482), .QN(n36995) );
  DFFRX1 u_lsu_mem_addr_q_reg_22_ ( .D(u_lsu_mem_addr_r[22]), .CK(n37876), 
        .RN(n44182), .Q(mmu_lsu_addr_w[22]), .QN(n8318) );
  DFFRX1 u_mmu_lsu_in_addr_q_reg_22_ ( .D(mmu_lsu_addr_w[22]), .CK(n37873), 
        .RN(n44182), .QN(n2483) );
  DFFRX1 u_mmu_itlb_va_addr_q_reg_22_ ( .D(n8436), .CK(clk_i), .RN(n44182), 
        .Q(u_mmu_itlb_va_addr_q[22]) );
  DFFRX1 u_mmu_dtlb_va_addr_q_reg_22_ ( .D(n8435), .CK(clk_i), .RN(n44206), 
        .Q(u_mmu_dtlb_va_addr_q[22]) );
  DFFRX1 u_decode_u_regfile_reg_r25_q_reg_22_ ( .D(u_decode_u_regfile_N1010), 
        .CK(n37837), .RN(n44092), .Q(n2485), .QN(n40854) );
  DFFRX1 u_decode_u_regfile_reg_r26_q_reg_22_ ( .D(u_decode_u_regfile_N1047), 
        .CK(n37836), .RN(n44091), .Q(n2486) );
  DFFRX1 u_decode_u_regfile_reg_r27_q_reg_22_ ( .D(u_decode_u_regfile_N1084), 
        .CK(n37835), .RN(n44092), .Q(n2487) );
  DFFRX1 u_decode_u_regfile_reg_r28_q_reg_22_ ( .D(u_decode_u_regfile_N1121), 
        .CK(n37834), .RN(n44092), .Q(n2488), .QN(n37011) );
  DFFRX1 u_decode_u_regfile_reg_r29_q_reg_22_ ( .D(u_decode_u_regfile_N1158), 
        .CK(n37833), .RN(n44092), .Q(n2489), .QN(n37014) );
  DFFRX1 u_decode_u_regfile_reg_r30_q_reg_22_ ( .D(u_decode_u_regfile_N1195), 
        .CK(n37832), .RN(n44092), .Q(n2490), .QN(n36989) );
  DFFRX1 u_decode_u_regfile_reg_r1_q_reg_22_ ( .D(u_decode_u_regfile_N122), 
        .CK(n37830), .RN(n44092), .Q(n2491) );
  DFFRX1 u_decode_u_regfile_reg_r31_q_reg_22_ ( .D(u_decode_u_regfile_N1232), 
        .CK(n37831), .RN(n44093), .Q(n2492) );
  DFFRX1 u_decode_u_regfile_reg_r2_q_reg_22_ ( .D(u_decode_u_regfile_N159), 
        .CK(n37829), .RN(n44091), .Q(n2493), .QN(n37005) );
  DFFRX1 u_decode_u_regfile_reg_r3_q_reg_22_ ( .D(u_decode_u_regfile_N196), 
        .CK(n37828), .RN(n44092), .Q(n2494) );
  DFFRX1 u_decode_u_regfile_reg_r4_q_reg_22_ ( .D(u_decode_u_regfile_N233), 
        .CK(n37827), .RN(n44092), .Q(n2495) );
  DFFRX1 u_decode_u_regfile_reg_r5_q_reg_22_ ( .D(u_decode_u_regfile_N270), 
        .CK(n37826), .RN(n44092), .Q(n2496), .QN(n37000) );
  DFFRX1 u_decode_u_regfile_reg_r6_q_reg_22_ ( .D(u_decode_u_regfile_N307), 
        .CK(n37825), .RN(n44092), .Q(n2497) );
  DFFRX1 u_decode_u_regfile_reg_r7_q_reg_22_ ( .D(u_decode_u_regfile_N344), 
        .CK(n37824), .RN(n44093), .Q(n2498), .QN(n37317) );
  DFFRX1 u_decode_u_regfile_reg_r8_q_reg_22_ ( .D(u_decode_u_regfile_N381), 
        .CK(n37823), .RN(n44091), .Q(n2499) );
  DFFRX1 u_decode_u_regfile_reg_r9_q_reg_22_ ( .D(u_decode_u_regfile_N418), 
        .CK(n37822), .RN(n44092), .Q(n2500) );
  DFFRX1 u_decode_u_regfile_reg_r10_q_reg_22_ ( .D(u_decode_u_regfile_N455), 
        .CK(n37821), .RN(n44091), .Q(n2501), .QN(n37009) );
  DFFRX1 u_decode_u_regfile_reg_r11_q_reg_22_ ( .D(u_decode_u_regfile_N492), 
        .CK(n37820), .RN(n44092), .Q(n2502) );
  DFFRX1 u_decode_u_regfile_reg_r12_q_reg_22_ ( .D(u_decode_u_regfile_N529), 
        .CK(n37819), .RN(n44092), .Q(n2503), .QN(n37016) );
  DFFRX1 u_decode_u_regfile_reg_r13_q_reg_22_ ( .D(u_decode_u_regfile_N566), 
        .CK(n37818), .RN(n44093), .Q(n2504), .QN(n37003) );
  DFFRX1 u_decode_u_regfile_reg_r14_q_reg_22_ ( .D(u_decode_u_regfile_N603), 
        .CK(n37817), .RN(n44092), .Q(n2505), .QN(n37008) );
  DFFRX1 u_decode_u_regfile_reg_r15_q_reg_22_ ( .D(u_decode_u_regfile_N640), 
        .CK(n37816), .RN(n44093), .Q(n2506) );
  DFFRX1 u_decode_u_regfile_reg_r16_q_reg_22_ ( .D(u_decode_u_regfile_N677), 
        .CK(n37815), .RN(n44091), .Q(n2507) );
  DFFRX1 u_decode_u_regfile_reg_r17_q_reg_22_ ( .D(u_decode_u_regfile_N714), 
        .CK(n37814), .RN(n44092), .Q(n2508) );
  DFFRX1 u_decode_u_regfile_reg_r18_q_reg_22_ ( .D(u_decode_u_regfile_N751), 
        .CK(n37813), .RN(n44091), .Q(n2509), .QN(n40856) );
  DFFRX1 u_decode_u_regfile_reg_r19_q_reg_22_ ( .D(u_decode_u_regfile_N788), 
        .CK(n37812), .RN(n44092), .Q(n2510), .QN(n37151) );
  DFFRX1 u_decode_u_regfile_reg_r20_q_reg_22_ ( .D(u_decode_u_regfile_N825), 
        .CK(n37811), .RN(n44092), .Q(n2511) );
  DFFRX1 u_decode_u_regfile_reg_r21_q_reg_22_ ( .D(u_decode_u_regfile_N862), 
        .CK(n37810), .RN(n44093), .Q(n2512), .QN(n37002) );
  DFFRX1 u_decode_u_regfile_reg_r22_q_reg_22_ ( .D(u_decode_u_regfile_N899), 
        .CK(n37809), .RN(n44092), .Q(n2513) );
  DFFRX1 u_decode_u_regfile_reg_r23_q_reg_22_ ( .D(u_decode_u_regfile_N936), 
        .CK(n37880), .RN(n44093), .Q(n2514), .QN(n36996) );
  DFFRX1 u_lsu_mem_data_wr_q_reg_22_ ( .D(u_lsu_N216), .CK(net1847), .RN(
        n44160), .QN(n2515) );
  DFFRX1 u_lsu_mem_addr_q_reg_16_ ( .D(u_lsu_mem_addr_r[16]), .CK(n37876), 
        .RN(n44184), .Q(mmu_lsu_addr_w[16]), .QN(n8304) );
  DFFRX1 u_mmu_lsu_in_addr_q_reg_16_ ( .D(mmu_lsu_addr_w[16]), .CK(n37873), 
        .RN(n44184), .QN(n2516) );
  DFFRX1 u_mmu_itlb_va_addr_q_reg_16_ ( .D(u_mmu_virt_addr_q[16]), .CK(n37871), 
        .RN(n44184), .Q(n2517) );
  DFFRX1 u_mmu_dtlb_va_addr_q_reg_16_ ( .D(u_mmu_virt_addr_q[16]), .CK(n37872), 
        .RN(n44207), .Q(u_mmu_dtlb_va_addr_q[16]) );
  DFFRX1 u_mmu_itlb_entry_q_reg_16_ ( .D(u_mmu_pte_entry_q[16]), .CK(net1792), 
        .RN(n44171), .Q(u_mmu_itlb_entry_q[16]) );
  DFFRX1 u_mmu_dtlb_entry_q_reg_16_ ( .D(u_mmu_pte_entry_q[16]), .CK(net1782), 
        .RN(n44196), .QN(n2518) );
  DFFRX1 u_muldiv_dividend_q_reg_16_ ( .D(u_muldiv_N248), .CK(net1913), .RN(
        n44160), .Q(u_muldiv_dividend_q[16]), .QN(n37451) );
  DFFRX1 u_decode_u_regfile_reg_r25_q_reg_16_ ( .D(u_decode_u_regfile_N1004), 
        .CK(n37837), .RN(n44097), .Q(n2519), .QN(n37170) );
  DFFRX1 u_decode_u_regfile_reg_r26_q_reg_16_ ( .D(u_decode_u_regfile_N1041), 
        .CK(n37836), .RN(n44097), .Q(n2520) );
  DFFRX1 u_decode_u_regfile_reg_r27_q_reg_16_ ( .D(u_decode_u_regfile_N1078), 
        .CK(n37835), .RN(n44098), .Q(n2521) );
  DFFRX1 u_decode_u_regfile_reg_r28_q_reg_16_ ( .D(u_decode_u_regfile_N1115), 
        .CK(n37834), .RN(n44097), .Q(n2522), .QN(n36874) );
  DFFRX1 u_decode_u_regfile_reg_r29_q_reg_16_ ( .D(u_decode_u_regfile_N1152), 
        .CK(n37833), .RN(n44098), .Q(n2523) );
  DFFRX1 u_decode_u_regfile_reg_r1_q_reg_16_ ( .D(u_decode_u_regfile_N116), 
        .CK(n37830), .RN(n44097), .Q(n2524), .QN(n37172) );
  DFFRX1 u_decode_u_regfile_reg_r30_q_reg_16_ ( .D(u_decode_u_regfile_N1189), 
        .CK(n37832), .RN(n44097), .Q(n2525), .QN(n36867) );
  DFFRX1 u_decode_u_regfile_reg_r31_q_reg_16_ ( .D(u_decode_u_regfile_N1226), 
        .CK(n37831), .RN(n44098), .Q(n2526), .QN(n36871) );
  DFFRX1 u_decode_u_regfile_reg_r2_q_reg_16_ ( .D(u_decode_u_regfile_N153), 
        .CK(n37829), .RN(n44097), .Q(n2527) );
  DFFRX1 u_decode_u_regfile_reg_r3_q_reg_16_ ( .D(u_decode_u_regfile_N190), 
        .CK(n37828), .RN(n44098), .Q(n2528), .QN(n37120) );
  DFFRX1 u_decode_u_regfile_reg_r4_q_reg_16_ ( .D(u_decode_u_regfile_N227), 
        .CK(n37827), .RN(n44097), .Q(n2529) );
  DFFRX1 u_decode_u_regfile_reg_r5_q_reg_16_ ( .D(u_decode_u_regfile_N264), 
        .CK(n37826), .RN(n44098), .Q(n2530) );
  DFFRX1 u_decode_u_regfile_reg_r6_q_reg_16_ ( .D(u_decode_u_regfile_N301), 
        .CK(n37825), .RN(n44097), .Q(n2531) );
  DFFRX1 u_decode_u_regfile_reg_r7_q_reg_16_ ( .D(u_decode_u_regfile_N338), 
        .CK(n37824), .RN(n44098), .QN(n36875) );
  DFFRX1 u_decode_u_regfile_reg_r8_q_reg_16_ ( .D(u_decode_u_regfile_N375), 
        .CK(n37823), .RN(n44097), .Q(n2533), .QN(n37164) );
  DFFRX1 u_decode_u_regfile_reg_r9_q_reg_16_ ( .D(u_decode_u_regfile_N412), 
        .CK(n37822), .RN(n44097), .Q(n2534), .QN(n37192) );
  DFFRX1 u_decode_u_regfile_reg_r10_q_reg_16_ ( .D(u_decode_u_regfile_N449), 
        .CK(n37821), .RN(n44097), .Q(n2535) );
  DFFRX1 u_decode_u_regfile_reg_r11_q_reg_16_ ( .D(u_decode_u_regfile_N486), 
        .CK(n37820), .RN(n44098), .Q(n2536), .QN(n37168) );
  DFFRX1 u_decode_u_regfile_reg_r12_q_reg_16_ ( .D(u_decode_u_regfile_N523), 
        .CK(n37819), .RN(n44097), .Q(n2537) );
  DFFRX1 u_decode_u_regfile_reg_r13_q_reg_16_ ( .D(u_decode_u_regfile_N560), 
        .CK(n37818), .RN(n44098), .Q(n2538) );
  DFFRX1 u_decode_u_regfile_reg_r14_q_reg_16_ ( .D(u_decode_u_regfile_N597), 
        .CK(n37817), .RN(n44097), .Q(n2539) );
  DFFRX1 u_decode_u_regfile_reg_r15_q_reg_16_ ( .D(u_decode_u_regfile_N634), 
        .CK(n37816), .RN(n44098), .Q(n2540), .QN(n36876) );
  DFFRX1 u_decode_u_regfile_reg_r16_q_reg_16_ ( .D(u_decode_u_regfile_N671), 
        .CK(n37815), .RN(n44096), .Q(n2541), .QN(n37154) );
  DFFRX1 u_decode_u_regfile_reg_r17_q_reg_16_ ( .D(u_decode_u_regfile_N708), 
        .CK(n37814), .RN(n44097), .Q(n2542), .QN(n37160) );
  DFFRX1 u_decode_u_regfile_reg_r18_q_reg_16_ ( .D(u_decode_u_regfile_N745), 
        .CK(n37813), .RN(n44097), .Q(n2543), .QN(n36879) );
  DFFRX1 u_decode_u_regfile_reg_r19_q_reg_16_ ( .D(u_decode_u_regfile_N782), 
        .CK(n37812), .RN(n44098), .Q(n2544), .QN(n37119) );
  DFFRX1 u_decode_u_regfile_reg_r20_q_reg_16_ ( .D(u_decode_u_regfile_N819), 
        .CK(n37811), .RN(n44097), .Q(n2545), .QN(n36872) );
  DFFRX1 u_decode_u_regfile_reg_r21_q_reg_16_ ( .D(u_decode_u_regfile_N856), 
        .CK(n37810), .RN(n44098), .Q(n2546) );
  DFFRX1 u_decode_u_regfile_reg_r22_q_reg_16_ ( .D(u_decode_u_regfile_N893), 
        .CK(n37809), .RN(n44097), .Q(n2547), .QN(n36865) );
  DFFRX1 u_decode_u_regfile_reg_r23_q_reg_16_ ( .D(u_decode_u_regfile_N930), 
        .CK(n37880), .RN(n44098), .Q(n2548) );
  DFFRX1 u_lsu_mem_addr_q_reg_21_ ( .D(u_lsu_mem_addr_r[21]), .CK(n37876), 
        .RN(n44184), .Q(mmu_lsu_addr_w[21]), .QN(n8316) );
  DFFRX1 u_mmu_lsu_in_addr_q_reg_21_ ( .D(mmu_lsu_addr_w[21]), .CK(n37873), 
        .RN(n44184), .QN(n2549) );
  DFFRX1 u_mmu_itlb_va_addr_q_reg_21_ ( .D(u_mmu_virt_addr_q[21]), .CK(n37871), 
        .RN(n44185), .Q(u_mmu_itlb_va_addr_q[21]) );
  DFFRX1 u_mmu_dtlb_va_addr_q_reg_21_ ( .D(n8434), .CK(clk_i), .RN(n44206), 
        .Q(u_mmu_dtlb_va_addr_q[21]) );
  DFFRX1 u_mmu_itlb_entry_q_reg_21_ ( .D(u_mmu_pte_entry_q[21]), .CK(net1792), 
        .RN(n44171), .Q(u_mmu_itlb_entry_q[21]) );
  DFFRX1 u_mmu_dtlb_entry_q_reg_21_ ( .D(u_mmu_pte_entry_q[21]), .CK(net1782), 
        .RN(n44197), .QN(n2550) );
  DFFRX1 u_decode_u_regfile_reg_r25_q_reg_21_ ( .D(u_decode_u_regfile_N1009), 
        .CK(n37837), .RN(n44090), .Q(n2551), .QN(n37142) );
  DFFRX1 u_decode_u_regfile_reg_r26_q_reg_21_ ( .D(u_decode_u_regfile_N1046), 
        .CK(n37836), .RN(n44090), .Q(n2552), .QN(n36962) );
  DFFRX1 u_decode_u_regfile_reg_r27_q_reg_21_ ( .D(u_decode_u_regfile_N1083), 
        .CK(n37835), .RN(n44090), .Q(n2553) );
  DFFRX1 u_decode_u_regfile_reg_r28_q_reg_21_ ( .D(u_decode_u_regfile_N1120), 
        .CK(n37834), .RN(n44090), .Q(n2554) );
  DFFRX1 u_decode_u_regfile_reg_r29_q_reg_21_ ( .D(u_decode_u_regfile_N1157), 
        .CK(n37833), .RN(n44091), .Q(n2555), .QN(n36986) );
  DFFRX1 u_decode_u_regfile_reg_r1_q_reg_21_ ( .D(u_decode_u_regfile_N121), 
        .CK(n37830), .RN(n44090), .Q(n2557) );
  DFFRX1 u_decode_u_regfile_reg_r31_q_reg_21_ ( .D(u_decode_u_regfile_N1231), 
        .CK(n37831), .RN(n44091), .Q(n2558) );
  DFFRX1 u_decode_u_regfile_reg_r2_q_reg_21_ ( .D(u_decode_u_regfile_N158), 
        .CK(n37829), .RN(n44090), .Q(n2559), .QN(n36979) );
  DFFRX1 u_decode_u_regfile_reg_r3_q_reg_21_ ( .D(u_decode_u_regfile_N195), 
        .CK(n37828), .RN(n44090), .Q(n2560) );
  DFFRX1 u_decode_u_regfile_reg_r4_q_reg_21_ ( .D(u_decode_u_regfile_N232), 
        .CK(n37827), .RN(n44090), .Q(n2561) );
  DFFRX1 u_decode_u_regfile_reg_r5_q_reg_21_ ( .D(u_decode_u_regfile_N269), 
        .CK(n37826), .RN(n44091), .Q(n2562), .QN(n36981) );
  DFFRX1 u_decode_u_regfile_reg_r6_q_reg_21_ ( .D(u_decode_u_regfile_N306), 
        .CK(n37825), .RN(n44090), .Q(n2563), .QN(n36990) );
  DFFRX1 u_decode_u_regfile_reg_r8_q_reg_21_ ( .D(u_decode_u_regfile_N380), 
        .CK(n37823), .RN(n44089), .Q(n2565), .QN(n37139) );
  DFFRX1 u_decode_u_regfile_reg_r9_q_reg_21_ ( .D(u_decode_u_regfile_N417), 
        .CK(n37822), .RN(n44090), .Q(n2566), .QN(n40846) );
  DFFRX1 u_decode_u_regfile_reg_r10_q_reg_21_ ( .D(u_decode_u_regfile_N454), 
        .CK(n37821), .RN(n44089), .Q(n2567), .QN(n36999) );
  DFFRX1 u_decode_u_regfile_reg_r11_q_reg_21_ ( .D(u_decode_u_regfile_N491), 
        .CK(n37820), .RN(n44091), .Q(n2568), .QN(n37130) );
  DFFRX1 u_decode_u_regfile_reg_r12_q_reg_21_ ( .D(u_decode_u_regfile_N528), 
        .CK(n37819), .RN(n44090), .Q(n2569), .QN(n36971) );
  DFFRX1 u_decode_u_regfile_reg_r13_q_reg_21_ ( .D(u_decode_u_regfile_N565), 
        .CK(n37818), .RN(n44091), .Q(n2570), .QN(n36973) );
  DFFRX1 u_decode_u_regfile_reg_r14_q_reg_21_ ( .D(u_decode_u_regfile_N602), 
        .CK(n37817), .RN(n44090), .Q(n2571), .QN(n36953) );
  DFFRX1 u_decode_u_regfile_reg_r15_q_reg_21_ ( .D(u_decode_u_regfile_N639), 
        .CK(n37816), .RN(n44091), .Q(n2572), .QN(n36948) );
  DFFRX1 u_decode_u_regfile_reg_r16_q_reg_21_ ( .D(u_decode_u_regfile_N676), 
        .CK(n37815), .RN(n44089), .Q(n2573), .QN(n37095) );
  DFFRX1 u_decode_u_regfile_reg_r17_q_reg_21_ ( .D(u_decode_u_regfile_N713), 
        .CK(n37814), .RN(n44090), .Q(n2574), .QN(n37137) );
  DFFRX1 u_decode_u_regfile_reg_r18_q_reg_21_ ( .D(u_decode_u_regfile_N750), 
        .CK(n37813), .RN(n44090), .Q(n2575) );
  DFFRX1 u_decode_u_regfile_reg_r19_q_reg_21_ ( .D(u_decode_u_regfile_N787), 
        .CK(n37812), .RN(n44090), .Q(n2576), .QN(n37136) );
  DFFRX1 u_decode_u_regfile_reg_r20_q_reg_21_ ( .D(u_decode_u_regfile_N824), 
        .CK(n37811), .RN(n44090), .Q(n2577) );
  DFFRX1 u_decode_u_regfile_reg_r21_q_reg_21_ ( .D(u_decode_u_regfile_N861), 
        .CK(n37810), .RN(n44091), .Q(n2578) );
  DFFRX1 u_decode_u_regfile_reg_r22_q_reg_21_ ( .D(u_decode_u_regfile_N898), 
        .CK(n37809), .RN(n44090), .Q(n2579) );
  DFFRX1 u_decode_u_regfile_reg_r23_q_reg_21_ ( .D(u_decode_u_regfile_N935), 
        .CK(n37880), .RN(n44091), .Q(n2580), .QN(n36959) );
  DFFRX1 u_lsu_mem_addr_q_reg_7_ ( .D(u_lsu_mem_addr_r[7]), .CK(n37869), .RN(
        n44199), .Q(mmu_lsu_addr_w[7]), .QN(n2581) );
  DFFRX1 u_mmu_lsu_in_addr_q_reg_7_ ( .D(mmu_lsu_addr_w[7]), .CK(n37875), .RN(
        n44199), .QN(n2582) );
  DFFRX1 u_muldiv_dividend_q_reg_7_ ( .D(u_muldiv_N239), .CK(net1908), .RN(
        n44160), .Q(u_muldiv_dividend_q[7]), .QN(n37426) );
  DFFRX1 u_decode_u_regfile_reg_r26_q_reg_7_ ( .D(u_decode_u_regfile_N1032), 
        .CK(n37864), .RN(n44140), .Q(n2583) );
  DFFRX1 u_decode_u_regfile_reg_r27_q_reg_7_ ( .D(u_decode_u_regfile_N1069), 
        .CK(n37863), .RN(n44141), .Q(n2584) );
  DFFRX1 u_decode_u_regfile_reg_r1_q_reg_7_ ( .D(u_decode_u_regfile_N107), 
        .CK(n37865), .RN(n44141), .Q(n2585), .QN(n37216) );
  DFFRX1 u_decode_u_regfile_reg_r28_q_reg_7_ ( .D(u_decode_u_regfile_N1106), 
        .CK(n37862), .RN(n44140), .Q(n2586), .QN(n36873) );
  DFFRX1 u_decode_u_regfile_reg_r29_q_reg_7_ ( .D(u_decode_u_regfile_N1143), 
        .CK(n37861), .RN(n44140), .Q(n2587) );
  DFFRX1 u_decode_u_regfile_reg_r30_q_reg_7_ ( .D(u_decode_u_regfile_N1180), 
        .CK(n37860), .RN(n44141), .Q(n2588), .QN(n36923) );
  DFFRX1 u_decode_u_regfile_reg_r31_q_reg_7_ ( .D(u_decode_u_regfile_N1217), 
        .CK(n37859), .RN(n44127), .Q(n2589), .QN(n36922) );
  DFFRX1 u_decode_u_regfile_reg_r2_q_reg_7_ ( .D(u_decode_u_regfile_N144), 
        .CK(n37858), .RN(n44140), .Q(n2590) );
  DFFRX1 u_decode_u_regfile_reg_r3_q_reg_7_ ( .D(u_decode_u_regfile_N181), 
        .CK(n37857), .RN(n44141), .Q(n2591), .QN(n37200) );
  DFFRX1 u_decode_u_regfile_reg_r4_q_reg_7_ ( .D(u_decode_u_regfile_N218), 
        .CK(n37856), .RN(n44140), .Q(n2592) );
  DFFRX1 u_decode_u_regfile_reg_r5_q_reg_7_ ( .D(u_decode_u_regfile_N255), 
        .CK(n37840), .RN(n44140), .Q(n2593) );
  DFFRX1 u_decode_u_regfile_reg_r6_q_reg_7_ ( .D(u_decode_u_regfile_N292), 
        .CK(n37855), .RN(n44140), .Q(n2594) );
  DFFRX1 u_decode_u_regfile_reg_r7_q_reg_7_ ( .D(u_decode_u_regfile_N329), 
        .CK(n37854), .RN(n44144), .QN(n36932) );
  DFFRX1 u_decode_u_regfile_reg_r8_q_reg_7_ ( .D(u_decode_u_regfile_N366), 
        .CK(n37839), .RN(n44141), .Q(n2596), .QN(n37202) );
  DFFRX1 u_decode_u_regfile_reg_r9_q_reg_7_ ( .D(u_decode_u_regfile_N403), 
        .CK(n37853), .RN(n44141), .Q(n2597), .QN(n37209) );
  DFFRX1 u_decode_u_regfile_reg_r10_q_reg_7_ ( .D(u_decode_u_regfile_N440), 
        .CK(n37852), .RN(n44140), .Q(n2598) );
  DFFRX1 u_decode_u_regfile_reg_r11_q_reg_7_ ( .D(u_decode_u_regfile_N477), 
        .CK(n37851), .RN(n44141), .Q(n2599), .QN(n37208) );
  DFFRX1 u_decode_u_regfile_reg_r12_q_reg_7_ ( .D(u_decode_u_regfile_N514), 
        .CK(n37850), .RN(n44141), .Q(n2600) );
  DFFRX1 u_decode_u_regfile_reg_r13_q_reg_7_ ( .D(u_decode_u_regfile_N551), 
        .CK(n37849), .RN(n44140), .Q(n2601) );
  DFFRX1 u_decode_u_regfile_reg_r14_q_reg_7_ ( .D(u_decode_u_regfile_N588), 
        .CK(n37848), .RN(n44141), .Q(n2602) );
  DFFRX1 u_decode_u_regfile_reg_r15_q_reg_7_ ( .D(u_decode_u_regfile_N625), 
        .CK(n37847), .RN(n44141), .Q(n2603) );
  DFFRX1 u_decode_u_regfile_reg_r16_q_reg_7_ ( .D(u_decode_u_regfile_N662), 
        .CK(n37846), .RN(n44141), .Q(n2604), .QN(n37207) );
  DFFRX1 u_decode_u_regfile_reg_r17_q_reg_7_ ( .D(u_decode_u_regfile_N699), 
        .CK(n37845), .RN(n44141), .Q(n2605), .QN(n37214) );
  DFFRX1 u_decode_u_regfile_reg_r18_q_reg_7_ ( .D(u_decode_u_regfile_N736), 
        .CK(n37844), .RN(n44140), .Q(n2606), .QN(n36934) );
  DFFRX1 u_decode_u_regfile_reg_r19_q_reg_7_ ( .D(u_decode_u_regfile_N773), 
        .CK(n37843), .RN(n44141), .Q(n2607), .QN(n37195) );
  DFFRX1 u_decode_u_regfile_reg_r20_q_reg_7_ ( .D(u_decode_u_regfile_N810), 
        .CK(n37842), .RN(n44140), .Q(n2608), .QN(n36925) );
  DFFRX1 u_decode_u_regfile_reg_r21_q_reg_7_ ( .D(u_decode_u_regfile_N847), 
        .CK(n37838), .RN(n44141), .Q(n2609), .QN(n36933) );
  DFFRX1 u_decode_u_regfile_reg_r22_q_reg_7_ ( .D(u_decode_u_regfile_N884), 
        .CK(n37841), .RN(n44140), .Q(n2610), .QN(n36916) );
  DFFRX1 u_decode_u_regfile_reg_r23_q_reg_7_ ( .D(u_decode_u_regfile_N921), 
        .CK(n37877), .RN(n44140), .Q(n2611), .QN(n38918) );
  DFFRX1 u_decode_u_regfile_reg_r24_q_reg_7_ ( .D(u_decode_u_regfile_N958), 
        .CK(n37878), .RN(n44141), .Q(n2612) );
  DFFRX1 u_lsu_mem_data_wr_q_reg_7_ ( .D(u_lsu_N201), .CK(n37874), .RN(n44200), 
        .QN(n2613) );
  DFFRX1 u_lsu_mem_data_wr_q_reg_15_ ( .D(u_lsu_N209), .CK(net1847), .RN(
        n44160), .QN(n2614) );
  DFFRX1 u_lsu_mem_data_wr_q_reg_23_ ( .D(u_lsu_N217), .CK(net1847), .RN(
        n44160), .QN(n2615) );
  DFFRX1 u_lsu_mem_data_wr_q_reg_31_ ( .D(u_lsu_N225), .CK(n37868), .RN(n44160), .QN(n2616) );
  DFFRX1 u_lsu_mem_addr_q_reg_26_ ( .D(u_lsu_mem_addr_r[26]), .CK(n37876), 
        .RN(n44116), .Q(mmu_lsu_addr_w[26]), .QN(n8326) );
  DFFRX1 u_mmu_lsu_in_addr_q_reg_26_ ( .D(mmu_lsu_addr_w[26]), .CK(n37873), 
        .RN(n44116), .QN(n2617) );
  DFFRX1 u_mmu_itlb_va_addr_q_reg_26_ ( .D(n8433), .CK(clk_i), .RN(n44189), 
        .Q(u_mmu_itlb_va_addr_q[26]) );
  DFFRX1 u_mmu_dtlb_va_addr_q_reg_26_ ( .D(n8432), .CK(clk_i), .RN(n44206), 
        .Q(u_mmu_dtlb_va_addr_q[26]) );
  DFFRX1 u_decode_u_regfile_reg_r25_q_reg_26_ ( .D(u_decode_u_regfile_N1014), 
        .CK(n37837), .RN(n44115), .Q(n2619), .QN(n37108) );
  DFFRX1 u_decode_u_regfile_reg_r26_q_reg_26_ ( .D(u_decode_u_regfile_N1051), 
        .CK(n37836), .RN(n44115), .Q(n2620) );
  DFFRX1 u_decode_u_regfile_reg_r27_q_reg_26_ ( .D(u_decode_u_regfile_N1088), 
        .CK(n37835), .RN(n44116), .Q(n2621), .QN(n42482) );
  DFFRX1 u_decode_u_regfile_reg_r28_q_reg_26_ ( .D(u_decode_u_regfile_N1125), 
        .CK(n37834), .RN(n44115), .Q(n2622) );
  DFFRX1 u_decode_u_regfile_reg_r29_q_reg_26_ ( .D(u_decode_u_regfile_N1162), 
        .CK(n37833), .RN(n44116), .Q(n2623), .QN(n40889) );
  DFFRX1 u_decode_u_regfile_reg_r30_q_reg_26_ ( .D(u_decode_u_regfile_N1199), 
        .CK(n37832), .RN(n44115), .Q(n2624), .QN(n36868) );
  DFFRX1 u_decode_u_regfile_reg_r31_q_reg_26_ ( .D(u_decode_u_regfile_N1236), 
        .CK(n37831), .RN(n44116), .Q(n2625), .QN(n42480) );
  DFFRX1 u_decode_u_regfile_reg_r1_q_reg_26_ ( .D(u_decode_u_regfile_N126), 
        .CK(n37830), .RN(n44115), .Q(n2626), .QN(n37022) );
  DFFRX1 u_decode_u_regfile_reg_r2_q_reg_26_ ( .D(u_decode_u_regfile_N163), 
        .CK(n37829), .RN(n44115), .Q(n2627), .QN(n36852) );
  DFFRX1 u_decode_u_regfile_reg_r3_q_reg_26_ ( .D(u_decode_u_regfile_N200), 
        .CK(n37828), .RN(n44116), .Q(n2628), .QN(n42483) );
  DFFRX1 u_decode_u_regfile_reg_r4_q_reg_26_ ( .D(u_decode_u_regfile_N237), 
        .CK(n37827), .RN(n44115), .Q(n2629), .QN(n36846) );
  DFFRX1 u_decode_u_regfile_reg_r5_q_reg_26_ ( .D(u_decode_u_regfile_N274), 
        .CK(n37826), .RN(n44116), .Q(n2630), .QN(n36817) );
  DFFRX1 u_decode_u_regfile_reg_r6_q_reg_26_ ( .D(u_decode_u_regfile_N311), 
        .CK(n37825), .RN(n44115), .Q(n2631), .QN(n40899) );
  DFFRX1 u_decode_u_regfile_reg_r7_q_reg_26_ ( .D(u_decode_u_regfile_N348), 
        .CK(n37824), .RN(n44116), .Q(n2632), .QN(n40904) );
  DFFRX1 u_decode_u_regfile_reg_r8_q_reg_26_ ( .D(u_decode_u_regfile_N385), 
        .CK(n37823), .RN(n44115), .Q(n2633) );
  DFFRX1 u_decode_u_regfile_reg_r9_q_reg_26_ ( .D(u_decode_u_regfile_N422), 
        .CK(n37822), .RN(n44115), .Q(n2634) );
  DFFRX1 u_decode_u_regfile_reg_r10_q_reg_26_ ( .D(u_decode_u_regfile_N459), 
        .CK(n37821), .RN(n44115), .Q(n2635) );
  DFFRX1 u_decode_u_regfile_reg_r11_q_reg_26_ ( .D(u_decode_u_regfile_N496), 
        .CK(n37820), .RN(n44116), .Q(n2636), .QN(n38744) );
  DFFRX1 u_decode_u_regfile_reg_r12_q_reg_26_ ( .D(u_decode_u_regfile_N533), 
        .CK(n37819), .RN(n44115), .Q(n2637) );
  DFFRX1 u_decode_u_regfile_reg_r13_q_reg_26_ ( .D(u_decode_u_regfile_N570), 
        .CK(n37818), .RN(n44116), .Q(n2638), .QN(n40891) );
  DFFRX1 u_decode_u_regfile_reg_r14_q_reg_26_ ( .D(u_decode_u_regfile_N607), 
        .CK(n37817), .RN(n44115), .Q(n2639), .QN(n40867) );
  DFFRX1 u_decode_u_regfile_reg_r15_q_reg_26_ ( .D(u_decode_u_regfile_N644), 
        .CK(n37816), .RN(n44116), .Q(n2640) );
  DFFRX1 u_decode_u_regfile_reg_r16_q_reg_26_ ( .D(u_decode_u_regfile_N681), 
        .CK(n37815), .RN(n44114), .Q(n2641) );
  DFFRX1 u_decode_u_regfile_reg_r17_q_reg_26_ ( .D(u_decode_u_regfile_N718), 
        .CK(n37814), .RN(n44115), .Q(n2642) );
  DFFRX1 u_decode_u_regfile_reg_r18_q_reg_26_ ( .D(u_decode_u_regfile_N755), 
        .CK(n37813), .RN(n44115), .Q(n2643) );
  DFFRX1 u_decode_u_regfile_reg_r19_q_reg_26_ ( .D(u_decode_u_regfile_N792), 
        .CK(n37812), .RN(n44116), .Q(n2644) );
  DFFRX1 u_decode_u_regfile_reg_r20_q_reg_26_ ( .D(u_decode_u_regfile_N829), 
        .CK(n37811), .RN(n44115), .Q(n2645) );
  DFFRX1 u_decode_u_regfile_reg_r22_q_reg_26_ ( .D(u_decode_u_regfile_N903), 
        .CK(n37809), .RN(n44115), .Q(n2647), .QN(n40859) );
  DFFRX1 u_decode_u_regfile_reg_r23_q_reg_26_ ( .D(u_decode_u_regfile_N940), 
        .CK(n37880), .RN(n44116), .Q(n2648), .QN(n36800) );
  DFFRX1 u_lsu_mem_data_wr_q_reg_26_ ( .D(u_lsu_N220), .CK(net1847), .RN(
        n44160), .QN(n2649) );
  DFFRX1 u_lsu_mem_addr_q_reg_18_ ( .D(u_lsu_mem_addr_r[18]), .CK(n37876), 
        .RN(n44186), .Q(mmu_lsu_addr_w[18]), .QN(n8308) );
  DFFRX1 u_mmu_lsu_in_addr_q_reg_18_ ( .D(mmu_lsu_addr_w[18]), .CK(n37873), 
        .RN(n44186), .QN(n2650) );
  DFFRX1 u_mmu_itlb_va_addr_q_reg_18_ ( .D(u_mmu_virt_addr_q[18]), .CK(n37871), 
        .RN(n44186), .QN(n17102) );
  DFFRX1 u_mmu_dtlb_va_addr_q_reg_18_ ( .D(u_mmu_virt_addr_q[18]), .CK(n37872), 
        .RN(n44205), .Q(u_mmu_dtlb_va_addr_q[18]) );
  DFFRX1 u_mmu_itlb_entry_q_reg_18_ ( .D(u_mmu_pte_entry_q[18]), .CK(net1792), 
        .RN(n44171), .Q(u_mmu_itlb_entry_q[18]) );
  DFFRX1 u_mmu_dtlb_entry_q_reg_18_ ( .D(u_mmu_pte_entry_q[18]), .CK(net1782), 
        .RN(n44196), .QN(n2651) );
  DFFRX1 u_muldiv_dividend_q_reg_18_ ( .D(u_muldiv_N250), .CK(net1913), .RN(
        n44160), .Q(u_muldiv_dividend_q[18]), .QN(n37461) );
  DFFRX1 u_decode_u_regfile_reg_r25_q_reg_18_ ( .D(u_decode_u_regfile_N1006), 
        .CK(n37837), .RN(n44101), .Q(n2652), .QN(n37123) );
  DFFRX1 u_decode_u_regfile_reg_r26_q_reg_18_ ( .D(u_decode_u_regfile_N1043), 
        .CK(n37836), .RN(n44100), .Q(n2653), .QN(n36931) );
  DFFRX1 u_decode_u_regfile_reg_r27_q_reg_18_ ( .D(u_decode_u_regfile_N1080), 
        .CK(n37835), .RN(n44101), .Q(n2654), .QN(n37124) );
  DFFRX1 u_decode_u_regfile_reg_r28_q_reg_18_ ( .D(u_decode_u_regfile_N1117), 
        .CK(n37834), .RN(n44101), .Q(n2655) );
  DFFRX1 u_decode_u_regfile_reg_r29_q_reg_18_ ( .D(u_decode_u_regfile_N1154), 
        .CK(n37833), .RN(n44101), .Q(n2656), .QN(n36926) );
  DFFRX1 u_decode_u_regfile_reg_r1_q_reg_18_ ( .D(u_decode_u_regfile_N118), 
        .CK(n37830), .RN(n44101), .Q(n2657), .QN(n37128) );
  DFFRX1 u_decode_u_regfile_reg_r30_q_reg_18_ ( .D(u_decode_u_regfile_N1191), 
        .CK(n37832), .RN(n44101), .Q(n2658) );
  DFFRX1 u_decode_u_regfile_reg_r31_q_reg_18_ ( .D(u_decode_u_regfile_N1228), 
        .CK(n37831), .RN(n44102), .Q(n2659) );
  DFFRX1 u_decode_u_regfile_reg_r2_q_reg_18_ ( .D(u_decode_u_regfile_N155), 
        .CK(n37829), .RN(n44100), .Q(n2660), .QN(n36915) );
  DFFRX1 u_decode_u_regfile_reg_r3_q_reg_18_ ( .D(u_decode_u_regfile_N192), 
        .CK(n37828), .RN(n44101), .Q(n2661), .QN(n37134) );
  DFFRX1 u_decode_u_regfile_reg_r4_q_reg_18_ ( .D(u_decode_u_regfile_N229), 
        .CK(n37827), .RN(n44101), .Q(n2662), .QN(n36939) );
  DFFRX1 u_decode_u_regfile_reg_r5_q_reg_18_ ( .D(u_decode_u_regfile_N266), 
        .CK(n37826), .RN(n44101), .Q(n2663), .QN(n36917) );
  DFFRX1 u_decode_u_regfile_reg_r6_q_reg_18_ ( .D(u_decode_u_regfile_N303), 
        .CK(n37825), .RN(n44101), .Q(n2664), .QN(n36911) );
  DFFRX1 u_decode_u_regfile_reg_r7_q_reg_18_ ( .D(u_decode_u_regfile_N340), 
        .CK(n37824), .RN(n44102), .Q(n2665), .QN(n37315) );
  DFFRX1 u_decode_u_regfile_reg_r8_q_reg_18_ ( .D(u_decode_u_regfile_N377), 
        .CK(n37823), .RN(n44100), .Q(n2666), .QN(n37125) );
  DFFRX1 u_decode_u_regfile_reg_r9_q_reg_18_ ( .D(u_decode_u_regfile_N414), 
        .CK(n37822), .RN(n44101), .Q(n2667), .QN(n37129) );
  DFFRX1 u_decode_u_regfile_reg_r10_q_reg_18_ ( .D(u_decode_u_regfile_N451), 
        .CK(n37821), .RN(n44100), .Q(n2668), .QN(n36927) );
  DFFRX1 u_decode_u_regfile_reg_r11_q_reg_18_ ( .D(u_decode_u_regfile_N488), 
        .CK(n37820), .RN(n44101), .Q(n2669), .QN(n37121) );
  DFFRX1 u_decode_u_regfile_reg_r12_q_reg_18_ ( .D(u_decode_u_regfile_N525), 
        .CK(n37819), .RN(n44101), .Q(n2670), .QN(n36918) );
  DFFRX1 u_decode_u_regfile_reg_r13_q_reg_18_ ( .D(u_decode_u_regfile_N562), 
        .CK(n37818), .RN(n44101), .Q(n2671), .QN(n36919) );
  DFFRX1 u_decode_u_regfile_reg_r14_q_reg_18_ ( .D(u_decode_u_regfile_N599), 
        .CK(n37817), .RN(n44101), .Q(n2672), .QN(n36908) );
  DFFRX1 u_decode_u_regfile_reg_r15_q_reg_18_ ( .D(u_decode_u_regfile_N636), 
        .CK(n37816), .RN(n44102), .Q(n2673), .QN(n36906) );
  DFFRX1 u_decode_u_regfile_reg_r16_q_reg_18_ ( .D(u_decode_u_regfile_N673), 
        .CK(n37815), .RN(n44100), .Q(n2674), .QN(n37131) );
  DFFRX1 u_decode_u_regfile_reg_r17_q_reg_18_ ( .D(u_decode_u_regfile_N710), 
        .CK(n37814), .RN(n44101), .Q(n2675), .QN(n37135) );
  DFFRX1 u_decode_u_regfile_reg_r18_q_reg_18_ ( .D(u_decode_u_regfile_N747), 
        .CK(n37813), .RN(n44100), .Q(n2676) );
  DFFRX1 u_decode_u_regfile_reg_r19_q_reg_18_ ( .D(u_decode_u_regfile_N784), 
        .CK(n37812), .RN(n44101), .Q(n2677), .QN(n37132) );
  DFFRX1 u_decode_u_regfile_reg_r20_q_reg_18_ ( .D(u_decode_u_regfile_N821), 
        .CK(n37811), .RN(n44100), .Q(n2678) );
  DFFRX1 u_decode_u_regfile_reg_r21_q_reg_18_ ( .D(u_decode_u_regfile_N858), 
        .CK(n37810), .RN(n44102), .Q(n2679) );
  DFFRX1 u_decode_u_regfile_reg_r22_q_reg_18_ ( .D(u_decode_u_regfile_N895), 
        .CK(n37809), .RN(n44101), .Q(n2680) );
  DFFRX1 u_decode_u_regfile_reg_r23_q_reg_18_ ( .D(u_decode_u_regfile_N932), 
        .CK(n37880), .RN(n44102), .Q(n2681), .QN(n36912) );
  DFFRX1 u_lsu_mem_data_wr_q_reg_18_ ( .D(u_lsu_N212), .CK(net1847), .RN(
        n44159), .QN(n2682) );
  DFFRX1 u_lsu_mem_addr_q_reg_12_ ( .D(u_lsu_mem_addr_r[12]), .CK(n37869), 
        .RN(n44185), .Q(mmu_lsu_addr_w[12]), .QN(n8296) );
  DFFRX1 u_mmu_lsu_in_addr_q_reg_12_ ( .D(mmu_lsu_addr_w[12]), .CK(n37875), 
        .RN(n44185), .QN(n2683) );
  DFFRX1 u_mmu_itlb_va_addr_q_reg_12_ ( .D(u_mmu_virt_addr_q[12]), .CK(n37871), 
        .RN(n44185), .Q(n2684) );
  DFFRX1 u_mmu_dtlb_va_addr_q_reg_12_ ( .D(u_mmu_virt_addr_q[12]), .CK(n37872), 
        .RN(n44205), .Q(u_mmu_dtlb_va_addr_q[12]) );
  DFFRX1 u_mmu_itlb_entry_q_reg_12_ ( .D(u_mmu_pte_entry_q[12]), .CK(net1792), 
        .RN(n44171), .Q(u_mmu_itlb_entry_q[12]) );
  DFFRX1 u_mmu_dtlb_entry_q_reg_12_ ( .D(u_mmu_pte_entry_q[12]), .CK(net1782), 
        .RN(n44210), .QN(n2685) );
  DFFRX1 u_muldiv_dividend_q_reg_12_ ( .D(u_muldiv_N244), .CK(net1908), .RN(
        n44159), .Q(u_muldiv_dividend_q[12]), .QN(n37441) );
  DFFRX1 u_decode_u_regfile_reg_r25_q_reg_12_ ( .D(u_decode_u_regfile_N1000), 
        .CK(n37879), .RN(n44139), .Q(n2686), .QN(n37210) );
  DFFRX1 u_decode_u_regfile_reg_r26_q_reg_12_ ( .D(u_decode_u_regfile_N1037), 
        .CK(n37864), .RN(n44138), .Q(n2687) );
  DFFRX1 u_decode_u_regfile_reg_r27_q_reg_12_ ( .D(u_decode_u_regfile_N1074), 
        .CK(n37863), .RN(n44139), .Q(n2688) );
  DFFRX1 u_decode_u_regfile_reg_r28_q_reg_12_ ( .D(u_decode_u_regfile_N1111), 
        .CK(n37862), .RN(n44138), .Q(n2689), .QN(n36937) );
  DFFRX1 u_decode_u_regfile_reg_r1_q_reg_12_ ( .D(u_decode_u_regfile_N112), 
        .CK(n37865), .RN(n44139), .Q(n2690), .QN(n37215) );
  DFFRX1 u_decode_u_regfile_reg_r29_q_reg_12_ ( .D(u_decode_u_regfile_N1148), 
        .CK(n37861), .RN(n44139), .Q(n2691) );
  DFFRX1 u_decode_u_regfile_reg_r30_q_reg_12_ ( .D(u_decode_u_regfile_N1185), 
        .CK(n37860), .RN(n44139), .Q(n2692), .QN(n36920) );
  DFFRX1 u_decode_u_regfile_reg_r31_q_reg_12_ ( .D(u_decode_u_regfile_N1222), 
        .CK(n37859), .RN(n44140), .Q(n2693), .QN(n36921) );
  DFFRX1 u_decode_u_regfile_reg_r2_q_reg_12_ ( .D(u_decode_u_regfile_N149), 
        .CK(n37858), .RN(n44138), .Q(n2694) );
  DFFRX1 u_decode_u_regfile_reg_r3_q_reg_12_ ( .D(u_decode_u_regfile_N186), 
        .CK(n37857), .RN(n44139), .Q(n2695), .QN(n37199) );
  DFFRX1 u_decode_u_regfile_reg_r4_q_reg_12_ ( .D(u_decode_u_regfile_N223), 
        .CK(n37856), .RN(n44138), .Q(n2696) );
  DFFRX1 u_decode_u_regfile_reg_r5_q_reg_12_ ( .D(u_decode_u_regfile_N260), 
        .CK(n37840), .RN(n44139), .Q(n2697) );
  DFFRX1 u_decode_u_regfile_reg_r6_q_reg_12_ ( .D(u_decode_u_regfile_N297), 
        .CK(n37855), .RN(n44139), .Q(n2698) );
  DFFRX1 u_decode_u_regfile_reg_r7_q_reg_12_ ( .D(u_decode_u_regfile_N334), 
        .CK(n37854), .RN(n44140), .QN(n36928) );
  DFFRX1 u_decode_u_regfile_reg_r8_q_reg_12_ ( .D(u_decode_u_regfile_N371), 
        .CK(n37839), .RN(n44138), .Q(n2700), .QN(n37197) );
  DFFRX1 u_decode_u_regfile_reg_r9_q_reg_12_ ( .D(u_decode_u_regfile_N408), 
        .CK(n37853), .RN(n44139), .Q(n2701), .QN(n37203) );
  DFFRX1 u_decode_u_regfile_reg_r10_q_reg_12_ ( .D(u_decode_u_regfile_N445), 
        .CK(n37852), .RN(n44138), .Q(n2702) );
  DFFRX1 u_decode_u_regfile_reg_r11_q_reg_12_ ( .D(u_decode_u_regfile_N482), 
        .CK(n37851), .RN(n44139), .Q(n2703), .QN(n37205) );
  DFFRX1 u_decode_u_regfile_reg_r12_q_reg_12_ ( .D(u_decode_u_regfile_N519), 
        .CK(n37850), .RN(n44138), .Q(n2704) );
  DFFRX1 u_decode_u_regfile_reg_r13_q_reg_12_ ( .D(u_decode_u_regfile_N556), 
        .CK(n37849), .RN(n44139), .Q(n2705) );
  DFFRX1 u_decode_u_regfile_reg_r14_q_reg_12_ ( .D(u_decode_u_regfile_N593), 
        .CK(n37848), .RN(n44139), .Q(n2706) );
  DFFRX1 u_decode_u_regfile_reg_r15_q_reg_12_ ( .D(u_decode_u_regfile_N630), 
        .CK(n37847), .RN(n44139), .Q(n2707) );
  DFFRX1 u_decode_u_regfile_reg_r16_q_reg_12_ ( .D(u_decode_u_regfile_N667), 
        .CK(n37846), .RN(n44138), .Q(n2708), .QN(n37204) );
  DFFRX1 u_decode_u_regfile_reg_r17_q_reg_12_ ( .D(u_decode_u_regfile_N704), 
        .CK(n37845), .RN(n44139), .Q(n2709), .QN(n37206) );
  DFFRX1 u_decode_u_regfile_reg_r18_q_reg_12_ ( .D(u_decode_u_regfile_N741), 
        .CK(n37844), .RN(n44138), .Q(n2710), .QN(n36930) );
  DFFRX1 u_decode_u_regfile_reg_r19_q_reg_12_ ( .D(u_decode_u_regfile_N778), 
        .CK(n37843), .RN(n44139), .Q(n2711), .QN(n37194) );
  DFFRX1 u_decode_u_regfile_reg_r20_q_reg_12_ ( .D(u_decode_u_regfile_N815), 
        .CK(n37842), .RN(n44138), .Q(n2712), .QN(n36924) );
  DFFRX1 u_decode_u_regfile_reg_r21_q_reg_12_ ( .D(u_decode_u_regfile_N852), 
        .CK(n37838), .RN(n44139), .Q(n2713), .QN(n36929) );
  DFFRX1 u_decode_u_regfile_reg_r22_q_reg_12_ ( .D(u_decode_u_regfile_N889), 
        .CK(n37841), .RN(n44139), .Q(n2714), .QN(n36914) );
  DFFRX1 u_decode_u_regfile_reg_r23_q_reg_12_ ( .D(u_decode_u_regfile_N926), 
        .CK(n37877), .RN(n44139), .Q(n2715) );
  DFFRX1 u_lsu_mem_addr_q_reg_8_ ( .D(u_lsu_mem_addr_r[8]), .CK(n37869), .RN(
        n44199), .Q(mmu_lsu_addr_w[8]), .QN(n2716) );
  DFFRX1 u_mmu_lsu_in_addr_q_reg_8_ ( .D(mmu_lsu_addr_w[8]), .CK(n37875), .RN(
        n44199), .QN(n2717) );
  DFFRX1 u_muldiv_dividend_q_reg_8_ ( .D(u_muldiv_N240), .CK(net1908), .RN(
        n44159), .Q(u_muldiv_dividend_q[8]), .QN(n37428) );
  DFFRX1 u_decode_u_regfile_reg_r26_q_reg_8_ ( .D(u_decode_u_regfile_N1033), 
        .CK(n37864), .RN(n44126), .Q(n2718), .QN(n42514) );
  DFFRX1 u_decode_u_regfile_reg_r27_q_reg_8_ ( .D(u_decode_u_regfile_N1070), 
        .CK(n37863), .RN(n44127), .Q(n2719) );
  DFFRX1 u_decode_u_regfile_reg_r1_q_reg_8_ ( .D(u_decode_u_regfile_N108), 
        .CK(n37865), .RN(n44127), .Q(n2720), .QN(n37250) );
  DFFRX1 u_decode_u_regfile_reg_r28_q_reg_8_ ( .D(u_decode_u_regfile_N1107), 
        .CK(n37862), .RN(n44126), .Q(n2721), .QN(n37072) );
  DFFRX1 u_decode_u_regfile_reg_r29_q_reg_8_ ( .D(u_decode_u_regfile_N1144), 
        .CK(n37861), .RN(n44127), .Q(n2722) );
  DFFRX1 u_decode_u_regfile_reg_r30_q_reg_8_ ( .D(u_decode_u_regfile_N1181), 
        .CK(n37860), .RN(n44126), .Q(n2723), .QN(n37056) );
  DFFRX1 u_decode_u_regfile_reg_r31_q_reg_8_ ( .D(u_decode_u_regfile_N1218), 
        .CK(n37859), .RN(n44127), .Q(n2724), .QN(n37058) );
  DFFRX1 u_decode_u_regfile_reg_r2_q_reg_8_ ( .D(u_decode_u_regfile_N145), 
        .CK(n37858), .RN(n44126), .Q(n2725) );
  DFFRX1 u_decode_u_regfile_reg_r3_q_reg_8_ ( .D(u_decode_u_regfile_N182), 
        .CK(n37857), .RN(n44127), .Q(n2726), .QN(n37243) );
  DFFRX1 u_decode_u_regfile_reg_r4_q_reg_8_ ( .D(u_decode_u_regfile_N219), 
        .CK(n37856), .RN(n44126), .Q(n2727) );
  DFFRX1 u_decode_u_regfile_reg_r5_q_reg_8_ ( .D(u_decode_u_regfile_N256), 
        .CK(n37840), .RN(n44127), .Q(n2728) );
  DFFRX1 u_decode_u_regfile_reg_r6_q_reg_8_ ( .D(u_decode_u_regfile_N293), 
        .CK(n37855), .RN(n44126), .Q(n2729) );
  DFFRX1 u_decode_u_regfile_reg_r7_q_reg_8_ ( .D(u_decode_u_regfile_N330), 
        .CK(n37854), .RN(n44127), .QN(n37066) );
  DFFRX1 u_decode_u_regfile_reg_r8_q_reg_8_ ( .D(u_decode_u_regfile_N367), 
        .CK(n37839), .RN(n44126), .Q(n2731), .QN(n37242) );
  DFFRX1 u_decode_u_regfile_reg_r9_q_reg_8_ ( .D(u_decode_u_regfile_N404), 
        .CK(n37853), .RN(n44127), .Q(n2732), .QN(n37246) );
  DFFRX1 u_decode_u_regfile_reg_r10_q_reg_8_ ( .D(u_decode_u_regfile_N441), 
        .CK(n37852), .RN(n44126), .Q(n2733) );
  DFFRX1 u_decode_u_regfile_reg_r11_q_reg_8_ ( .D(u_decode_u_regfile_N478), 
        .CK(n37851), .RN(n44127), .Q(n2734), .QN(n37244) );
  DFFRX1 u_decode_u_regfile_reg_r12_q_reg_8_ ( .D(u_decode_u_regfile_N515), 
        .CK(n37850), .RN(n44126), .Q(n2735) );
  DFFRX1 u_decode_u_regfile_reg_r13_q_reg_8_ ( .D(u_decode_u_regfile_N552), 
        .CK(n37849), .RN(n44127), .Q(n2736) );
  DFFRX1 u_decode_u_regfile_reg_r14_q_reg_8_ ( .D(u_decode_u_regfile_N589), 
        .CK(n37848), .RN(n44126), .Q(n2737) );
  DFFRX1 u_decode_u_regfile_reg_r15_q_reg_8_ ( .D(u_decode_u_regfile_N626), 
        .CK(n37847), .RN(n44127), .Q(n2738) );
  DFFRX1 u_decode_u_regfile_reg_r16_q_reg_8_ ( .D(u_decode_u_regfile_N663), 
        .CK(n37846), .RN(n44126), .Q(n2739), .QN(n37245) );
  DFFRX1 u_decode_u_regfile_reg_r17_q_reg_8_ ( .D(u_decode_u_regfile_N700), 
        .CK(n37845), .RN(n44127), .Q(n2740), .QN(n37248) );
  DFFRX1 u_decode_u_regfile_reg_r18_q_reg_8_ ( .D(u_decode_u_regfile_N737), 
        .CK(n37844), .RN(n44126), .Q(n2741), .QN(n37065) );
  DFFRX1 u_decode_u_regfile_reg_r19_q_reg_8_ ( .D(u_decode_u_regfile_N774), 
        .CK(n37843), .RN(n44127), .Q(n2742), .QN(n37241) );
  DFFRX1 u_decode_u_regfile_reg_r20_q_reg_8_ ( .D(u_decode_u_regfile_N811), 
        .CK(n37842), .RN(n44126), .Q(n2743), .QN(n37059) );
  DFFRX1 u_decode_u_regfile_reg_r21_q_reg_8_ ( .D(u_decode_u_regfile_N848), 
        .CK(n37838), .RN(n44127), .Q(n2744), .QN(n37063) );
  DFFRX1 u_decode_u_regfile_reg_r22_q_reg_8_ ( .D(u_decode_u_regfile_N885), 
        .CK(n37841), .RN(n44126), .Q(n2745), .QN(n37049) );
  DFFRX1 u_decode_u_regfile_reg_r23_q_reg_8_ ( .D(u_decode_u_regfile_N922), 
        .CK(n37877), .RN(n44127), .Q(n2746) );
  DFFRX1 u_decode_u_regfile_reg_r24_q_reg_8_ ( .D(u_decode_u_regfile_N959), 
        .CK(n37878), .RN(n44126), .Q(n2747), .QN(n37249) );
  DFFRX1 u_lsu_mem_data_wr_q_reg_4_ ( .D(u_lsu_N198), .CK(n37874), .RN(n44200), 
        .QN(n2748) );
  DFFRX1 u_lsu_mem_data_wr_q_reg_12_ ( .D(u_lsu_N206), .CK(n37874), .RN(n44159), .QN(n2749) );
  DFFRX1 u_lsu_mem_data_wr_q_reg_20_ ( .D(u_lsu_N214), .CK(net1847), .RN(
        n44159), .QN(n2750) );
  DFFRX1 u_lsu_mem_data_wr_q_reg_1_ ( .D(u_lsu_N195), .CK(n37874), .RN(n44200), 
        .QN(n2751) );
  DFFRX1 u_lsu_mem_data_wr_q_reg_9_ ( .D(u_lsu_N203), .CK(n37874), .RN(n44159), 
        .QN(n2752) );
  DFFRX1 u_lsu_mem_addr_q_reg_13_ ( .D(u_lsu_mem_addr_r[13]), .CK(n37876), 
        .RN(n44186), .Q(mmu_lsu_addr_w[13]), .QN(n8298) );
  DFFRX1 u_mmu_lsu_in_addr_q_reg_13_ ( .D(mmu_lsu_addr_w[13]), .CK(n37875), 
        .RN(n44186), .QN(n2753) );
  DFFRX1 u_mmu_itlb_va_addr_q_reg_13_ ( .D(u_mmu_virt_addr_q[13]), .CK(n37871), 
        .RN(n44186), .QN(n16237) );
  DFFRX1 u_mmu_dtlb_va_addr_q_reg_13_ ( .D(u_mmu_virt_addr_q[13]), .CK(n37872), 
        .RN(n44206), .Q(u_mmu_dtlb_va_addr_q[13]) );
  DFFRX1 u_mmu_itlb_entry_q_reg_13_ ( .D(u_mmu_pte_entry_q[13]), .CK(net1792), 
        .RN(n44171), .Q(u_mmu_itlb_entry_q[13]) );
  DFFRX1 u_mmu_dtlb_entry_q_reg_13_ ( .D(u_mmu_pte_entry_q[13]), .CK(net1782), 
        .RN(n44210), .QN(n2754) );
  DFFRX1 u_muldiv_dividend_q_reg_13_ ( .D(u_muldiv_N245), .CK(net1908), .RN(
        n44159), .Q(u_muldiv_dividend_q[13]) );
  DFFRX1 u_decode_u_regfile_reg_r25_q_reg_13_ ( .D(u_decode_u_regfile_N1001), 
        .CK(n37879), .RN(n44122), .Q(n2755), .QN(n37190) );
  DFFRX1 u_decode_u_regfile_reg_r26_q_reg_13_ ( .D(u_decode_u_regfile_N1038), 
        .CK(n37864), .RN(n44122), .Q(n2756) );
  DFFRX1 u_decode_u_regfile_reg_r27_q_reg_13_ ( .D(u_decode_u_regfile_N1075), 
        .CK(n37863), .RN(n44123), .Q(n2757) );
  DFFRX1 u_decode_u_regfile_reg_r28_q_reg_13_ ( .D(u_decode_u_regfile_N1112), 
        .CK(n37862), .RN(n44122), .Q(n2758), .QN(n36861) );
  DFFRX1 u_decode_u_regfile_reg_r1_q_reg_13_ ( .D(u_decode_u_regfile_N113), 
        .CK(n37865), .RN(n44122), .Q(n2759), .QN(n37193) );
  DFFRX1 u_decode_u_regfile_reg_r29_q_reg_13_ ( .D(u_decode_u_regfile_N1149), 
        .CK(n37861), .RN(n44123), .Q(n2760) );
  DFFRX1 u_decode_u_regfile_reg_r30_q_reg_13_ ( .D(u_decode_u_regfile_N1186), 
        .CK(n37860), .RN(n44122), .Q(n2761), .QN(n36850) );
  DFFRX1 u_decode_u_regfile_reg_r31_q_reg_13_ ( .D(u_decode_u_regfile_N1223), 
        .CK(n37859), .RN(n44123), .Q(n2762), .QN(n36844) );
  DFFRX1 u_decode_u_regfile_reg_r2_q_reg_13_ ( .D(u_decode_u_regfile_N150), 
        .CK(n37858), .RN(n44122), .Q(n2763) );
  DFFRX1 u_decode_u_regfile_reg_r3_q_reg_13_ ( .D(u_decode_u_regfile_N187), 
        .CK(n37857), .RN(n44123), .Q(n2764), .QN(n37183) );
  DFFRX1 u_decode_u_regfile_reg_r4_q_reg_13_ ( .D(u_decode_u_regfile_N224), 
        .CK(n37856), .RN(n44122), .Q(n2765) );
  DFFRX1 u_decode_u_regfile_reg_r5_q_reg_13_ ( .D(u_decode_u_regfile_N261), 
        .CK(n37840), .RN(n44123), .Q(n2766) );
  DFFRX1 u_decode_u_regfile_reg_r6_q_reg_13_ ( .D(u_decode_u_regfile_N298), 
        .CK(n37855), .RN(n44122), .Q(n2767) );
  DFFRX1 u_decode_u_regfile_reg_r7_q_reg_13_ ( .D(u_decode_u_regfile_N335), 
        .CK(n37854), .RN(n44123), .QN(n36853) );
  DFFRX1 u_decode_u_regfile_reg_r8_q_reg_13_ ( .D(u_decode_u_regfile_N372), 
        .CK(n37839), .RN(n44122), .Q(n2769), .QN(n37184) );
  DFFRX1 u_decode_u_regfile_reg_r9_q_reg_13_ ( .D(u_decode_u_regfile_N409), 
        .CK(n37853), .RN(n44122), .Q(n2770), .QN(n37186) );
  DFFRX1 u_decode_u_regfile_reg_r10_q_reg_13_ ( .D(u_decode_u_regfile_N446), 
        .CK(n37852), .RN(n44122), .Q(n2771) );
  DFFRX1 u_decode_u_regfile_reg_r11_q_reg_13_ ( .D(u_decode_u_regfile_N483), 
        .CK(n37851), .RN(n44123), .Q(n2772), .QN(n37187) );
  DFFRX1 u_decode_u_regfile_reg_r12_q_reg_13_ ( .D(u_decode_u_regfile_N520), 
        .CK(n37850), .RN(n44122), .Q(n2773) );
  DFFRX1 u_decode_u_regfile_reg_r13_q_reg_13_ ( .D(u_decode_u_regfile_N557), 
        .CK(n37849), .RN(n44123), .Q(n2774) );
  DFFRX1 u_decode_u_regfile_reg_r14_q_reg_13_ ( .D(u_decode_u_regfile_N594), 
        .CK(n37848), .RN(n44122), .Q(n2775) );
  DFFRX1 u_decode_u_regfile_reg_r15_q_reg_13_ ( .D(u_decode_u_regfile_N631), 
        .CK(n37847), .RN(n44123), .Q(n2776) );
  DFFRX1 u_decode_u_regfile_reg_r16_q_reg_13_ ( .D(u_decode_u_regfile_N668), 
        .CK(n37846), .RN(n44122), .Q(n2777), .QN(n37185) );
  DFFRX1 u_decode_u_regfile_reg_r17_q_reg_13_ ( .D(u_decode_u_regfile_N705), 
        .CK(n37845), .RN(n44123), .Q(n2778), .QN(n37189) );
  DFFRX1 u_decode_u_regfile_reg_r18_q_reg_13_ ( .D(u_decode_u_regfile_N742), 
        .CK(n37844), .RN(n44122), .Q(n2779), .QN(n36856) );
  DFFRX1 u_decode_u_regfile_reg_r19_q_reg_13_ ( .D(u_decode_u_regfile_N779), 
        .CK(n37843), .RN(n44123), .Q(n2780), .QN(n37182) );
  DFFRX1 u_decode_u_regfile_reg_r20_q_reg_13_ ( .D(u_decode_u_regfile_N816), 
        .CK(n37842), .RN(n44122), .Q(n2781), .QN(n36849) );
  DFFRX1 u_decode_u_regfile_reg_r21_q_reg_13_ ( .D(u_decode_u_regfile_N853), 
        .CK(n37838), .RN(n44123), .Q(n2782), .QN(n36855) );
  DFFRX1 u_decode_u_regfile_reg_r22_q_reg_13_ ( .D(u_decode_u_regfile_N890), 
        .CK(n37841), .RN(n44122), .Q(n2783), .QN(n36838) );
  DFFRX1 u_decode_u_regfile_reg_r23_q_reg_13_ ( .D(u_decode_u_regfile_N927), 
        .CK(n37877), .RN(n44123), .Q(n2784), .QN(n38666) );
  DFFRX1 u_lsu_mem_addr_q_reg_27_ ( .D(u_lsu_mem_addr_r[27]), .CK(n37876), 
        .RN(n44183), .Q(mmu_lsu_addr_w[27]), .QN(n8328) );
  DFFRX1 u_mmu_lsu_in_addr_q_reg_27_ ( .D(mmu_lsu_addr_w[27]), .CK(n37873), 
        .RN(n44183), .QN(n2785) );
  DFFRX1 u_decode_u_regfile_reg_r25_q_reg_27_ ( .D(u_decode_u_regfile_N1015), 
        .CK(n37837), .RN(n44190), .Q(n2786), .QN(n37020) );
  DFFRX1 u_decode_u_regfile_reg_r26_q_reg_27_ ( .D(u_decode_u_regfile_N1052), 
        .CK(n37836), .RN(n44189), .Q(n2787), .QN(n38716) );
  DFFRX1 u_decode_u_regfile_reg_r27_q_reg_27_ ( .D(u_decode_u_regfile_N1089), 
        .CK(n37835), .RN(n44190), .Q(n2788), .QN(n37027) );
  DFFRX1 u_decode_u_regfile_reg_r28_q_reg_27_ ( .D(u_decode_u_regfile_N1126), 
        .CK(n37834), .RN(n44189), .Q(n2789) );
  DFFRX1 u_decode_u_regfile_reg_r29_q_reg_27_ ( .D(u_decode_u_regfile_N1163), 
        .CK(n37833), .RN(n44190), .Q(n2790), .QN(n36842) );
  DFFRX1 u_decode_u_regfile_reg_r30_q_reg_27_ ( .D(u_decode_u_regfile_N1200), 
        .CK(n37832), .RN(n44190), .Q(n2791), .QN(n36837) );
  DFFRX1 u_decode_u_regfile_reg_r31_q_reg_27_ ( .D(u_decode_u_regfile_N1237), 
        .CK(n37831), .RN(n44191), .Q(n2792), .QN(n36836) );
  DFFRX1 u_decode_u_regfile_reg_r1_q_reg_27_ ( .D(u_decode_u_regfile_N127), 
        .CK(n37830), .RN(n44190), .Q(n2793), .QN(n37021) );
  DFFRX1 u_decode_u_regfile_reg_r2_q_reg_27_ ( .D(u_decode_u_regfile_N164), 
        .CK(n37829), .RN(n44189), .Q(n2794), .QN(n36798) );
  DFFRX1 u_decode_u_regfile_reg_r3_q_reg_27_ ( .D(u_decode_u_regfile_N201), 
        .CK(n37828), .RN(n44190), .Q(n2795), .QN(n37036) );
  DFFRX1 u_decode_u_regfile_reg_r4_q_reg_27_ ( .D(u_decode_u_regfile_N238), 
        .CK(n37827), .RN(n44189), .Q(n2796), .QN(n36840) );
  DFFRX1 u_decode_u_regfile_reg_r5_q_reg_27_ ( .D(u_decode_u_regfile_N275), 
        .CK(n37826), .RN(n44190), .Q(n2797), .QN(n36845) );
  DFFRX1 u_decode_u_regfile_reg_r6_q_reg_27_ ( .D(u_decode_u_regfile_N312), 
        .CK(n37825), .RN(n44190), .Q(n2798), .QN(n36851) );
  DFFRX1 u_decode_u_regfile_reg_r7_q_reg_27_ ( .D(u_decode_u_regfile_N349), 
        .CK(n37824), .RN(n44191), .Q(n2799), .QN(n37323) );
  DFFRX1 u_decode_u_regfile_reg_r8_q_reg_27_ ( .D(u_decode_u_regfile_N386), 
        .CK(n37823), .RN(n44189), .Q(n2800), .QN(n37033) );
  DFFRX1 u_decode_u_regfile_reg_r9_q_reg_27_ ( .D(u_decode_u_regfile_N423), 
        .CK(n37822), .RN(n44190), .Q(n2801), .QN(n37023) );
  DFFRX1 u_decode_u_regfile_reg_r10_q_reg_27_ ( .D(u_decode_u_regfile_N460), 
        .CK(n37821), .RN(n44189), .Q(n2802) );
  DFFRX1 u_decode_u_regfile_reg_r11_q_reg_27_ ( .D(u_decode_u_regfile_N497), 
        .CK(n37820), .RN(n44190), .Q(n2803), .QN(n37064) );
  DFFRX1 u_decode_u_regfile_reg_r12_q_reg_27_ ( .D(u_decode_u_regfile_N534), 
        .CK(n37819), .RN(n44189), .Q(n2804), .QN(n42532) );
  DFFRX1 u_decode_u_regfile_reg_r13_q_reg_27_ ( .D(u_decode_u_regfile_N571), 
        .CK(n37818), .RN(n44190), .Q(n2805), .QN(n42529) );
  DFFRX1 u_decode_u_regfile_reg_r14_q_reg_27_ ( .D(u_decode_u_regfile_N608), 
        .CK(n37817), .RN(n44190), .Q(n2806), .QN(n36839) );
  DFFRX1 u_decode_u_regfile_reg_r15_q_reg_27_ ( .D(u_decode_u_regfile_N645), 
        .CK(n37816), .RN(n44190), .Q(n2807), .QN(n42531) );
  DFFRX1 u_decode_u_regfile_reg_r16_q_reg_27_ ( .D(u_decode_u_regfile_N682), 
        .CK(n37815), .RN(n44189), .Q(n2808), .QN(n42528) );
  DFFRX1 u_decode_u_regfile_reg_r17_q_reg_27_ ( .D(u_decode_u_regfile_N719), 
        .CK(n37814), .RN(n44190), .Q(n2809), .QN(n37019) );
  DFFRX1 u_decode_u_regfile_reg_r18_q_reg_27_ ( .D(u_decode_u_regfile_N756), 
        .CK(n37813), .RN(n44189), .Q(n2810) );
  DFFRX1 u_decode_u_regfile_reg_r19_q_reg_27_ ( .D(u_decode_u_regfile_N793), 
        .CK(n37812), .RN(n44190), .Q(n2811), .QN(n37025) );
  DFFRX1 u_decode_u_regfile_reg_r20_q_reg_27_ ( .D(u_decode_u_regfile_N830), 
        .CK(n37811), .RN(n44189), .Q(n2812) );
  DFFRX1 u_decode_u_regfile_reg_r21_q_reg_27_ ( .D(u_decode_u_regfile_N867), 
        .CK(n37810), .RN(n44190), .Q(n2813), .QN(n42530) );
  DFFRX1 u_decode_u_regfile_reg_r22_q_reg_27_ ( .D(u_decode_u_regfile_N904), 
        .CK(n37809), .RN(n44190), .Q(n2814) );
  DFFRX1 u_decode_u_regfile_reg_r23_q_reg_27_ ( .D(u_decode_u_regfile_N941), 
        .CK(n37880), .RN(n44190), .Q(n2815) );
  DFFRX1 u_lsu_mem_data_wr_q_reg_27_ ( .D(u_lsu_N221), .CK(net1847), .RN(
        n44159), .QN(n2816) );
  DFFRX1 u_lsu_mem_addr_q_reg_25_ ( .D(u_lsu_mem_addr_r[25]), .CK(n37876), 
        .RN(n44183), .Q(mmu_lsu_addr_w[25]), .QN(n8324) );
  DFFRX1 u_mmu_lsu_in_addr_q_reg_25_ ( .D(mmu_lsu_addr_w[25]), .CK(n37873), 
        .RN(n44183), .QN(n2817) );
  DFFRX1 u_mmu_itlb_va_addr_q_reg_25_ ( .D(n8431), .CK(clk_i), .RN(n44183), 
        .Q(u_mmu_itlb_va_addr_q[25]) );
  DFFRX1 u_mmu_dtlb_va_addr_q_reg_25_ ( .D(n8430), .CK(clk_i), .RN(n44206), 
        .Q(u_mmu_dtlb_va_addr_q[25]) );
  DFFRX1 u_decode_u_regfile_reg_r25_q_reg_25_ ( .D(u_decode_u_regfile_N1013), 
        .CK(n37837), .RN(n44113), .Q(n2819), .QN(n37018) );
  DFFRX1 u_decode_u_regfile_reg_r26_q_reg_25_ ( .D(u_decode_u_regfile_N1050), 
        .CK(n37836), .RN(n44113), .Q(n2820) );
  DFFRX1 u_decode_u_regfile_reg_r27_q_reg_25_ ( .D(u_decode_u_regfile_N1087), 
        .CK(n37835), .RN(n44114), .Q(n2821) );
  DFFRX1 u_decode_u_regfile_reg_r28_q_reg_25_ ( .D(u_decode_u_regfile_N1124), 
        .CK(n37834), .RN(n44113), .Q(n2822), .QN(n42491) );
  DFFRX1 u_decode_u_regfile_reg_r29_q_reg_25_ ( .D(u_decode_u_regfile_N1161), 
        .CK(n37833), .RN(n44114), .Q(n2823), .QN(n42506) );
  DFFRX1 u_decode_u_regfile_reg_r30_q_reg_25_ ( .D(u_decode_u_regfile_N1198), 
        .CK(n37832), .RN(n44113), .Q(n2824), .QN(n36831) );
  DFFRX1 u_decode_u_regfile_reg_r31_q_reg_25_ ( .D(u_decode_u_regfile_N1235), 
        .CK(n37831), .RN(n44114), .Q(n2825), .QN(n36830) );
  DFFRX1 u_decode_u_regfile_reg_r1_q_reg_25_ ( .D(u_decode_u_regfile_N125), 
        .CK(n37830), .RN(n44114), .Q(n2826) );
  DFFRX1 u_decode_u_regfile_reg_r2_q_reg_25_ ( .D(u_decode_u_regfile_N162), 
        .CK(n37829), .RN(n44113), .Q(n2827) );
  DFFRX1 u_decode_u_regfile_reg_r3_q_reg_25_ ( .D(u_decode_u_regfile_N199), 
        .CK(n37828), .RN(n44114), .Q(n2828) );
  DFFRX1 u_decode_u_regfile_reg_r4_q_reg_25_ ( .D(u_decode_u_regfile_N236), 
        .CK(n37827), .RN(n44113), .Q(n2829) );
  DFFRX1 u_decode_u_regfile_reg_r5_q_reg_25_ ( .D(u_decode_u_regfile_N273), 
        .CK(n37826), .RN(n44114), .Q(n2830), .QN(n42508) );
  DFFRX1 u_decode_u_regfile_reg_r6_q_reg_25_ ( .D(u_decode_u_regfile_N310), 
        .CK(n37825), .RN(n44113), .Q(n2831), .QN(n36835) );
  DFFRX1 u_decode_u_regfile_reg_r7_q_reg_25_ ( .D(u_decode_u_regfile_N347), 
        .CK(n37824), .RN(n44114), .Q(n2832), .QN(n37322) );
  DFFRX1 u_decode_u_regfile_reg_r8_q_reg_25_ ( .D(u_decode_u_regfile_N384), 
        .CK(n37823), .RN(n44113), .Q(n2833), .QN(n38743) );
  DFFRX1 u_decode_u_regfile_reg_r9_q_reg_25_ ( .D(u_decode_u_regfile_N421), 
        .CK(n37822), .RN(n44114), .Q(n2834) );
  DFFRX1 u_decode_u_regfile_reg_r10_q_reg_25_ ( .D(u_decode_u_regfile_N458), 
        .CK(n37821), .RN(n44113), .Q(n2835) );
  DFFRX1 u_decode_u_regfile_reg_r11_q_reg_25_ ( .D(u_decode_u_regfile_N495), 
        .CK(n37820), .RN(n44114), .Q(n2836) );
  DFFRX1 u_decode_u_regfile_reg_r12_q_reg_25_ ( .D(u_decode_u_regfile_N532), 
        .CK(n37819), .RN(n44113), .Q(n2837) );
  DFFRX1 u_decode_u_regfile_reg_r13_q_reg_25_ ( .D(u_decode_u_regfile_N569), 
        .CK(n37818), .RN(n44114), .Q(n2838) );
  DFFRX1 u_decode_u_regfile_reg_r14_q_reg_25_ ( .D(u_decode_u_regfile_N606), 
        .CK(n37817), .RN(n44113), .Q(n2839), .QN(n36816) );
  DFFRX1 u_decode_u_regfile_reg_r15_q_reg_25_ ( .D(u_decode_u_regfile_N643), 
        .CK(n37816), .RN(n44114), .Q(n2840), .QN(n36833) );
  DFFRX1 u_decode_u_regfile_reg_r16_q_reg_25_ ( .D(u_decode_u_regfile_N680), 
        .CK(n37815), .RN(n44113), .Q(n2841) );
  DFFRX1 u_decode_u_regfile_reg_r17_q_reg_25_ ( .D(u_decode_u_regfile_N717), 
        .CK(n37814), .RN(n44114), .Q(n2842), .QN(n37017) );
  DFFRX1 u_decode_u_regfile_reg_r18_q_reg_25_ ( .D(u_decode_u_regfile_N754), 
        .CK(n37813), .RN(n44113), .Q(n2843) );
  DFFRX1 u_decode_u_regfile_reg_r19_q_reg_25_ ( .D(u_decode_u_regfile_N791), 
        .CK(n37812), .RN(n44114), .Q(n2844), .QN(n37071) );
  DFFRX1 u_decode_u_regfile_reg_r20_q_reg_25_ ( .D(u_decode_u_regfile_N828), 
        .CK(n37811), .RN(n44113), .Q(n2845) );
  DFFRX1 u_decode_u_regfile_reg_r21_q_reg_25_ ( .D(u_decode_u_regfile_N865), 
        .CK(n37810), .RN(n44114), .Q(n2846) );
  DFFRX1 u_decode_u_regfile_reg_r22_q_reg_25_ ( .D(u_decode_u_regfile_N902), 
        .CK(n37809), .RN(n44113), .Q(n2847), .QN(n36829) );
  DFFRX1 u_decode_u_regfile_reg_r23_q_reg_25_ ( .D(u_decode_u_regfile_N939), 
        .CK(n37880), .RN(n44114), .Q(n2848), .QN(n40903) );
  DFFRX1 u_lsu_mem_data_wr_q_reg_25_ ( .D(u_lsu_N219), .CK(net1847), .RN(
        n44159), .QN(n2849) );
  DFFRX1 u_lsu_mem_addr_q_reg_24_ ( .D(u_lsu_mem_addr_r[24]), .CK(n37876), 
        .RN(n44184), .Q(mmu_lsu_addr_w[24]), .QN(n8322) );
  DFFRX1 u_mmu_lsu_in_addr_q_reg_24_ ( .D(mmu_lsu_addr_w[24]), .CK(n37873), 
        .RN(n44184), .QN(n2850) );
  DFFRX1 u_mmu_itlb_va_addr_q_reg_24_ ( .D(n8429), .CK(clk_i), .RN(n44184), 
        .Q(u_mmu_itlb_va_addr_q[24]) );
  DFFRX1 u_mmu_dtlb_va_addr_q_reg_24_ ( .D(n8428), .CK(clk_i), .RN(n44206), 
        .Q(u_mmu_dtlb_va_addr_q[24]) );
  DFFRX1 u_decode_u_regfile_reg_r25_q_reg_24_ ( .D(u_decode_u_regfile_N1012), 
        .CK(n37837), .RN(n44112), .Q(n2852), .QN(n42476) );
  DFFRX1 u_decode_u_regfile_reg_r26_q_reg_24_ ( .D(u_decode_u_regfile_N1049), 
        .CK(n37836), .RN(n44111), .Q(n2853), .QN(n36822) );
  DFFRX1 u_decode_u_regfile_reg_r27_q_reg_24_ ( .D(u_decode_u_regfile_N1086), 
        .CK(n37835), .RN(n44112), .Q(n2854) );
  DFFRX1 u_decode_u_regfile_reg_r28_q_reg_24_ ( .D(u_decode_u_regfile_N1123), 
        .CK(n37834), .RN(n44111), .Q(n2855) );
  DFFRX1 u_decode_u_regfile_reg_r29_q_reg_24_ ( .D(u_decode_u_regfile_N1160), 
        .CK(n37833), .RN(n44112), .Q(n2856), .QN(n36997) );
  DFFRX1 u_decode_u_regfile_reg_r30_q_reg_24_ ( .D(u_decode_u_regfile_N1197), 
        .CK(n37832), .RN(n44112), .Q(n2857), .QN(n36975) );
  DFFRX1 u_decode_u_regfile_reg_r31_q_reg_24_ ( .D(u_decode_u_regfile_N1234), 
        .CK(n37831), .RN(n44112), .Q(n2858) );
  DFFRX1 u_decode_u_regfile_reg_r1_q_reg_24_ ( .D(u_decode_u_regfile_N124), 
        .CK(n37830), .RN(n44112), .Q(n2859) );
  DFFRX1 u_decode_u_regfile_reg_r2_q_reg_24_ ( .D(u_decode_u_regfile_N161), 
        .CK(n37829), .RN(n44111), .Q(n2860), .QN(n36825) );
  DFFRX1 u_decode_u_regfile_reg_r3_q_reg_24_ ( .D(u_decode_u_regfile_N198), 
        .CK(n37828), .RN(n44112), .Q(n2861), .QN(n40373) );
  DFFRX1 u_decode_u_regfile_reg_r4_q_reg_24_ ( .D(u_decode_u_regfile_N235), 
        .CK(n37827), .RN(n44111), .Q(n2862), .QN(n37001) );
  DFFRX1 u_decode_u_regfile_reg_r5_q_reg_24_ ( .D(u_decode_u_regfile_N272), 
        .CK(n37826), .RN(n44112), .Q(n2863), .QN(n37012) );
  DFFRX1 u_decode_u_regfile_reg_r6_q_reg_24_ ( .D(u_decode_u_regfile_N309), 
        .CK(n37825), .RN(n44112), .Q(n2864), .QN(n36957) );
  DFFRX1 u_decode_u_regfile_reg_r7_q_reg_24_ ( .D(u_decode_u_regfile_N346), 
        .CK(n37824), .RN(n44113), .Q(n2865), .QN(n37321) );
  DFFRX1 u_decode_u_regfile_reg_r8_q_reg_24_ ( .D(u_decode_u_regfile_N383), 
        .CK(n37823), .RN(n44095), .Q(n2866), .QN(n40600) );
  DFFRX1 u_decode_u_regfile_reg_r9_q_reg_24_ ( .D(u_decode_u_regfile_N420), 
        .CK(n37822), .RN(n44112), .Q(n2867) );
  DFFRX1 u_decode_u_regfile_reg_r10_q_reg_24_ ( .D(u_decode_u_regfile_N457), 
        .CK(n37821), .RN(n44095), .Q(n2868), .QN(n36826) );
  DFFRX1 u_decode_u_regfile_reg_r11_q_reg_24_ ( .D(u_decode_u_regfile_N494), 
        .CK(n37820), .RN(n44112), .Q(n2869) );
  DFFRX1 u_decode_u_regfile_reg_r12_q_reg_24_ ( .D(u_decode_u_regfile_N531), 
        .CK(n37819), .RN(n44111), .Q(n2870), .QN(n36985) );
  DFFRX1 u_decode_u_regfile_reg_r13_q_reg_24_ ( .D(u_decode_u_regfile_N568), 
        .CK(n37818), .RN(n44112), .Q(n2871), .QN(n37010) );
  DFFRX1 u_decode_u_regfile_reg_r14_q_reg_24_ ( .D(u_decode_u_regfile_N605), 
        .CK(n37817), .RN(n44112), .Q(n2872), .QN(n36992) );
  DFFRX1 u_decode_u_regfile_reg_r15_q_reg_24_ ( .D(u_decode_u_regfile_N642), 
        .CK(n37816), .RN(n44112), .Q(n2873), .QN(n36983) );
  DFFRX1 u_decode_u_regfile_reg_r16_q_reg_24_ ( .D(u_decode_u_regfile_N679), 
        .CK(n37815), .RN(n44095), .Q(n2874) );
  DFFRX1 u_decode_u_regfile_reg_r17_q_reg_24_ ( .D(u_decode_u_regfile_N716), 
        .CK(n37814), .RN(n44112), .Q(n2875) );
  DFFRX1 u_decode_u_regfile_reg_r18_q_reg_24_ ( .D(u_decode_u_regfile_N753), 
        .CK(n37813), .RN(n44115), .Q(n2876), .QN(n36821) );
  DFFRX1 u_decode_u_regfile_reg_r19_q_reg_24_ ( .D(u_decode_u_regfile_N790), 
        .CK(n37812), .RN(n44112), .Q(n2877), .QN(n40861) );
  DFFRX1 u_decode_u_regfile_reg_r20_q_reg_24_ ( .D(u_decode_u_regfile_N827), 
        .CK(n37811), .RN(n44111), .Q(n2878), .QN(n37013) );
  DFFRX1 u_decode_u_regfile_reg_r21_q_reg_24_ ( .D(u_decode_u_regfile_N864), 
        .CK(n37810), .RN(n44112), .Q(n2879) );
  DFFRX1 u_decode_u_regfile_reg_r22_q_reg_24_ ( .D(u_decode_u_regfile_N901), 
        .CK(n37809), .RN(n44111), .Q(n2880), .QN(n36998) );
  DFFRX1 u_decode_u_regfile_reg_r23_q_reg_24_ ( .D(u_decode_u_regfile_N938), 
        .CK(n37880), .RN(n44112), .Q(n2881), .QN(n36980) );
  DFFRX1 u_lsu_mem_addr_q_reg_17_ ( .D(u_lsu_mem_addr_r[17]), .CK(n37876), 
        .RN(n44183), .Q(mmu_lsu_addr_w[17]), .QN(n8306) );
  DFFRX1 u_mmu_lsu_in_addr_q_reg_17_ ( .D(mmu_lsu_addr_w[17]), .CK(n37873), 
        .RN(n44183), .QN(n2882) );
  DFFRX1 u_mmu_itlb_va_addr_q_reg_17_ ( .D(u_mmu_virt_addr_q[17]), .CK(n37871), 
        .RN(n44184), .Q(n2883) );
  DFFRX1 u_mmu_dtlb_va_addr_q_reg_17_ ( .D(u_mmu_virt_addr_q[17]), .CK(n37872), 
        .RN(n44206), .Q(u_mmu_dtlb_va_addr_q[17]) );
  DFFRX1 u_mmu_itlb_entry_q_reg_17_ ( .D(u_mmu_pte_entry_q[17]), .CK(net1792), 
        .RN(n44171), .Q(u_mmu_itlb_entry_q[17]) );
  DFFRX1 u_mmu_dtlb_entry_q_reg_17_ ( .D(u_mmu_pte_entry_q[17]), .CK(net1782), 
        .RN(n44196), .QN(n2884) );
  DFFRX1 u_muldiv_dividend_q_reg_17_ ( .D(u_muldiv_N249), .CK(net1913), .RN(
        n44158), .Q(u_muldiv_dividend_q[17]) );
  DFFRX1 u_decode_u_regfile_reg_r25_q_reg_17_ ( .D(u_decode_u_regfile_N1005), 
        .CK(n37837), .RN(n44099), .Q(n2885), .QN(n37165) );
  DFFRX1 u_decode_u_regfile_reg_r26_q_reg_17_ ( .D(u_decode_u_regfile_N1042), 
        .CK(n37836), .RN(n44099), .Q(n2886), .QN(n37004) );
  DFFRX1 u_decode_u_regfile_reg_r27_q_reg_17_ ( .D(u_decode_u_regfile_N1079), 
        .CK(n37835), .RN(n44099), .Q(n2887) );
  DFFRX1 u_decode_u_regfile_reg_r28_q_reg_17_ ( .D(u_decode_u_regfile_N1116), 
        .CK(n37834), .RN(n44099), .Q(n2888) );
  DFFRX1 u_decode_u_regfile_reg_r29_q_reg_17_ ( .D(u_decode_u_regfile_N1153), 
        .CK(n37833), .RN(n44100), .Q(n2889), .QN(n37006) );
  DFFRX1 u_decode_u_regfile_reg_r1_q_reg_17_ ( .D(u_decode_u_regfile_N117), 
        .CK(n37830), .RN(n44099), .Q(n2890), .QN(n37169) );
  DFFRX1 u_decode_u_regfile_reg_r30_q_reg_17_ ( .D(u_decode_u_regfile_N1190), 
        .CK(n37832), .RN(n44099), .Q(n2891) );
  DFFRX1 u_decode_u_regfile_reg_r31_q_reg_17_ ( .D(u_decode_u_regfile_N1227), 
        .CK(n37831), .RN(n44100), .Q(n2892) );
  DFFRX1 u_decode_u_regfile_reg_r2_q_reg_17_ ( .D(u_decode_u_regfile_N154), 
        .CK(n37829), .RN(n44099), .Q(n2893), .QN(n36988) );
  DFFRX1 u_decode_u_regfile_reg_r3_q_reg_17_ ( .D(u_decode_u_regfile_N191), 
        .CK(n37828), .RN(n44099), .Q(n2894), .QN(n37156) );
  DFFRX1 u_decode_u_regfile_reg_r4_q_reg_17_ ( .D(u_decode_u_regfile_N228), 
        .CK(n37827), .RN(n44099), .Q(n2895), .QN(n37015) );
  DFFRX1 u_decode_u_regfile_reg_r5_q_reg_17_ ( .D(u_decode_u_regfile_N265), 
        .CK(n37826), .RN(n44100), .Q(n2896), .QN(n36987) );
  DFFRX1 u_decode_u_regfile_reg_r6_q_reg_17_ ( .D(u_decode_u_regfile_N302), 
        .CK(n37825), .RN(n44099), .Q(n2897), .QN(n36960) );
  DFFRX1 u_decode_u_regfile_reg_r7_q_reg_17_ ( .D(u_decode_u_regfile_N339), 
        .CK(n37824), .RN(n44100), .Q(n2898), .QN(n37314) );
  DFFRX1 u_decode_u_regfile_reg_r8_q_reg_17_ ( .D(u_decode_u_regfile_N376), 
        .CK(n37823), .RN(n44098), .Q(n2899), .QN(n37155) );
  DFFRX1 u_decode_u_regfile_reg_r9_q_reg_17_ ( .D(u_decode_u_regfile_N413), 
        .CK(n37822), .RN(n44099), .Q(n2900), .QN(n37152) );
  DFFRX1 u_decode_u_regfile_reg_r10_q_reg_17_ ( .D(u_decode_u_regfile_N450), 
        .CK(n37821), .RN(n44098), .Q(n2901), .QN(n37007) );
  DFFRX1 u_decode_u_regfile_reg_r11_q_reg_17_ ( .D(u_decode_u_regfile_N487), 
        .CK(n37820), .RN(n44100), .Q(n2902), .QN(n37159) );
  DFFRX1 u_decode_u_regfile_reg_r12_q_reg_17_ ( .D(u_decode_u_regfile_N524), 
        .CK(n37819), .RN(n44099), .Q(n2903), .QN(n36991) );
  DFFRX1 u_decode_u_regfile_reg_r13_q_reg_17_ ( .D(u_decode_u_regfile_N561), 
        .CK(n37818), .RN(n44100), .Q(n2904), .QN(n36993) );
  DFFRX1 u_decode_u_regfile_reg_r14_q_reg_17_ ( .D(u_decode_u_regfile_N598), 
        .CK(n37817), .RN(n44099), .Q(n2905), .QN(n36964) );
  DFFRX1 u_decode_u_regfile_reg_r15_q_reg_17_ ( .D(u_decode_u_regfile_N635), 
        .CK(n37816), .RN(n44100), .Q(n2906), .QN(n36954) );
  DFFRX1 u_decode_u_regfile_reg_r16_q_reg_17_ ( .D(u_decode_u_regfile_N672), 
        .CK(n37815), .RN(n44098), .Q(n2907) );
  DFFRX1 u_decode_u_regfile_reg_r17_q_reg_17_ ( .D(u_decode_u_regfile_N709), 
        .CK(n37814), .RN(n44099), .Q(n2908) );
  DFFRX1 u_decode_u_regfile_reg_r18_q_reg_17_ ( .D(u_decode_u_regfile_N746), 
        .CK(n37813), .RN(n44098), .Q(n2909) );
  DFFRX1 u_decode_u_regfile_reg_r19_q_reg_17_ ( .D(u_decode_u_regfile_N783), 
        .CK(n37812), .RN(n44099), .Q(n2910), .QN(n37150) );
  DFFRX1 u_decode_u_regfile_reg_r20_q_reg_17_ ( .D(u_decode_u_regfile_N820), 
        .CK(n37811), .RN(n44099), .Q(n2911) );
  DFFRX1 u_decode_u_regfile_reg_r21_q_reg_17_ ( .D(u_decode_u_regfile_N857), 
        .CK(n37810), .RN(n44100), .Q(n2912) );
  DFFRX1 u_decode_u_regfile_reg_r22_q_reg_17_ ( .D(u_decode_u_regfile_N894), 
        .CK(n37809), .RN(n44099), .Q(n2913) );
  DFFRX1 u_decode_u_regfile_reg_r23_q_reg_17_ ( .D(u_decode_u_regfile_N931), 
        .CK(n37880), .RN(n44100), .Q(n2914), .QN(n36972) );
  DFFRX1 u_lsu_mem_data_wr_q_reg_17_ ( .D(u_lsu_N211), .CK(net1847), .RN(
        n44158), .QN(n2915) );
  DFFRX1 u_fetch_branch_pc_q_reg_31_ ( .D(net2317), .CK(n37866), .RN(n44183), 
        .QN(n2916) );
  DFFRX1 u_decode_u_regfile_reg_r25_q_reg_31_ ( .D(u_decode_u_regfile_N1019), 
        .CK(n37837), .RN(n44188), .Q(n2917), .QN(n40897) );
  DFFRX1 u_decode_u_regfile_reg_r26_q_reg_31_ ( .D(u_decode_u_regfile_N1056), 
        .CK(n37836), .RN(n44203), .Q(n2918) );
  DFFRX1 u_decode_u_regfile_reg_r27_q_reg_31_ ( .D(u_decode_u_regfile_N1093), 
        .CK(n37835), .RN(n44187), .Q(n2919), .QN(n36880) );
  DFFRX1 u_decode_u_regfile_reg_r28_q_reg_31_ ( .D(u_decode_u_regfile_N1130), 
        .CK(n37834), .RN(n44207), .Q(n2920), .QN(n36795) );
  DFFRX1 u_decode_u_regfile_reg_r29_q_reg_31_ ( .D(u_decode_u_regfile_N1167), 
        .CK(n37833), .RN(n44203), .Q(n2921) );
  DFFRX1 u_decode_u_regfile_reg_r30_q_reg_31_ ( .D(u_decode_u_regfile_N1204), 
        .CK(n37832), .RN(n44203), .Q(n2922), .QN(n40884) );
  DFFRX1 u_decode_u_regfile_reg_r31_q_reg_31_ ( .D(u_decode_u_regfile_N1241), 
        .CK(n37831), .RN(n44204), .Q(n2923) );
  DFFRX1 u_decode_u_regfile_reg_r1_q_reg_31_ ( .D(u_decode_u_regfile_N131), 
        .CK(n37830), .RN(n44187), .Q(n2924), .QN(n36832) );
  DFFRX1 u_decode_u_regfile_reg_r2_q_reg_31_ ( .D(u_decode_u_regfile_N168), 
        .CK(n37829), .RN(n44203), .Q(n2925) );
  DFFRX1 u_decode_u_regfile_reg_r3_q_reg_31_ ( .D(u_decode_u_regfile_N205), 
        .CK(n37828), .RN(n44187), .Q(n2926), .QN(n36877) );
  DFFRX1 u_decode_u_regfile_reg_r4_q_reg_31_ ( .D(u_decode_u_regfile_N242), 
        .CK(n37827), .RN(n44203), .Q(n2927), .QN(n36797) );
  DFFRX1 u_decode_u_regfile_reg_r5_q_reg_31_ ( .D(u_decode_u_regfile_N279), 
        .CK(n37826), .RN(n44204), .Q(n2928), .QN(n40908) );
  DFFRX1 u_decode_u_regfile_reg_r6_q_reg_31_ ( .D(u_decode_u_regfile_N316), 
        .CK(n37825), .RN(n44203), .Q(n2929), .QN(n40906) );
  DFFRX1 u_decode_u_regfile_reg_r7_q_reg_31_ ( .D(u_decode_u_regfile_N353), 
        .CK(n37824), .RN(n44204), .QN(n36796) );
  DFFRX1 u_decode_u_regfile_reg_r8_q_reg_31_ ( .D(u_decode_u_regfile_N390), 
        .CK(n37823), .RN(n44187), .Q(n2931), .QN(n36818) );
  DFFRX1 u_decode_u_regfile_reg_r9_q_reg_31_ ( .D(u_decode_u_regfile_N427), 
        .CK(n37822), .RN(n44188), .Q(n2932), .QN(n40885) );
  DFFRX1 u_decode_u_regfile_reg_r10_q_reg_31_ ( .D(u_decode_u_regfile_N464), 
        .CK(n37821), .RN(n44203), .Q(n2933) );
  DFFRX1 u_decode_u_regfile_reg_r11_q_reg_31_ ( .D(u_decode_u_regfile_N501), 
        .CK(n37820), .RN(n44187), .Q(n2934), .QN(n37067) );
  DFFRX1 u_decode_u_regfile_reg_r12_q_reg_31_ ( .D(u_decode_u_regfile_N538), 
        .CK(n37819), .RN(n44204), .Q(n2935) );
  DFFRX1 u_decode_u_regfile_reg_r13_q_reg_31_ ( .D(u_decode_u_regfile_N575), 
        .CK(n37818), .RN(n44203), .Q(n2936), .QN(n40877) );
  DFFRX1 u_decode_u_regfile_reg_r14_q_reg_31_ ( .D(u_decode_u_regfile_N612), 
        .CK(n37817), .RN(n44204), .Q(n2937), .QN(n36843) );
  DFFRX1 u_decode_u_regfile_reg_r15_q_reg_31_ ( .D(u_decode_u_regfile_N649), 
        .CK(n37816), .RN(n44204), .Q(n2938), .QN(n40875) );
  DFFRX1 u_decode_u_regfile_reg_r16_q_reg_31_ ( .D(u_decode_u_regfile_N686), 
        .CK(n37815), .RN(n44187), .Q(n2939), .QN(n37074) );
  DFFRX1 u_decode_u_regfile_reg_r17_q_reg_31_ ( .D(u_decode_u_regfile_N723), 
        .CK(n37814), .RN(n44187), .Q(n2940) );
  DFFRX1 u_decode_u_regfile_reg_r18_q_reg_31_ ( .D(u_decode_u_regfile_N760), 
        .CK(n37813), .RN(n44204), .Q(n2941) );
  DFFRX1 u_decode_u_regfile_reg_r19_q_reg_31_ ( .D(u_decode_u_regfile_N797), 
        .CK(n37812), .RN(n44187), .Q(n2942) );
  DFFRX1 u_decode_u_regfile_reg_r20_q_reg_31_ ( .D(u_decode_u_regfile_N834), 
        .CK(n37811), .RN(n44203), .Q(n2943) );
  DFFRX1 u_decode_u_regfile_reg_r21_q_reg_31_ ( .D(u_decode_u_regfile_N871), 
        .CK(n37810), .RN(n44203), .Q(n2944) );
  DFFRX1 u_decode_u_regfile_reg_r22_q_reg_31_ ( .D(u_decode_u_regfile_N908), 
        .CK(n37809), .RN(n44204), .Q(n2945) );
  DFFRX1 u_lsu_mem_data_wr_q_reg_5_ ( .D(u_lsu_N199), .CK(n37874), .RN(n44200), 
        .QN(n2946) );
  DFFRX1 u_lsu_mem_data_wr_q_reg_13_ ( .D(u_lsu_N207), .CK(net1847), .RN(
        n44158), .QN(n2947) );
  DFFRX1 u_lsu_mem_data_wr_q_reg_21_ ( .D(u_lsu_N215), .CK(net1847), .RN(
        n44158), .QN(n2948) );
  DFFRX1 u_lsu_mem_data_wr_q_reg_0_ ( .D(u_lsu_N194), .CK(n37874), .RN(n44200), 
        .QN(n2949) );
  DFFRX1 u_lsu_mem_data_wr_q_reg_8_ ( .D(u_lsu_N202), .CK(n37874), .RN(n44158), 
        .QN(n2950) );
  DFFRX1 u_lsu_mem_data_wr_q_reg_16_ ( .D(u_lsu_N210), .CK(net1847), .RN(
        n44158), .QN(n2951) );
  DFFRX1 u_lsu_mem_data_wr_q_reg_24_ ( .D(u_lsu_N218), .CK(net1847), .RN(
        n44158), .QN(n2952) );
  DFFRX1 u_lsu_mem_data_wr_q_reg_28_ ( .D(u_lsu_N222), .CK(net1847), .RN(
        n44158), .QN(n2953) );
  DFFRX1 u_decode_u_regfile_reg_r25_q_reg_30_ ( .D(u_decode_u_regfile_N1018), 
        .CK(n37837), .RN(n44181), .Q(n2954), .QN(n42510) );
  DFFRX1 u_decode_u_regfile_reg_r26_q_reg_30_ ( .D(u_decode_u_regfile_N1055), 
        .CK(n37836), .RN(n44180), .Q(n2955), .QN(n36792) );
  DFFRX1 u_decode_u_regfile_reg_r27_q_reg_30_ ( .D(u_decode_u_regfile_N1092), 
        .CK(n37835), .RN(n44181), .Q(n2956) );
  DFFRX1 u_decode_u_regfile_reg_r28_q_reg_30_ ( .D(u_decode_u_regfile_N1129), 
        .CK(n37834), .RN(n44180), .Q(n2957), .QN(n40850) );
  DFFRX1 u_decode_u_regfile_reg_r29_q_reg_30_ ( .D(u_decode_u_regfile_N1166), 
        .CK(n37833), .RN(n44181), .Q(n2958) );
  DFFRX1 u_decode_u_regfile_reg_r30_q_reg_30_ ( .D(u_decode_u_regfile_N1203), 
        .CK(n37832), .RN(n44181), .Q(n2959), .QN(n36794) );
  DFFRX1 u_decode_u_regfile_reg_r31_q_reg_30_ ( .D(u_decode_u_regfile_N1240), 
        .CK(n37831), .RN(n44181), .Q(n2960), .QN(n40852) );
  DFFRX1 u_decode_u_regfile_reg_r1_q_reg_30_ ( .D(u_decode_u_regfile_N130), 
        .CK(n37830), .RN(n44181), .Q(n2961) );
  DFFRX1 u_decode_u_regfile_reg_r2_q_reg_30_ ( .D(u_decode_u_regfile_N167), 
        .CK(n37829), .RN(n44180), .Q(n2962) );
  DFFRX1 u_decode_u_regfile_reg_r3_q_reg_30_ ( .D(u_decode_u_regfile_N204), 
        .CK(n37828), .RN(n44181), .Q(n2963), .QN(n42505) );
  DFFRX1 u_decode_u_regfile_reg_r4_q_reg_30_ ( .D(u_decode_u_regfile_N241), 
        .CK(n37827), .RN(n44180), .Q(n2964), .QN(n36827) );
  DFFRX1 u_decode_u_regfile_reg_r5_q_reg_30_ ( .D(u_decode_u_regfile_N278), 
        .CK(n37826), .RN(n44181), .Q(n2965), .QN(n40895) );
  DFFRX1 u_decode_u_regfile_reg_r6_q_reg_30_ ( .D(u_decode_u_regfile_N315), 
        .CK(n37825), .RN(n44181), .Q(n2966), .QN(n40887) );
  DFFRX1 u_decode_u_regfile_reg_r7_q_reg_30_ ( .D(u_decode_u_regfile_N352), 
        .CK(n37824), .RN(n44182), .QN(n36823) );
  DFFRX1 u_decode_u_regfile_reg_r8_q_reg_30_ ( .D(u_decode_u_regfile_N389), 
        .CK(n37823), .RN(n44180), .Q(n2968) );
  DFFRX1 u_decode_u_regfile_reg_r9_q_reg_30_ ( .D(u_decode_u_regfile_N426), 
        .CK(n37822), .RN(n44181), .Q(n2969) );
  DFFRX1 u_decode_u_regfile_reg_r10_q_reg_30_ ( .D(u_decode_u_regfile_N463), 
        .CK(n37821), .RN(n44180), .Q(n2970) );
  DFFRX1 u_decode_u_regfile_reg_r11_q_reg_30_ ( .D(u_decode_u_regfile_N500), 
        .CK(n37820), .RN(n44181), .Q(n2971) );
  DFFRX1 u_decode_u_regfile_reg_r12_q_reg_30_ ( .D(u_decode_u_regfile_N537), 
        .CK(n37819), .RN(n44180), .Q(n2972), .QN(n36834) );
  DFFRX1 u_decode_u_regfile_reg_r13_q_reg_30_ ( .D(u_decode_u_regfile_N574), 
        .CK(n37818), .RN(n44181), .Q(n2973) );
  DFFRX1 u_decode_u_regfile_reg_r14_q_reg_30_ ( .D(u_decode_u_regfile_N611), 
        .CK(n37817), .RN(n44181), .Q(n2974), .QN(n36793) );
  DFFRX1 u_decode_u_regfile_reg_r15_q_reg_30_ ( .D(u_decode_u_regfile_N648), 
        .CK(n37816), .RN(n44181), .Q(n2975) );
  DFFRX1 u_decode_u_regfile_reg_r16_q_reg_30_ ( .D(u_decode_u_regfile_N685), 
        .CK(n37815), .RN(n44180), .Q(n2976), .QN(n42511) );
  DFFRX1 u_decode_u_regfile_reg_r17_q_reg_30_ ( .D(u_decode_u_regfile_N722), 
        .CK(n37814), .RN(n44181), .Q(n2977) );
  DFFRX1 u_decode_u_regfile_reg_r19_q_reg_30_ ( .D(u_decode_u_regfile_N796), 
        .CK(n37812), .RN(n44181), .Q(n2979), .QN(n42507) );
  DFFRX1 u_decode_u_regfile_reg_r20_q_reg_30_ ( .D(u_decode_u_regfile_N833), 
        .CK(n37811), .RN(n44180), .Q(n2980) );
  DFFRX1 u_decode_u_regfile_reg_r22_q_reg_30_ ( .D(u_decode_u_regfile_N907), 
        .CK(n37809), .RN(n44180), .Q(n2982), .QN(n36824) );
  DFFRX1 u_decode_u_regfile_reg_r25_q_reg_29_ ( .D(u_decode_u_regfile_N1017), 
        .CK(n37837), .RN(n44195), .Q(n2983), .QN(n36940) );
  DFFRX1 u_decode_u_regfile_reg_r26_q_reg_29_ ( .D(u_decode_u_regfile_N1054), 
        .CK(n37836), .RN(n44194), .Q(n2984), .QN(n36848) );
  DFFRX1 u_decode_u_regfile_reg_r27_q_reg_29_ ( .D(u_decode_u_regfile_N1091), 
        .CK(n37835), .RN(n44195), .Q(n2985), .QN(n36935) );
  DFFRX1 u_decode_u_regfile_reg_r28_q_reg_29_ ( .D(u_decode_u_regfile_N1128), 
        .CK(n37834), .RN(n44194), .Q(n2986) );
  DFFRX1 u_decode_u_regfile_reg_r29_q_reg_29_ ( .D(u_decode_u_regfile_N1165), 
        .CK(n37833), .RN(n44195), .Q(n2987) );
  DFFRX1 u_decode_u_regfile_reg_r30_q_reg_29_ ( .D(u_decode_u_regfile_N1202), 
        .CK(n37832), .RN(n44194), .Q(n2988) );
  DFFRX1 u_decode_u_regfile_reg_r31_q_reg_29_ ( .D(u_decode_u_regfile_N1239), 
        .CK(n37831), .RN(n44195), .Q(n2989) );
  DFFRX1 u_decode_u_regfile_reg_r1_q_reg_29_ ( .D(u_decode_u_regfile_N129), 
        .CK(n37830), .RN(n44195), .Q(n2990) );
  DFFRX1 u_decode_u_regfile_reg_r2_q_reg_29_ ( .D(u_decode_u_regfile_N166), 
        .CK(n37829), .RN(n44194), .Q(n2991), .QN(n40865) );
  DFFRX1 u_decode_u_regfile_reg_r3_q_reg_29_ ( .D(u_decode_u_regfile_N203), 
        .CK(n37828), .RN(n44195), .Q(n2992), .QN(n37037) );
  DFFRX1 u_decode_u_regfile_reg_r4_q_reg_29_ ( .D(u_decode_u_regfile_N240), 
        .CK(n37827), .RN(n44194), .Q(n2993) );
  DFFRX1 u_decode_u_regfile_reg_r5_q_reg_29_ ( .D(u_decode_u_regfile_N277), 
        .CK(n37826), .RN(n44195), .Q(n2994) );
  DFFRX1 u_decode_u_regfile_reg_r6_q_reg_29_ ( .D(u_decode_u_regfile_N314), 
        .CK(n37825), .RN(n44194), .Q(n2995) );
  DFFRX1 u_decode_u_regfile_reg_r7_q_reg_29_ ( .D(u_decode_u_regfile_N351), 
        .CK(n37824), .RN(n44195), .Q(n2996), .QN(n37324) );
  DFFRX1 u_decode_u_regfile_reg_r8_q_reg_29_ ( .D(u_decode_u_regfile_N388), 
        .CK(n37823), .RN(n44194), .Q(n2997), .QN(n37034) );
  DFFRX1 u_decode_u_regfile_reg_r9_q_reg_29_ ( .D(u_decode_u_regfile_N425), 
        .CK(n37822), .RN(n44195), .Q(n2998), .QN(n37045) );
  DFFRX1 u_decode_u_regfile_reg_r10_q_reg_29_ ( .D(u_decode_u_regfile_N462), 
        .CK(n37821), .RN(n44194), .Q(n2999), .QN(n40869) );
  DFFRX1 u_decode_u_regfile_reg_r11_q_reg_29_ ( .D(u_decode_u_regfile_N499), 
        .CK(n37820), .RN(n44195), .Q(n3000), .QN(n37094) );
  DFFRX1 u_decode_u_regfile_reg_r12_q_reg_29_ ( .D(u_decode_u_regfile_N536), 
        .CK(n37819), .RN(n44194), .Q(n3001) );
  DFFRX1 u_decode_u_regfile_reg_r13_q_reg_29_ ( .D(u_decode_u_regfile_N573), 
        .CK(n37818), .RN(n44195), .Q(n3002) );
  DFFRX1 u_decode_u_regfile_reg_r14_q_reg_29_ ( .D(u_decode_u_regfile_N610), 
        .CK(n37817), .RN(n44194), .Q(n3003) );
  DFFRX1 u_decode_u_regfile_reg_r15_q_reg_29_ ( .D(u_decode_u_regfile_N647), 
        .CK(n37816), .RN(n44195), .Q(n3004) );
  DFFRX1 u_decode_u_regfile_reg_r16_q_reg_29_ ( .D(u_decode_u_regfile_N684), 
        .CK(n37815), .RN(n44194), .Q(n3005) );
  DFFRX1 u_decode_u_regfile_reg_r17_q_reg_29_ ( .D(u_decode_u_regfile_N721), 
        .CK(n37814), .RN(n44195), .Q(n3006), .QN(n37048) );
  DFFRX1 u_decode_u_regfile_reg_r18_q_reg_29_ ( .D(u_decode_u_regfile_N758), 
        .CK(n37813), .RN(n44194), .Q(n3007), .QN(n36841) );
  DFFRX1 u_decode_u_regfile_reg_r19_q_reg_29_ ( .D(u_decode_u_regfile_N795), 
        .CK(n37812), .RN(n44195), .Q(n3008), .QN(n37029) );
  DFFRX1 u_decode_u_regfile_reg_r22_q_reg_29_ ( .D(u_decode_u_regfile_N906), 
        .CK(n37809), .RN(n44194), .Q(n3011) );
  DFFRX1 u_lsu_mem_data_wr_q_reg_29_ ( .D(u_lsu_N223), .CK(n37868), .RN(n44158), .QN(n3012) );
  DFFRX1 u_muldiv_divisor_q_reg_58_ ( .D(u_muldiv_N323), .CK(net1898), .RN(
        n44158), .Q(u_muldiv_divisor_q[58]) );
  DFFRX1 u_muldiv_divisor_q_reg_57_ ( .D(u_muldiv_N322), .CK(net1898), .RN(
        n44158), .Q(u_muldiv_divisor_q[57]) );
  DFFRX1 u_muldiv_divisor_q_reg_56_ ( .D(u_muldiv_N321), .CK(net1898), .RN(
        n44158), .Q(u_muldiv_divisor_q[56]) );
  DFFRX1 u_muldiv_divisor_q_reg_55_ ( .D(u_muldiv_N320), .CK(net1898), .RN(
        n44158), .Q(u_muldiv_divisor_q[55]) );
  DFFRX1 u_muldiv_divisor_q_reg_54_ ( .D(u_muldiv_N319), .CK(net1898), .RN(
        n44157), .Q(u_muldiv_divisor_q[54]) );
  DFFRX1 u_muldiv_divisor_q_reg_53_ ( .D(u_muldiv_N318), .CK(net1898), .RN(
        n44157), .Q(u_muldiv_divisor_q[53]) );
  DFFRX1 u_muldiv_divisor_q_reg_52_ ( .D(u_muldiv_N317), .CK(net1898), .RN(
        n44157), .Q(u_muldiv_divisor_q[52]) );
  DFFRX1 u_muldiv_divisor_q_reg_51_ ( .D(u_muldiv_N316), .CK(net1898), .RN(
        n44157), .Q(u_muldiv_divisor_q[51]) );
  DFFRX1 u_muldiv_divisor_q_reg_50_ ( .D(u_muldiv_N315), .CK(net1898), .RN(
        n44157), .Q(u_muldiv_divisor_q[50]) );
  DFFRX1 u_muldiv_divisor_q_reg_49_ ( .D(u_muldiv_N314), .CK(net1898), .RN(
        n44157), .Q(u_muldiv_divisor_q[49]) );
  DFFRX1 u_muldiv_divisor_q_reg_48_ ( .D(u_muldiv_N313), .CK(net1898), .RN(
        n44157), .Q(u_muldiv_divisor_q[48]) );
  DFFRX1 u_muldiv_divisor_q_reg_47_ ( .D(u_muldiv_N312), .CK(net1893), .RN(
        n44157), .Q(u_muldiv_divisor_q[47]) );
  DFFRX1 u_decode_u_regfile_reg_r25_q_reg_14_ ( .D(u_decode_u_regfile_N1002), 
        .CK(n37879), .RN(n44096), .Q(n3013), .QN(n37177) );
  DFFRX1 u_decode_u_regfile_reg_r26_q_reg_14_ ( .D(u_decode_u_regfile_N1039), 
        .CK(n37864), .RN(n44095), .Q(n3014) );
  DFFRX1 u_decode_u_regfile_reg_r27_q_reg_14_ ( .D(u_decode_u_regfile_N1076), 
        .CK(n37863), .RN(n44096), .Q(n3015) );
  DFFRX1 u_decode_u_regfile_reg_r28_q_reg_14_ ( .D(u_decode_u_regfile_N1113), 
        .CK(n37862), .RN(n44095), .Q(n3016), .QN(n36869) );
  DFFRX1 u_decode_u_regfile_reg_r1_q_reg_14_ ( .D(u_decode_u_regfile_N114), 
        .CK(n37865), .RN(n44096), .Q(n3017), .QN(n37181) );
  DFFRX1 u_decode_u_regfile_reg_r29_q_reg_14_ ( .D(u_decode_u_regfile_N1150), 
        .CK(n37861), .RN(n44096), .Q(n3018) );
  DFFRX1 u_decode_u_regfile_reg_r30_q_reg_14_ ( .D(u_decode_u_regfile_N1187), 
        .CK(n37860), .RN(n44095), .Q(n3019), .QN(n36854) );
  DFFRX1 u_decode_u_regfile_reg_r31_q_reg_14_ ( .D(u_decode_u_regfile_N1224), 
        .CK(n37859), .RN(n44096), .Q(n3020), .QN(n36858) );
  DFFRX1 u_decode_u_regfile_reg_r2_q_reg_14_ ( .D(u_decode_u_regfile_N151), 
        .CK(n37858), .RN(n44095), .Q(n3021), .QN(n40642) );
  DFFRX1 u_decode_u_regfile_reg_r3_q_reg_14_ ( .D(u_decode_u_regfile_N188), 
        .CK(n37857), .RN(n44096), .Q(n3022), .QN(n37144) );
  DFFRX1 u_decode_u_regfile_reg_r4_q_reg_14_ ( .D(u_decode_u_regfile_N225), 
        .CK(n37856), .RN(n44095), .Q(n3023) );
  DFFRX1 u_decode_u_regfile_reg_r5_q_reg_14_ ( .D(u_decode_u_regfile_N262), 
        .CK(n37840), .RN(n44096), .Q(n3024) );
  DFFRX1 u_decode_u_regfile_reg_r6_q_reg_14_ ( .D(u_decode_u_regfile_N299), 
        .CK(n37855), .RN(n44095), .Q(n3025) );
  DFFRX1 u_decode_u_regfile_reg_r7_q_reg_14_ ( .D(u_decode_u_regfile_N336), 
        .CK(n37854), .RN(n44096), .QN(n36864) );
  DFFRX1 u_decode_u_regfile_reg_r8_q_reg_14_ ( .D(u_decode_u_regfile_N373), 
        .CK(n37839), .RN(n44103), .Q(n3027), .QN(n37178) );
  DFFRX1 u_decode_u_regfile_reg_r9_q_reg_14_ ( .D(u_decode_u_regfile_N410), 
        .CK(n37853), .RN(n44096), .Q(n3028), .QN(n37176) );
  DFFRX1 u_decode_u_regfile_reg_r10_q_reg_14_ ( .D(u_decode_u_regfile_N447), 
        .CK(n37852), .RN(n44099), .Q(n3029) );
  DFFRX1 u_decode_u_regfile_reg_r11_q_reg_14_ ( .D(u_decode_u_regfile_N484), 
        .CK(n37851), .RN(n44096), .Q(n3030), .QN(n37175) );
  DFFRX1 u_decode_u_regfile_reg_r12_q_reg_14_ ( .D(u_decode_u_regfile_N521), 
        .CK(n37850), .RN(n44095), .Q(n3031) );
  DFFRX1 u_decode_u_regfile_reg_r13_q_reg_14_ ( .D(u_decode_u_regfile_N558), 
        .CK(n37849), .RN(n44096), .Q(n3032) );
  DFFRX1 u_decode_u_regfile_reg_r14_q_reg_14_ ( .D(u_decode_u_regfile_N595), 
        .CK(n37848), .RN(n44095), .Q(n3033) );
  DFFRX1 u_decode_u_regfile_reg_r15_q_reg_14_ ( .D(u_decode_u_regfile_N632), 
        .CK(n37847), .RN(n44096), .Q(n3034) );
  DFFRX1 u_decode_u_regfile_reg_r16_q_reg_14_ ( .D(u_decode_u_regfile_N669), 
        .CK(n37846), .RN(n44140), .Q(n3035), .QN(n37174) );
  DFFRX1 u_decode_u_regfile_reg_r17_q_reg_14_ ( .D(u_decode_u_regfile_N706), 
        .CK(n37845), .RN(n44096), .Q(n3036), .QN(n37148) );
  DFFRX1 u_decode_u_regfile_reg_r18_q_reg_14_ ( .D(u_decode_u_regfile_N743), 
        .CK(n37844), .RN(n44095), .Q(n3037), .QN(n36863) );
  DFFRX1 u_decode_u_regfile_reg_r19_q_reg_14_ ( .D(u_decode_u_regfile_N780), 
        .CK(n37843), .RN(n44096), .Q(n3038), .QN(n37173) );
  DFFRX1 u_decode_u_regfile_reg_r20_q_reg_14_ ( .D(u_decode_u_regfile_N817), 
        .CK(n37842), .RN(n44095), .Q(n3039), .QN(n36857) );
  DFFRX1 u_decode_u_regfile_reg_r21_q_reg_14_ ( .D(u_decode_u_regfile_N854), 
        .CK(n37838), .RN(n44096), .Q(n3040), .QN(n36859) );
  DFFRX1 u_decode_u_regfile_reg_r22_q_reg_14_ ( .D(u_decode_u_regfile_N891), 
        .CK(n37841), .RN(n44095), .Q(n3041), .QN(n36847) );
  DFFRX1 u_lsu_mem_data_wr_q_reg_14_ ( .D(u_lsu_N208), .CK(net1847), .RN(
        n44157), .QN(n3042) );
  DFFRX1 u_lsu_mem_data_wr_q_reg_30_ ( .D(u_lsu_N224), .CK(n37868), .RN(n44157), .QN(n3043) );
  DFFRX1 u_mmu_itlb_va_addr_q_reg_30_ ( .D(n8427), .CK(clk_i), .RN(n44182), 
        .Q(u_mmu_itlb_va_addr_q[30]) );
  DFFRX1 u_mmu_dtlb_va_addr_q_reg_30_ ( .D(n8426), .CK(clk_i), .RN(n44206), 
        .Q(u_mmu_dtlb_va_addr_q[30]) );
  DFFRX1 u_mmu_itlb_va_addr_q_reg_31_ ( .D(n8425), .CK(clk_i), .RN(n44183), 
        .Q(u_mmu_itlb_va_addr_q[31]) );
  DFFRX1 u_mmu_dtlb_va_addr_q_reg_31_ ( .D(n8424), .CK(clk_i), .RN(n44206), 
        .Q(u_mmu_dtlb_va_addr_q[31]) );
  DFFRX1 u_mmu_dtlb_va_addr_q_reg_29_ ( .D(n8423), .CK(clk_i), .RN(n44207), 
        .Q(u_mmu_dtlb_va_addr_q[29]) );
  DFFRX1 u_mmu_pte_addr_q_reg_12_ ( .D(U1_U6_Z_12), .CK(n37884), .RN(n44210), 
        .QN(n3044) );
  DFFRX1 u_mmu_pte_addr_q_reg_13_ ( .D(U1_U6_Z_13), .CK(n37884), .RN(n44210), 
        .QN(n3045) );
  DFFRX1 u_mmu_pte_addr_q_reg_14_ ( .D(U1_U6_Z_14), .CK(n37884), .RN(n44211), 
        .QN(n3046) );
  DFFRX1 u_mmu_pte_addr_q_reg_15_ ( .D(U1_U6_Z_15), .CK(n37884), .RN(n44211), 
        .QN(n3047) );
  DFFRX1 u_mmu_pte_addr_q_reg_16_ ( .D(U1_U6_Z_16), .CK(n37808), .RN(n44211), 
        .QN(n3048) );
  DFFRX1 u_mmu_pte_addr_q_reg_17_ ( .D(U1_U6_Z_17), .CK(n37808), .RN(n44196), 
        .QN(n3049) );
  DFFRX1 u_mmu_pte_addr_q_reg_18_ ( .D(U1_U6_Z_18), .CK(n37808), .RN(n44196), 
        .QN(n3050) );
  DFFRX1 u_mmu_pte_addr_q_reg_19_ ( .D(U1_U6_Z_19), .CK(n37808), .RN(n44196), 
        .QN(n3051) );
  DFFRX1 u_mmu_pte_addr_q_reg_20_ ( .D(U1_U6_Z_20), .CK(n37808), .RN(n44197), 
        .QN(n3052) );
  DFFRX1 u_mmu_pte_addr_q_reg_21_ ( .D(U1_U6_Z_21), .CK(n37808), .RN(n44197), 
        .QN(n3053) );
  DFFRX1 u_mmu_pte_addr_q_reg_22_ ( .D(U1_U6_Z_22), .CK(n37808), .RN(n44197), 
        .QN(n3054) );
  DFFRX1 u_mmu_pte_addr_q_reg_23_ ( .D(U1_U6_Z_23), .CK(n37808), .RN(n44197), 
        .QN(n3055) );
  DFFRX1 u_mmu_pte_addr_q_reg_24_ ( .D(U1_U6_Z_24), .CK(n37808), .RN(n44197), 
        .QN(n3056) );
  DFFRX1 u_mmu_pte_addr_q_reg_25_ ( .D(U1_U6_Z_25), .CK(n37808), .RN(n44197), 
        .QN(n3057) );
  DFFRX1 u_mmu_pte_addr_q_reg_26_ ( .D(U1_U6_Z_26), .CK(n37808), .RN(n44198), 
        .QN(n3058) );
  DFFRX1 u_mmu_pte_addr_q_reg_27_ ( .D(U1_U6_Z_27), .CK(n37808), .RN(n44198), 
        .QN(n3059) );
  DFFRX1 u_mmu_pte_addr_q_reg_28_ ( .D(U1_U6_Z_28), .CK(n37808), .RN(n44198), 
        .QN(n3060) );
  DFFRX1 u_mmu_pte_addr_q_reg_29_ ( .D(U1_U6_Z_29), .CK(n37808), .RN(n44198), 
        .QN(n3061) );
  DFFRX1 u_mmu_pte_addr_q_reg_30_ ( .D(U1_U6_Z_30), .CK(n37808), .RN(n44198), 
        .QN(n3062) );
  DFFRX1 u_mmu_pte_addr_q_reg_31_ ( .D(U1_U6_Z_31), .CK(n37808), .RN(n44198), 
        .QN(n3063) );
  DFFRX1 u_exec_result_q_reg_14_ ( .D(u_exec_alu_p_w[14]), .CK(clk_i), .RN(
        n44140), .Q(writeback_exec_value_w[14]), .QN(n37678) );
  DFFRX1 u_exec_result_q_reg_29_ ( .D(u_exec_alu_p_w[29]), .CK(clk_i), .RN(
        n44194), .Q(writeback_exec_value_w[29]), .QN(n37686) );
  DFFRX1 u_exec_result_q_reg_15_ ( .D(u_exec_alu_p_w[15]), .CK(clk_i), .RN(
        n44123), .Q(writeback_exec_value_w[15]), .QN(n37671) );
  DFFRX1 u_exec_result_q_reg_11_ ( .D(u_exec_alu_p_w[11]), .CK(clk_i), .RN(
        n44136), .Q(writeback_exec_value_w[11]), .QN(n37676) );
  DFFRX1 u_exec_result_q_reg_19_ ( .D(u_exec_alu_p_w[19]), .CK(clk_i), .RN(
        n44102), .Q(writeback_exec_value_w[19]), .QN(n37593) );
  DFFRX1 u_exec_result_q_reg_6_ ( .D(u_exec_alu_p_w[6]), .CK(clk_i), .RN(
        n44141), .Q(writeback_exec_value_w[6]), .QN(n37667) );
  DFFRX1 u_exec_result_q_reg_2_ ( .D(u_exec_alu_p_w[2]), .CK(clk_i), .RN(
        n44205), .Q(writeback_exec_value_w[2]), .QN(n37687) );
  DFFRX1 u_exec_result_q_reg_10_ ( .D(u_exec_alu_p_w[10]), .CK(clk_i), .RN(
        n44134), .Q(writeback_exec_value_w[10]), .QN(n37675) );
  DFFRX1 u_exec_result_q_reg_20_ ( .D(u_exec_alu_p_w[20]), .CK(clk_i), .RN(
        n44088), .Q(writeback_exec_value_w[20]), .QN(n37594) );
  DFFRX1 u_exec_result_q_reg_3_ ( .D(u_exec_alu_p_w[3]), .CK(clk_i), .RN(
        n44128), .Q(writeback_exec_value_w[3]), .QN(n37664) );
  DFFRX1 u_exec_result_q_reg_9_ ( .D(u_exec_alu_p_w[9]), .CK(clk_i), .RN(
        n44132), .Q(writeback_exec_value_w[9]), .QN(n37674) );
  DFFRX1 u_exec_result_q_reg_23_ ( .D(u_exec_alu_p_w[23]), .CK(clk_i), .RN(
        n44093), .Q(writeback_exec_value_w[23]), .QN(n37684) );
  DFFRX1 u_exec_result_q_reg_22_ ( .D(u_exec_alu_p_w[22]), .CK(clk_i), .RN(
        n44091), .Q(writeback_exec_value_w[22]), .QN(n37683) );
  DFFRX1 u_exec_result_q_reg_16_ ( .D(u_exec_alu_p_w[16]), .CK(clk_i), .RN(
        n44096), .Q(writeback_exec_value_w[16]), .QN(n37679) );
  DFFRX1 u_exec_result_q_reg_21_ ( .D(u_exec_alu_p_w[21]), .CK(clk_i), .RN(
        n44089), .Q(writeback_exec_value_w[21]), .QN(n37682) );
  DFFRX1 u_exec_result_q_reg_7_ ( .D(u_exec_alu_p_w[7]), .CK(clk_i), .RN(
        n44127), .Q(writeback_exec_value_w[7]), .QN(n37673) );
  DFFRX1 u_exec_result_q_reg_18_ ( .D(u_exec_alu_p_w[18]), .CK(clk_i), .RN(
        n44100), .Q(writeback_exec_value_w[18]), .QN(n37681) );
  DFFRX1 u_exec_result_q_reg_12_ ( .D(u_exec_alu_p_w[12]), .CK(clk_i), .RN(
        n44138), .Q(writeback_exec_value_w[12]), .QN(n37677) );
  DFFRX1 u_exec_result_q_reg_8_ ( .D(u_exec_alu_p_w[8]), .CK(clk_i), .RN(
        n44126), .Q(writeback_exec_value_w[8]), .QN(n37672) );
  DFFRX1 u_exec_result_q_reg_4_ ( .D(u_exec_alu_p_w[4]), .CK(clk_i), .RN(
        n44187), .Q(writeback_exec_value_w[4]), .QN(n37669) );
  DFFRX1 u_exec_result_q_reg_1_ ( .D(u_exec_alu_p_w[1]), .CK(clk_i), .RN(
        n44119), .Q(writeback_exec_value_w[1]), .QN(n37666) );
  DFFRX1 u_exec_result_q_reg_13_ ( .D(u_exec_alu_p_w[13]), .CK(clk_i), .RN(
        n44121), .Q(writeback_exec_value_w[13]), .QN(n37670) );
  DFFRX1 u_exec_result_q_reg_25_ ( .D(u_exec_alu_p_w[25]), .CK(clk_i), .RN(
        n44113), .Q(writeback_exec_value_w[25]), .QN(n37596) );
  DFFRX1 u_exec_result_q_reg_24_ ( .D(u_exec_alu_p_w[24]), .CK(clk_i), .RN(
        n44095), .Q(writeback_exec_value_w[24]), .QN(n37595) );
  DFFRX1 u_exec_result_q_reg_17_ ( .D(u_exec_alu_p_w[17]), .CK(clk_i), .RN(
        n44098), .Q(writeback_exec_value_w[17]), .QN(n37680) );
  DFFRX1 u_exec_result_q_reg_5_ ( .D(u_exec_alu_p_w[5]), .CK(clk_i), .RN(
        n44143), .Q(writeback_exec_value_w[5]), .QN(n37668) );
  DFFRX1 u_exec_result_q_reg_0_ ( .D(u_exec_alu_p_w[0]), .CK(clk_i), .RN(
        n44205), .Q(writeback_exec_value_w[0]), .QN(n37665) );
  DFFRX1 u_exec_result_q_reg_28_ ( .D(u_exec_alu_p_w[28]), .CK(clk_i), .RN(
        n44191), .Q(writeback_exec_value_w[28]), .QN(n37685) );
  DFFRX1 u_muldiv_wb_result_q_reg_8_ ( .D(u_muldiv_N529), .CK(clk_i), .RN(
        n44157), .Q(writeback_muldiv_value_w[8]), .QN(n37606) );
  DFFRX1 u_muldiv_wb_result_q_reg_7_ ( .D(u_muldiv_N528), .CK(clk_i), .RN(
        n44157), .Q(writeback_muldiv_value_w[7]), .QN(n37605) );
  DFFRX1 u_muldiv_wb_result_q_reg_9_ ( .D(u_muldiv_N530), .CK(clk_i), .RN(
        n44157), .Q(writeback_muldiv_value_w[9]), .QN(n37607) );
  DFFRX1 u_muldiv_wb_result_q_reg_10_ ( .D(u_muldiv_N531), .CK(clk_i), .RN(
        n44157), .Q(writeback_muldiv_value_w[10]), .QN(n37608) );
  DFFRX1 u_muldiv_wb_result_q_reg_6_ ( .D(u_muldiv_N527), .CK(clk_i), .RN(
        n44157), .Q(writeback_muldiv_value_w[6]), .QN(n37633) );
  DFFRX1 u_muldiv_wb_result_q_reg_11_ ( .D(u_muldiv_N532), .CK(clk_i), .RN(
        n44157), .Q(writeback_muldiv_value_w[11]), .QN(n37609) );
  DFFRX1 u_muldiv_wb_result_q_reg_2_ ( .D(u_muldiv_N523), .CK(clk_i), .RN(
        n44157), .Q(writeback_muldiv_value_w[2]), .QN(n37629) );
  DFFRX1 u_muldiv_wb_result_q_reg_3_ ( .D(u_muldiv_N524), .CK(clk_i), .RN(
        n44156), .Q(writeback_muldiv_value_w[3]), .QN(n37630) );
  DFFRX1 u_muldiv_wb_result_q_reg_4_ ( .D(u_muldiv_N525), .CK(clk_i), .RN(
        n44156), .Q(writeback_muldiv_value_w[4]), .QN(n37631) );
  DFFRX1 u_muldiv_wb_result_q_reg_1_ ( .D(u_muldiv_N522), .CK(clk_i), .RN(
        n44156), .Q(writeback_muldiv_value_w[1]), .QN(n37601) );
  DFFRX1 u_muldiv_wb_result_q_reg_5_ ( .D(u_muldiv_N526), .CK(clk_i), .RN(
        n44156), .Q(writeback_muldiv_value_w[5]), .QN(n37632) );
  DFFRX1 u_muldiv_wb_result_q_reg_0_ ( .D(u_muldiv_N521), .CK(clk_i), .RN(
        n44156), .Q(writeback_muldiv_value_w[0]), .QN(n37600) );
  DFFRX1 u_muldiv_wb_result_q_reg_17_ ( .D(u_muldiv_N538), .CK(clk_i), .RN(
        n44156), .Q(writeback_muldiv_value_w[17]), .QN(n37615) );
  DFFRX1 u_muldiv_wb_result_q_reg_24_ ( .D(u_muldiv_N545), .CK(clk_i), .RN(
        n44156), .Q(writeback_muldiv_value_w[24]), .QN(n37621) );
  DFFRX1 u_muldiv_wb_result_q_reg_25_ ( .D(u_muldiv_N546), .CK(clk_i), .RN(
        n44156), .Q(writeback_muldiv_value_w[25]), .QN(n37622) );
  DFFRX1 u_muldiv_wb_result_q_reg_27_ ( .D(u_muldiv_N548), .CK(clk_i), .RN(
        n44156), .Q(writeback_muldiv_value_w[27]), .QN(n37624) );
  DFFRX1 u_muldiv_wb_result_q_reg_13_ ( .D(u_muldiv_N534), .CK(clk_i), .RN(
        n44156), .Q(writeback_muldiv_value_w[13]), .QN(n37611) );
  DFFRX1 u_muldiv_wb_result_q_reg_12_ ( .D(u_muldiv_N533), .CK(clk_i), .RN(
        n44156), .Q(writeback_muldiv_value_w[12]), .QN(n37610) );
  DFFRX1 u_muldiv_wb_result_q_reg_18_ ( .D(u_muldiv_N539), .CK(clk_i), .RN(
        n44156), .Q(writeback_muldiv_value_w[18]), .QN(n37616) );
  DFFRX1 u_muldiv_wb_result_q_reg_26_ ( .D(u_muldiv_N547), .CK(clk_i), .RN(
        n44156), .Q(writeback_muldiv_value_w[26]), .QN(n37623) );
  DFFRX1 u_muldiv_wb_result_q_reg_21_ ( .D(u_muldiv_N542), .CK(clk_i), .RN(
        n44156), .Q(writeback_muldiv_value_w[21]), .QN(n37618) );
  DFFRX1 u_muldiv_wb_result_q_reg_16_ ( .D(u_muldiv_N537), .CK(clk_i), .RN(
        n44156), .Q(writeback_muldiv_value_w[16]), .QN(n37614) );
  DFFRX1 u_muldiv_wb_result_q_reg_22_ ( .D(u_muldiv_N543), .CK(clk_i), .RN(
        n44156), .Q(writeback_muldiv_value_w[22]), .QN(n37619) );
  DFFRX1 u_muldiv_wb_result_q_reg_23_ ( .D(u_muldiv_N544), .CK(clk_i), .RN(
        n44156), .Q(writeback_muldiv_value_w[23]), .QN(n37620) );
  DFFRX1 u_muldiv_wb_result_q_reg_20_ ( .D(u_muldiv_N541), .CK(clk_i), .RN(
        n44156), .Q(writeback_muldiv_value_w[20]), .QN(n37599) );
  DFFRX1 u_muldiv_wb_result_q_reg_19_ ( .D(u_muldiv_N540), .CK(clk_i), .RN(
        n44155), .Q(writeback_muldiv_value_w[19]), .QN(n37617) );
  DFFRX1 u_muldiv_wb_result_q_reg_28_ ( .D(u_muldiv_N549), .CK(clk_i), .RN(
        n44155), .Q(writeback_muldiv_value_w[28]), .QN(n37625) );
  DFFRX1 u_muldiv_wb_result_q_reg_29_ ( .D(u_muldiv_N550), .CK(clk_i), .RN(
        n44155), .Q(writeback_muldiv_value_w[29]), .QN(n37626) );
  DFFRX1 u_muldiv_wb_result_q_reg_14_ ( .D(u_muldiv_N535), .CK(clk_i), .RN(
        n44155), .Q(writeback_muldiv_value_w[14]), .QN(n37612) );
  DFFRX1 u_muldiv_wb_result_q_reg_15_ ( .D(u_muldiv_N536), .CK(clk_i), .RN(
        n44155), .Q(writeback_muldiv_value_w[15]), .QN(n37613) );
  DFFRX1 u_muldiv_wb_result_q_reg_31_ ( .D(u_muldiv_N552), .CK(clk_i), .RN(
        n44155), .Q(writeback_muldiv_value_w[31]), .QN(n37628) );
  DFFRX1 u_muldiv_wb_result_q_reg_30_ ( .D(u_muldiv_N551), .CK(clk_i), .RN(
        n44155), .Q(writeback_muldiv_value_w[30]), .QN(n37627) );
  DFFRX1 u_csr_writeback_value_q_reg_8_ ( .D(u_csr_result_r[8]), .CK(net1857), 
        .RN(n44155), .Q(writeback_csr_value_w[8]), .QN(n37635) );
  DFFRX1 u_csr_writeback_value_q_reg_7_ ( .D(u_csr_result_r[7]), .CK(net1857), 
        .RN(n44159), .Q(writeback_csr_value_w[7]), .QN(n37634) );
  DFFRX1 u_csr_writeback_value_q_reg_9_ ( .D(u_csr_result_r[9]), .CK(net1857), 
        .RN(n44163), .Q(writeback_csr_value_w[9]), .QN(n37636) );
  DFFRX1 u_csr_writeback_value_q_reg_10_ ( .D(u_csr_result_r[10]), .CK(net1857), .RN(n44203), .Q(writeback_csr_value_w[10]), .QN(n37637) );
  DFFRX1 u_csr_writeback_value_q_reg_6_ ( .D(u_csr_result_r[6]), .CK(net1857), 
        .RN(n44203), .Q(writeback_csr_value_w[6]), .QN(n37662) );
  DFFRX1 u_csr_writeback_value_q_reg_11_ ( .D(u_csr_result_r[11]), .CK(net1857), .RN(n44203), .Q(writeback_csr_value_w[11]), .QN(n37638) );
  DFFRX1 u_csr_writeback_value_q_reg_5_ ( .D(u_csr_result_r[5]), .CK(net1857), 
        .RN(n44203), .Q(writeback_csr_value_w[5]), .QN(n37661) );
  DFFRX1 u_csr_writeback_value_q_reg_4_ ( .D(u_csr_result_r[4]), .CK(net1857), 
        .RN(n44203), .Q(writeback_csr_value_w[4]), .QN(n37660) );
  DFFRX1 u_csr_writeback_value_q_reg_3_ ( .D(u_csr_result_r[3]), .CK(net1857), 
        .RN(n44203), .Q(writeback_csr_value_w[3]), .QN(n37659) );
  DFFRX1 u_csr_writeback_value_q_reg_2_ ( .D(u_csr_result_r[2]), .CK(net1857), 
        .RN(n44203), .Q(writeback_csr_value_w[2]), .QN(n37658) );
  DFFRX1 u_csr_writeback_value_q_reg_1_ ( .D(u_csr_result_r[1]), .CK(net1857), 
        .RN(n44203), .Q(writeback_csr_value_w[1]), .QN(n37604) );
  DFFRX1 u_csr_writeback_value_q_reg_0_ ( .D(u_csr_result_r[0]), .CK(net1857), 
        .RN(n44202), .Q(writeback_csr_value_w[0]), .QN(n37603) );
  DFFRX1 u_csr_writeback_value_q_reg_31_ ( .D(u_csr_result_r[31]), .CK(net1862), .RN(n44202), .Q(writeback_csr_value_w[31]), .QN(n37657) );
  DFFRX1 u_csr_writeback_value_q_reg_17_ ( .D(u_csr_result_r[17]), .CK(net1862), .RN(n44202), .Q(writeback_csr_value_w[17]), .QN(n37644) );
  DFFRX1 u_csr_writeback_value_q_reg_24_ ( .D(u_csr_result_r[24]), .CK(net1862), .RN(n44202), .Q(writeback_csr_value_w[24]), .QN(n37650) );
  DFFRX1 u_csr_writeback_value_q_reg_25_ ( .D(u_csr_result_r[25]), .CK(net1862), .RN(n44202), .Q(writeback_csr_value_w[25]), .QN(n37651) );
  DFFRX1 u_csr_writeback_value_q_reg_27_ ( .D(u_csr_result_r[27]), .CK(net1862), .RN(n44202), .Q(writeback_csr_value_w[27]), .QN(n37653) );
  DFFRX1 u_csr_writeback_value_q_reg_13_ ( .D(u_csr_result_r[13]), .CK(net1857), .RN(n44202), .Q(writeback_csr_value_w[13]), .QN(n37640) );
  DFFRX1 u_csr_writeback_value_q_reg_12_ ( .D(u_csr_result_r[12]), .CK(net1857), .RN(n44202), .Q(writeback_csr_value_w[12]), .QN(n37639) );
  DFFRX1 u_csr_writeback_value_q_reg_18_ ( .D(u_csr_result_r[18]), .CK(net1862), .RN(n44202), .Q(writeback_csr_value_w[18]), .QN(n37645) );
  DFFRX1 u_csr_writeback_value_q_reg_26_ ( .D(u_csr_result_r[26]), .CK(net1862), .RN(n44202), .Q(writeback_csr_value_w[26]), .QN(n37652) );
  DFFRX1 u_csr_writeback_value_q_reg_21_ ( .D(u_csr_result_r[21]), .CK(net1862), .RN(n44202), .Q(writeback_csr_value_w[21]), .QN(n37647) );
  DFFRX1 u_csr_writeback_value_q_reg_16_ ( .D(u_csr_result_r[16]), .CK(net1862), .RN(n44202), .Q(writeback_csr_value_w[16]), .QN(n37643) );
  DFFRX1 u_csr_writeback_value_q_reg_22_ ( .D(u_csr_result_r[22]), .CK(net1862), .RN(n44202), .Q(writeback_csr_value_w[22]), .QN(n37648) );
  DFFRX1 u_csr_writeback_value_q_reg_23_ ( .D(u_csr_result_r[23]), .CK(net1862), .RN(n44202), .Q(writeback_csr_value_w[23]), .QN(n37649) );
  DFFRX1 u_csr_writeback_value_q_reg_20_ ( .D(u_csr_result_r[20]), .CK(net1862), .RN(n44202), .Q(writeback_csr_value_w[20]), .QN(n37602) );
  DFFRX1 u_csr_writeback_value_q_reg_19_ ( .D(u_csr_result_r[19]), .CK(net1862), .RN(n44202), .Q(writeback_csr_value_w[19]), .QN(n37646) );
  DFFRX1 u_csr_writeback_value_q_reg_28_ ( .D(u_csr_result_r[28]), .CK(net1862), .RN(n44202), .Q(writeback_csr_value_w[28]), .QN(n37654) );
  DFFRX1 u_csr_writeback_value_q_reg_29_ ( .D(u_csr_result_r[29]), .CK(net1862), .RN(n44202), .Q(writeback_csr_value_w[29]), .QN(n37655) );
  DFFRX1 u_csr_writeback_value_q_reg_14_ ( .D(u_csr_result_r[14]), .CK(net1857), .RN(n44201), .Q(writeback_csr_value_w[14]), .QN(n37641) );
  DFFRX1 u_csr_writeback_value_q_reg_15_ ( .D(u_csr_result_r[15]), .CK(net1857), .RN(n44201), .Q(writeback_csr_value_w[15]), .QN(n37642) );
  DFFRX1 u_csr_writeback_value_q_reg_30_ ( .D(u_csr_result_r[30]), .CK(net1862), .RN(n44201), .Q(writeback_csr_value_w[30]), .QN(n37656) );
  DFFRX1 u_csr_pc_m_q_reg_2_ ( .D(opcode_pc_w[2]), .CK(net1867), .RN(n44116), 
        .Q(n3064) );
  DFFRX1 u_csr_pc_m_q_reg_3_ ( .D(opcode_pc_w[3]), .CK(net1867), .RN(n44117), 
        .QN(n37764) );
  DFFSHQX1 u_csr_reset_q_reg ( .D(1'b0), .CK(clk_i), .SN(n44087), .Q(n8572) );
  DFFSHQX1 u_csr_csr_mpriv_q_reg_1_ ( .D(n36340), .CK(clk_i), .SN(n44087), .Q(
        u_csr_N3162) );
  DFFSHQX1 u_csr_csr_mpriv_q_reg_0_ ( .D(n36341), .CK(clk_i), .SN(n44087), .Q(
        u_csr_N3161) );
  INVX1 U4 ( .A(n8572), .Y(n8805) );
  INVX1 U52 ( .A(n16954), .Y(n48) );
  INVX1 U53 ( .A(n15627), .Y(n49) );
  INVX1 U54 ( .A(n15735), .Y(n50) );
  INVX1 U55 ( .A(n16351), .Y(n51) );
  INVX1 U56 ( .A(n16407), .Y(n52) );
  INVX1 U57 ( .A(n15884), .Y(n53) );
  INVX1 U58 ( .A(n15887), .Y(n54) );
  INVX1 U59 ( .A(n16299), .Y(n55) );
  INVX1 U183 ( .A(n16298), .Y(n179) );
  INVX1 U184 ( .A(n16233), .Y(n180) );
  INVX1 U219 ( .A(n15501), .Y(n215) );
  INVX1 U220 ( .A(n16961), .Y(n216) );
  INVX1 U230 ( .A(n17106), .Y(n226) );
  INVX1 U231 ( .A(n16910), .Y(n227) );
  INVX1 U233 ( .A(n15836), .Y(n229) );
  INVX1 U259 ( .A(n16958), .Y(n255) );
  INVX1 U260 ( .A(n16864), .Y(n256) );
  INVX1 U261 ( .A(n16640), .Y(n257) );
  INVX1 U304 ( .A(n16165), .Y(n300) );
  INVX1 U313 ( .A(n16234), .Y(n309) );
  INVX1 U344 ( .A(n15404), .Y(n340) );
  INVX1 U372 ( .A(n15965), .Y(n368) );
  INVX1 U373 ( .A(n15829), .Y(n369) );
  INVX1 U375 ( .A(n15966), .Y(n371) );
  INVX1 U377 ( .A(mem_d_data_rd_i[28]), .Y(n373) );
  INVX1 U379 ( .A(n27352), .Y(n375) );
  INVX1 U382 ( .A(n16113), .Y(n378) );
  INVX1 U388 ( .A(mem_d_data_rd_i[27]), .Y(n384) );
  INVX1 U392 ( .A(n25699), .Y(n388) );
  INVX1 U395 ( .A(n26959), .Y(n391) );
  INVX1 U399 ( .A(mem_d_data_rd_i[26]), .Y(n395) );
  INVX1 U414 ( .A(n26978), .Y(n410) );
  INVX1 U415 ( .A(n26331), .Y(n411) );
  INVX1 U433 ( .A(mem_d_data_rd_i[15]), .Y(n429) );
  INVX1 U434 ( .A(mem_d_data_rd_i[9]), .Y(n430) );
  INVX1 U435 ( .A(mem_d_data_rd_i[8]), .Y(n431) );
  INVX1 U436 ( .A(mem_d_data_rd_i[4]), .Y(n432) );
  INVX1 U440 ( .A(mem_d_data_rd_i[3]), .Y(n436) );
  INVX1 U441 ( .A(mem_d_data_rd_i[2]), .Y(n437) );
  INVX1 U442 ( .A(mem_d_data_rd_i[1]), .Y(n438) );
  INVX1 U444 ( .A(mem_d_accept_i), .Y(n440) );
  INVX1 U445 ( .A(u_muldiv_N264), .Y(n441) );
  INVX1 U455 ( .A(n26917), .Y(n451) );
  INVX1 U461 ( .A(n40682), .Y(n457) );
  INVX1 U462 ( .A(n25409), .Y(n458) );
  INVX1 U463 ( .A(n26294), .Y(n459) );
  INVX1 U465 ( .A(n27390), .Y(n461) );
  INVX1 U466 ( .A(n26913), .Y(n462) );
  INVX1 U467 ( .A(n28515), .Y(n463) );
  INVX1 U469 ( .A(n28163), .Y(n465) );
  INVX1 U470 ( .A(n28032), .Y(n466) );
  INVX1 U473 ( .A(n26272), .Y(n469) );
  INVX1 U474 ( .A(n26285), .Y(n470) );
  INVX1 U491 ( .A(mem_d_ack_i), .Y(n487) );
  INVX1 U495 ( .A(n29231), .Y(n491) );
  INVX1 U496 ( .A(n21240), .Y(n492) );
  INVX1 U498 ( .A(n29248), .Y(n494) );
  INVX1 U500 ( .A(n29281), .Y(n496) );
  INVX1 U502 ( .A(n29264), .Y(n498) );
  INVX1 U506 ( .A(n29240), .Y(n502) );
  INVX1 U508 ( .A(n29273), .Y(n504) );
  INVX1 U516 ( .A(n29294), .Y(n512) );
  INVX1 U517 ( .A(n19867), .Y(n513) );
  INVX1 U521 ( .A(n29107), .Y(n517) );
  INVX1 U522 ( .A(n24101), .Y(n518) );
  INVX1 U523 ( .A(n29304), .Y(n519) );
  INVX1 U524 ( .A(n19670), .Y(n520) );
  INVX1 U527 ( .A(n29085), .Y(n523) );
  INVX1 U528 ( .A(n18296), .Y(n524) );
  INVX1 U530 ( .A(n29162), .Y(n526) );
  INVX1 U532 ( .A(n29182), .Y(n528) );
  INVX1 U534 ( .A(n29203), .Y(n530) );
  INVX1 U538 ( .A(n29339), .Y(n534) );
  INVX1 U542 ( .A(n29033), .Y(n538) );
  INVX1 U544 ( .A(n19475), .Y(n540) );
  INVX1 U545 ( .A(n19472), .Y(n541) );
  INVX1 U546 ( .A(n29316), .Y(n542) );
  INVX1 U548 ( .A(n29129), .Y(n544) );
  INVX1 U550 ( .A(n29047), .Y(n546) );
  INVX1 U552 ( .A(n29099), .Y(n548) );
  INVX1 U554 ( .A(n29073), .Y(n550) );
  INVX1 U555 ( .A(n29118), .Y(n551) );
  INVX1 U557 ( .A(n24179), .Y(n553) );
  INVX1 U558 ( .A(n29139), .Y(n554) );
  INVX1 U562 ( .A(n29349), .Y(n558) );
  INVX1 U566 ( .A(n29328), .Y(n562) );
  INVX1 U568 ( .A(n29059), .Y(n564) );
  INVX1 U570 ( .A(n29173), .Y(n566) );
  INVX1 U573 ( .A(n24134), .Y(n569) );
  INVX1 U574 ( .A(n29212), .Y(n570) );
  INVX1 U576 ( .A(n29193), .Y(n572) );
  INVX1 U579 ( .A(mem_d_error_i), .Y(n575) );
  INVX1 U580 ( .A(mem_d_resp_tag_i[9]), .Y(n576) );
  INVX1 U581 ( .A(n33678), .Y(n577) );
  INVX1 U585 ( .A(n33681), .Y(n581) );
  INVX1 U586 ( .A(mem_d_resp_tag_i[8]), .Y(n582) );
  INVX1 U587 ( .A(n33543), .Y(n583) );
  INVX1 U588 ( .A(n32009), .Y(n584) );
  INVX1 U589 ( .A(mem_d_resp_tag_i[7]), .Y(n585) );
  INVX1 U590 ( .A(mem_d_resp_tag_i[6]), .Y(n586) );
  INVX1 U591 ( .A(mem_d_resp_tag_i[5]), .Y(n587) );
  INVX1 U600 ( .A(n24440), .Y(n596) );
  INVX1 U615 ( .A(n24574), .Y(n611) );
  INVX1 U616 ( .A(n24573), .Y(n612) );
  INVX1 U659 ( .A(n28102), .Y(n655) );
  INVX1 U696 ( .A(n28735), .Y(n692) );
  INVX1 U701 ( .A(mem_d_addr_o[28]), .Y(n697) );
  INVX1 U712 ( .A(n14474), .Y(n708) );
  INVX1 U713 ( .A(n13846), .Y(n709) );
  INVX1 U714 ( .A(n14137), .Y(n710) );
  INVX1 U716 ( .A(n14127), .Y(n712) );
  INVX1 U717 ( .A(n14468), .Y(n713) );
  INVX1 U718 ( .A(n14473), .Y(n714) );
  INVX1 U719 ( .A(n14488), .Y(n715) );
  INVX1 U720 ( .A(n14502), .Y(n716) );
  INVX1 U721 ( .A(n14516), .Y(n717) );
  INVX1 U722 ( .A(n14544), .Y(n718) );
  INVX1 U723 ( .A(n14558), .Y(n719) );
  INVX1 U724 ( .A(n14572), .Y(n720) );
  INVX1 U725 ( .A(n14600), .Y(n721) );
  INVX1 U726 ( .A(n14614), .Y(n722) );
  INVX1 U727 ( .A(n14628), .Y(n723) );
  INVX1 U728 ( .A(n14656), .Y(n724) );
  INVX1 U729 ( .A(n14670), .Y(n725) );
  INVX1 U730 ( .A(n14684), .Y(n726) );
  INVX1 U731 ( .A(n14712), .Y(n727) );
  INVX1 U732 ( .A(n14726), .Y(n728) );
  INVX1 U733 ( .A(n14740), .Y(n729) );
  INVX1 U734 ( .A(n14768), .Y(n730) );
  INVX1 U735 ( .A(n14782), .Y(n731) );
  INVX1 U736 ( .A(n14796), .Y(n732) );
  INVX1 U768 ( .A(n13987), .Y(n764) );
  INVX1 U803 ( .A(n14005), .Y(n799) );
  INVX1 U809 ( .A(u_muldiv_dividend_q[28]), .Y(n805) );
  INVX1 U821 ( .A(n14119), .Y(n817) );
  INVX1 U837 ( .A(n14101), .Y(n833) );
  INVX1 U851 ( .A(n14164), .Y(n847) );
  INVX1 U852 ( .A(n14163), .Y(n848) );
  INVX1 U853 ( .A(n14162), .Y(n849) );
  INVX1 U854 ( .A(n14161), .Y(n850) );
  INVX1 U855 ( .A(n14160), .Y(n851) );
  INVX1 U856 ( .A(n14159), .Y(n852) );
  INVX1 U857 ( .A(n14158), .Y(n853) );
  INVX1 U858 ( .A(n14157), .Y(n854) );
  INVX1 U859 ( .A(n14156), .Y(n855) );
  INVX1 U860 ( .A(n14155), .Y(n856) );
  INVX1 U861 ( .A(n14154), .Y(n857) );
  INVX1 U862 ( .A(n14153), .Y(n858) );
  INVX1 U863 ( .A(n14152), .Y(n859) );
  INVX1 U864 ( .A(n14151), .Y(n860) );
  INVX1 U865 ( .A(n14150), .Y(n861) );
  INVX1 U866 ( .A(n14149), .Y(n862) );
  INVX1 U867 ( .A(n14148), .Y(n863) );
  INVX1 U872 ( .A(n14081), .Y(n868) );
  INVX1 U873 ( .A(n14063), .Y(n869) );
  INVX1 U874 ( .A(n14043), .Y(n870) );
  INVX1 U875 ( .A(n14025), .Y(n871) );
  INVX1 U876 ( .A(n13967), .Y(n872) );
  INVX1 U877 ( .A(n13949), .Y(n873) );
  INVX1 U878 ( .A(n13929), .Y(n874) );
  INVX1 U879 ( .A(n13911), .Y(n875) );
  INVX1 U880 ( .A(n13891), .Y(n876) );
  INVX1 U881 ( .A(n13873), .Y(n877) );
  INVX1 U887 ( .A(n28214), .Y(n883) );
  INVX1 U888 ( .A(n27370), .Y(n884) );
  INVX1 U889 ( .A(n27371), .Y(n885) );
  INVX1 U977 ( .A(n27096), .Y(n973) );
  INVX1 U984 ( .A(n42968), .Y(n980) );
  INVX1 U1058 ( .A(n24231), .Y(n1054) );
  INVX1 U1061 ( .A(n29275), .Y(n1057) );
  INVX1 U1066 ( .A(n29040), .Y(n1062) );
  INVX1 U1067 ( .A(n29283), .Y(n1063) );
  INVX1 U1069 ( .A(n29214), .Y(n1065) );
  INVX1 U1086 ( .A(n28166), .Y(n1082) );
  INVX1 U1087 ( .A(n28175), .Y(n1083) );
  INVX1 U1089 ( .A(n28195), .Y(n1085) );
  INVX1 U1090 ( .A(n29591), .Y(n1086) );
  INVX1 U1141 ( .A(u_csr_csr_sscratch_q[6]), .Y(n1137) );
  INVX1 U1142 ( .A(u_csr_csr_sscratch_q[5]), .Y(n1138) );
  INVX1 U1143 ( .A(u_csr_csr_sscratch_q[4]), .Y(n1139) );
  INVX1 U1144 ( .A(u_csr_csr_sscratch_q[3]), .Y(n1140) );
  INVX1 U1145 ( .A(u_csr_csr_sscratch_q[31]), .Y(n1141) );
  INVX1 U1146 ( .A(u_csr_csr_sscratch_q[30]), .Y(n1142) );
  INVX1 U1147 ( .A(u_csr_csr_sscratch_q[2]), .Y(n1143) );
  INVX1 U1148 ( .A(u_csr_csr_sscratch_q[29]), .Y(n1144) );
  INVX1 U1149 ( .A(u_csr_csr_sscratch_q[28]), .Y(n1145) );
  INVX1 U1150 ( .A(u_csr_csr_sscratch_q[27]), .Y(n1146) );
  INVX1 U1151 ( .A(u_csr_csr_sscratch_q[26]), .Y(n1147) );
  INVX1 U1152 ( .A(u_csr_csr_sscratch_q[25]), .Y(n1148) );
  INVX1 U1153 ( .A(u_csr_csr_sscratch_q[24]), .Y(n1149) );
  INVX1 U1154 ( .A(u_csr_csr_sscratch_q[23]), .Y(n1150) );
  INVX1 U1155 ( .A(u_csr_csr_sscratch_q[22]), .Y(n1151) );
  INVX1 U1156 ( .A(u_csr_csr_sscratch_q[21]), .Y(n1152) );
  INVX1 U1157 ( .A(u_csr_csr_sscratch_q[20]), .Y(n1153) );
  INVX1 U1158 ( .A(u_csr_csr_sscratch_q[1]), .Y(n1154) );
  INVX1 U1159 ( .A(u_csr_csr_sscratch_q[19]), .Y(n1155) );
  INVX1 U1160 ( .A(u_csr_csr_sscratch_q[18]), .Y(n1156) );
  INVX1 U1161 ( .A(u_csr_csr_sscratch_q[17]), .Y(n1157) );
  INVX1 U1162 ( .A(u_csr_csr_sscratch_q[16]), .Y(n1158) );
  INVX1 U1163 ( .A(u_csr_csr_sscratch_q[15]), .Y(n1159) );
  INVX1 U1164 ( .A(u_csr_csr_sscratch_q[14]), .Y(n1160) );
  INVX1 U1165 ( .A(u_csr_csr_sscratch_q[13]), .Y(n1161) );
  INVX1 U1166 ( .A(u_csr_csr_sscratch_q[12]), .Y(n1162) );
  INVX1 U1167 ( .A(u_csr_csr_sscratch_q[10]), .Y(n1163) );
  INVX1 U1168 ( .A(u_csr_csr_sscratch_q[0]), .Y(n1164) );
  INVX1 U1169 ( .A(u_csr_csr_stvec_q[9]), .Y(n1165) );
  INVX1 U1170 ( .A(u_csr_csr_stvec_q[8]), .Y(n1166) );
  INVX1 U1171 ( .A(u_csr_csr_stvec_q[7]), .Y(n1167) );
  INVX1 U1172 ( .A(u_csr_csr_stvec_q[6]), .Y(n1168) );
  INVX1 U1173 ( .A(u_csr_csr_stvec_q[5]), .Y(n1169) );
  INVX1 U1176 ( .A(u_csr_csr_stvec_q[31]), .Y(n1172) );
  INVX1 U1177 ( .A(u_csr_csr_stvec_q[30]), .Y(n1173) );
  INVX1 U1179 ( .A(u_csr_csr_stvec_q[29]), .Y(n1175) );
  INVX1 U1180 ( .A(u_csr_csr_stvec_q[28]), .Y(n1176) );
  INVX1 U1181 ( .A(u_csr_csr_stvec_q[27]), .Y(n1177) );
  INVX1 U1182 ( .A(u_csr_csr_stvec_q[26]), .Y(n1178) );
  INVX1 U1183 ( .A(u_csr_csr_stvec_q[25]), .Y(n1179) );
  INVX1 U1184 ( .A(u_csr_csr_stvec_q[24]), .Y(n1180) );
  INVX1 U1185 ( .A(u_csr_csr_stvec_q[23]), .Y(n1181) );
  INVX1 U1186 ( .A(u_csr_csr_stvec_q[22]), .Y(n1182) );
  INVX1 U1187 ( .A(u_csr_csr_stvec_q[21]), .Y(n1183) );
  INVX1 U1188 ( .A(u_csr_csr_stvec_q[20]), .Y(n1184) );
  INVX1 U1190 ( .A(u_csr_csr_stvec_q[19]), .Y(n1186) );
  INVX1 U1191 ( .A(u_csr_csr_stvec_q[18]), .Y(n1187) );
  INVX1 U1192 ( .A(u_csr_csr_stvec_q[17]), .Y(n1188) );
  INVX1 U1193 ( .A(u_csr_csr_stvec_q[16]), .Y(n1189) );
  INVX1 U1194 ( .A(u_csr_csr_stvec_q[15]), .Y(n1190) );
  INVX1 U1195 ( .A(u_csr_csr_stvec_q[14]), .Y(n1191) );
  INVX1 U1196 ( .A(u_csr_csr_stvec_q[13]), .Y(n1192) );
  INVX1 U1197 ( .A(u_csr_csr_stvec_q[12]), .Y(n1193) );
  INVX1 U1198 ( .A(u_csr_csr_stvec_q[10]), .Y(n1194) );
  INVX1 U1228 ( .A(u_csr_csr_sscratch_q[11]), .Y(n1224) );
  INVX1 U1229 ( .A(u_csr_csr_stvec_q[11]), .Y(n1225) );
  INVX1 U1413 ( .A(u_muldiv_dividend_q[19]), .Y(n1409) );
  INVX1 U1443 ( .A(u_muldiv_dividend_q[20]), .Y(n1439) );
  INVX1 U1463 ( .A(u_muldiv_dividend_q[23]), .Y(n1459) );
  INVX1 U1475 ( .A(u_muldiv_dividend_q[22]), .Y(n1471) );
  INVX1 U1515 ( .A(u_muldiv_dividend_q[26]), .Y(n1511) );
  INVX1 U1565 ( .A(u_muldiv_dividend_q[27]), .Y(n1561) );
  INVX1 U1586 ( .A(u_muldiv_dividend_q[24]), .Y(n1582) );
  INVX1 U1633 ( .A(u_muldiv_divisor_q[60]), .Y(n1629) );
  INVX1 U1634 ( .A(u_muldiv_dividend_q[29]), .Y(n1630) );
  INVX1 U1755 ( .A(n8805), .Y(n1751) );
  NAND2X1 U8905 ( .A(n10607), .B(n10608), .Y(u_muldiv_result_r[0]) );
  NAND2X1 U12310 ( .A(n13840), .B(n13841), .Y(u_muldiv_N552) );
  NOR2X1 U12312 ( .A(n13843), .B(n13844), .Y(n13840) );
  AND2X1 U12313 ( .A(n13845), .B(n13846), .Y(n13844) );
  NOR2X1 U12314 ( .A(n13847), .B(n44630), .Y(n13843) );
  XNOR2X1 U12315 ( .A(n13845), .B(n13849), .Y(n13847) );
  NAND2X1 U12316 ( .A(n13850), .B(n13851), .Y(n13849) );
  NAND2X1 U12317 ( .A(n13852), .B(n13853), .Y(n13845) );
  NAND2X1 U12318 ( .A(u_muldiv_dividend_q[31]), .B(n37586), .Y(n13853) );
  NAND2X1 U12319 ( .A(u_muldiv_quotient_q[31]), .B(n44823), .Y(n13852) );
  NAND2X1 U12320 ( .A(n13854), .B(n13855), .Y(u_muldiv_N551) );
  NOR2X1 U12322 ( .A(n13856), .B(n13857), .Y(n13854) );
  NOR2X1 U12323 ( .A(n13850), .B(n709), .Y(n13857) );
  NOR2X1 U12324 ( .A(n13858), .B(n44630), .Y(n13856) );
  XNOR2X1 U12325 ( .A(n13850), .B(n13851), .Y(n13858) );
  NOR2X1 U12326 ( .A(n13859), .B(n13860), .Y(n13851) );
  AND2X1 U12327 ( .A(n13861), .B(n13862), .Y(n13850) );
  NAND2X1 U12328 ( .A(u_muldiv_dividend_q[30]), .B(n37586), .Y(n13862) );
  NAND2X1 U12329 ( .A(u_muldiv_quotient_q[30]), .B(n44823), .Y(n13861) );
  NAND2X1 U12330 ( .A(n13863), .B(n13864), .Y(u_muldiv_N550) );
  NOR2X1 U12332 ( .A(n13865), .B(n13866), .Y(n13863) );
  AND2X1 U12333 ( .A(n13860), .B(n13846), .Y(n13866) );
  NOR2X1 U12334 ( .A(n13867), .B(n44630), .Y(n13865) );
  XNOR2X1 U12335 ( .A(n13859), .B(n13860), .Y(n13867) );
  NAND2X1 U12336 ( .A(n13868), .B(n13869), .Y(n13860) );
  NAND2X1 U12337 ( .A(u_muldiv_dividend_q[29]), .B(n37586), .Y(n13869) );
  NAND2X1 U12338 ( .A(u_muldiv_quotient_q[29]), .B(n44823), .Y(n13868) );
  NAND2X1 U12339 ( .A(n13870), .B(n13871), .Y(n13859) );
  NOR2X1 U12340 ( .A(n13872), .B(n13873), .Y(n13870) );
  NAND2X1 U12341 ( .A(n13874), .B(n13875), .Y(u_muldiv_N549) );
  NOR2X1 U12343 ( .A(n13876), .B(n13877), .Y(n13874) );
  AND2X1 U12344 ( .A(n13872), .B(n13846), .Y(n13877) );
  NOR2X1 U12345 ( .A(n13878), .B(n44630), .Y(n13876) );
  XNOR2X1 U12346 ( .A(n13872), .B(n13879), .Y(n13878) );
  NAND2X1 U12347 ( .A(n13871), .B(n877), .Y(n13879) );
  NAND2X1 U12348 ( .A(n13880), .B(n13881), .Y(n13872) );
  NAND2X1 U12349 ( .A(u_muldiv_dividend_q[28]), .B(n37586), .Y(n13881) );
  NAND2X1 U12350 ( .A(u_muldiv_quotient_q[28]), .B(n44823), .Y(n13880) );
  NAND2X1 U12351 ( .A(n13882), .B(n13883), .Y(u_muldiv_N548) );
  NOR2X1 U12353 ( .A(n13884), .B(n13885), .Y(n13882) );
  NOR2X1 U12354 ( .A(n877), .B(n709), .Y(n13885) );
  NOR2X1 U12355 ( .A(n13886), .B(n44629), .Y(n13884) );
  XNOR2X1 U12356 ( .A(n13871), .B(n877), .Y(n13886) );
  NAND2X1 U12357 ( .A(n13887), .B(n13888), .Y(n13873) );
  NAND2X1 U12358 ( .A(u_muldiv_dividend_q[27]), .B(n37586), .Y(n13888) );
  NAND2X1 U12359 ( .A(u_muldiv_quotient_q[27]), .B(n44823), .Y(n13887) );
  NOR2X1 U12360 ( .A(n13889), .B(n13890), .Y(n13871) );
  OR2X1 U12361 ( .A(n13891), .B(n13892), .Y(n13889) );
  NAND2X1 U12362 ( .A(n13893), .B(n13894), .Y(u_muldiv_N547) );
  NOR2X1 U12364 ( .A(n13895), .B(n13896), .Y(n13893) );
  NOR2X1 U12365 ( .A(n876), .B(n709), .Y(n13896) );
  NOR2X1 U12366 ( .A(n13897), .B(n44629), .Y(n13895) );
  XNOR2X1 U12367 ( .A(n876), .B(n13898), .Y(n13897) );
  NOR2X1 U12368 ( .A(n13892), .B(n13890), .Y(n13898) );
  NAND2X1 U12369 ( .A(n13899), .B(n13900), .Y(n13891) );
  NAND2X1 U12370 ( .A(u_muldiv_dividend_q[26]), .B(n37586), .Y(n13900) );
  NAND2X1 U12371 ( .A(u_muldiv_quotient_q[26]), .B(n44823), .Y(n13899) );
  NAND2X1 U12372 ( .A(n13901), .B(n13902), .Y(u_muldiv_N546) );
  NOR2X1 U12374 ( .A(n13903), .B(n13904), .Y(n13901) );
  AND2X1 U12375 ( .A(n13892), .B(n13846), .Y(n13904) );
  NOR2X1 U12376 ( .A(n13905), .B(n44629), .Y(n13903) );
  XNOR2X1 U12377 ( .A(n13890), .B(n13892), .Y(n13905) );
  NAND2X1 U12378 ( .A(n13906), .B(n13907), .Y(n13892) );
  NAND2X1 U12379 ( .A(u_muldiv_dividend_q[25]), .B(n44824), .Y(n13907) );
  NAND2X1 U12380 ( .A(u_muldiv_quotient_q[25]), .B(n44823), .Y(n13906) );
  NAND2X1 U12381 ( .A(n13908), .B(n13909), .Y(n13890) );
  NOR2X1 U12382 ( .A(n13910), .B(n13911), .Y(n13908) );
  NAND2X1 U12383 ( .A(n13912), .B(n13913), .Y(u_muldiv_N545) );
  NOR2X1 U12385 ( .A(n13914), .B(n13915), .Y(n13912) );
  AND2X1 U12386 ( .A(n13910), .B(n13846), .Y(n13915) );
  NOR2X1 U12387 ( .A(n13916), .B(n44629), .Y(n13914) );
  XNOR2X1 U12388 ( .A(n13910), .B(n13917), .Y(n13916) );
  NAND2X1 U12389 ( .A(n13909), .B(n875), .Y(n13917) );
  NAND2X1 U12390 ( .A(n13918), .B(n13919), .Y(n13910) );
  NAND2X1 U12391 ( .A(u_muldiv_dividend_q[24]), .B(n44824), .Y(n13919) );
  NAND2X1 U12392 ( .A(u_muldiv_quotient_q[24]), .B(n44823), .Y(n13918) );
  NAND2X1 U12393 ( .A(n13920), .B(n13921), .Y(u_muldiv_N544) );
  NOR2X1 U12395 ( .A(n13922), .B(n13923), .Y(n13920) );
  NOR2X1 U12396 ( .A(n875), .B(n709), .Y(n13923) );
  NOR2X1 U12397 ( .A(n13924), .B(n44629), .Y(n13922) );
  XNOR2X1 U12398 ( .A(n13909), .B(n875), .Y(n13924) );
  NAND2X1 U12399 ( .A(n13925), .B(n13926), .Y(n13911) );
  NAND2X1 U12400 ( .A(u_muldiv_dividend_q[23]), .B(n44824), .Y(n13926) );
  NAND2X1 U12401 ( .A(u_muldiv_quotient_q[23]), .B(n44822), .Y(n13925) );
  NOR2X1 U12402 ( .A(n13927), .B(n13928), .Y(n13909) );
  OR2X1 U12403 ( .A(n13929), .B(n13930), .Y(n13927) );
  NAND2X1 U12404 ( .A(n13931), .B(n13932), .Y(u_muldiv_N543) );
  NOR2X1 U12406 ( .A(n13933), .B(n13934), .Y(n13931) );
  NOR2X1 U12407 ( .A(n874), .B(n709), .Y(n13934) );
  NOR2X1 U12408 ( .A(n13935), .B(n44629), .Y(n13933) );
  XNOR2X1 U12409 ( .A(n874), .B(n13936), .Y(n13935) );
  NOR2X1 U12410 ( .A(n13930), .B(n13928), .Y(n13936) );
  NAND2X1 U12411 ( .A(n13937), .B(n13938), .Y(n13929) );
  NAND2X1 U12412 ( .A(u_muldiv_dividend_q[22]), .B(n44825), .Y(n13938) );
  NAND2X1 U12413 ( .A(u_muldiv_quotient_q[22]), .B(n44822), .Y(n13937) );
  NAND2X1 U12414 ( .A(n13939), .B(n13940), .Y(u_muldiv_N542) );
  NOR2X1 U12416 ( .A(n13941), .B(n13942), .Y(n13939) );
  AND2X1 U12417 ( .A(n13930), .B(n13846), .Y(n13942) );
  NOR2X1 U12418 ( .A(n13943), .B(n44629), .Y(n13941) );
  XNOR2X1 U12419 ( .A(n13928), .B(n13930), .Y(n13943) );
  NAND2X1 U12420 ( .A(n13944), .B(n13945), .Y(n13930) );
  NAND2X1 U12421 ( .A(u_muldiv_dividend_q[21]), .B(n44825), .Y(n13945) );
  NAND2X1 U12422 ( .A(u_muldiv_quotient_q[21]), .B(n44822), .Y(n13944) );
  NAND2X1 U12423 ( .A(n13946), .B(n13947), .Y(n13928) );
  NOR2X1 U12424 ( .A(n13948), .B(n13949), .Y(n13946) );
  NAND2X1 U12425 ( .A(n13950), .B(n13951), .Y(u_muldiv_N541) );
  NOR2X1 U12427 ( .A(n13952), .B(n13953), .Y(n13950) );
  AND2X1 U12428 ( .A(n13948), .B(n13846), .Y(n13953) );
  NOR2X1 U12429 ( .A(n13954), .B(n44629), .Y(n13952) );
  XNOR2X1 U12430 ( .A(n13948), .B(n13955), .Y(n13954) );
  NAND2X1 U12431 ( .A(n13947), .B(n873), .Y(n13955) );
  NAND2X1 U12432 ( .A(n13956), .B(n13957), .Y(n13948) );
  NAND2X1 U12433 ( .A(u_muldiv_dividend_q[20]), .B(n44825), .Y(n13957) );
  NAND2X1 U12434 ( .A(u_muldiv_quotient_q[20]), .B(n44822), .Y(n13956) );
  NAND2X1 U12435 ( .A(n13958), .B(n13959), .Y(u_muldiv_N540) );
  NOR2X1 U12437 ( .A(n13960), .B(n13961), .Y(n13958) );
  NOR2X1 U12438 ( .A(n873), .B(n709), .Y(n13961) );
  NOR2X1 U12439 ( .A(n13962), .B(n44629), .Y(n13960) );
  XNOR2X1 U12440 ( .A(n13947), .B(n873), .Y(n13962) );
  NAND2X1 U12441 ( .A(n13963), .B(n13964), .Y(n13949) );
  NAND2X1 U12442 ( .A(u_muldiv_dividend_q[19]), .B(n44826), .Y(n13964) );
  NAND2X1 U12443 ( .A(u_muldiv_quotient_q[19]), .B(n44822), .Y(n13963) );
  NOR2X1 U12444 ( .A(n13965), .B(n13966), .Y(n13947) );
  OR2X1 U12445 ( .A(n13967), .B(n13968), .Y(n13965) );
  NAND2X1 U12446 ( .A(n13969), .B(n13970), .Y(u_muldiv_N539) );
  NOR2X1 U12448 ( .A(n13971), .B(n13972), .Y(n13969) );
  NOR2X1 U12449 ( .A(n872), .B(n709), .Y(n13972) );
  NOR2X1 U12450 ( .A(n13973), .B(n44629), .Y(n13971) );
  XNOR2X1 U12451 ( .A(n872), .B(n13974), .Y(n13973) );
  NOR2X1 U12452 ( .A(n13968), .B(n13966), .Y(n13974) );
  NAND2X1 U12453 ( .A(n13975), .B(n13976), .Y(n13967) );
  NAND2X1 U12454 ( .A(u_muldiv_dividend_q[18]), .B(n44826), .Y(n13976) );
  NAND2X1 U12455 ( .A(u_muldiv_quotient_q[18]), .B(n44822), .Y(n13975) );
  NAND2X1 U12456 ( .A(n13977), .B(n13978), .Y(u_muldiv_N538) );
  NOR2X1 U12458 ( .A(n13979), .B(n13980), .Y(n13977) );
  AND2X1 U12459 ( .A(n13968), .B(n13846), .Y(n13980) );
  NOR2X1 U12460 ( .A(n13981), .B(n44629), .Y(n13979) );
  XNOR2X1 U12461 ( .A(n13966), .B(n13968), .Y(n13981) );
  NAND2X1 U12462 ( .A(n13982), .B(n13983), .Y(n13968) );
  NAND2X1 U12463 ( .A(u_muldiv_dividend_q[17]), .B(n44826), .Y(n13983) );
  NAND2X1 U12464 ( .A(u_muldiv_quotient_q[17]), .B(n44822), .Y(n13982) );
  NAND2X1 U12465 ( .A(n13984), .B(n13985), .Y(n13966) );
  NOR2X1 U12466 ( .A(n13986), .B(n13987), .Y(n13984) );
  NAND2X1 U12467 ( .A(n13988), .B(n13989), .Y(u_muldiv_N537) );
  NOR2X1 U12469 ( .A(n13990), .B(n13991), .Y(n13988) );
  AND2X1 U12470 ( .A(n13986), .B(n13846), .Y(n13991) );
  NOR2X1 U12471 ( .A(n13992), .B(n44629), .Y(n13990) );
  XNOR2X1 U12472 ( .A(n13986), .B(n13993), .Y(n13992) );
  NAND2X1 U12473 ( .A(n13985), .B(n764), .Y(n13993) );
  NAND2X1 U12474 ( .A(n13994), .B(n13995), .Y(n13986) );
  NAND2X1 U12475 ( .A(u_muldiv_dividend_q[16]), .B(n44827), .Y(n13995) );
  NAND2X1 U12476 ( .A(u_muldiv_quotient_q[16]), .B(n44822), .Y(n13994) );
  NAND2X1 U12477 ( .A(n13996), .B(n13997), .Y(u_muldiv_N536) );
  NOR2X1 U12479 ( .A(n13998), .B(n13999), .Y(n13996) );
  NOR2X1 U12480 ( .A(n764), .B(n709), .Y(n13999) );
  NOR2X1 U12481 ( .A(n14000), .B(n44629), .Y(n13998) );
  XNOR2X1 U12482 ( .A(n13985), .B(n764), .Y(n14000) );
  NAND2X1 U12483 ( .A(n14001), .B(n14002), .Y(n13987) );
  NAND2X1 U12484 ( .A(u_muldiv_dividend_q[15]), .B(n44827), .Y(n14002) );
  NAND2X1 U12485 ( .A(u_muldiv_quotient_q[15]), .B(n44822), .Y(n14001) );
  NOR2X1 U12486 ( .A(n14003), .B(n14004), .Y(n13985) );
  OR2X1 U12487 ( .A(n14005), .B(n14006), .Y(n14003) );
  NAND2X1 U12488 ( .A(n14007), .B(n14008), .Y(u_muldiv_N535) );
  NOR2X1 U12490 ( .A(n14009), .B(n14010), .Y(n14007) );
  NOR2X1 U12491 ( .A(n799), .B(n709), .Y(n14010) );
  NOR2X1 U12492 ( .A(n14011), .B(n44629), .Y(n14009) );
  XNOR2X1 U12493 ( .A(n799), .B(n14012), .Y(n14011) );
  NOR2X1 U12494 ( .A(n14006), .B(n14004), .Y(n14012) );
  NAND2X1 U12495 ( .A(n14013), .B(n14014), .Y(n14005) );
  NAND2X1 U12496 ( .A(u_muldiv_dividend_q[14]), .B(n44827), .Y(n14014) );
  NAND2X1 U12497 ( .A(u_muldiv_quotient_q[14]), .B(n44822), .Y(n14013) );
  NAND2X1 U12498 ( .A(n14015), .B(n14016), .Y(u_muldiv_N534) );
  NOR2X1 U12500 ( .A(n14017), .B(n14018), .Y(n14015) );
  AND2X1 U12501 ( .A(n14006), .B(n13846), .Y(n14018) );
  NOR2X1 U12502 ( .A(n14019), .B(n44628), .Y(n14017) );
  XNOR2X1 U12503 ( .A(n14004), .B(n14006), .Y(n14019) );
  NAND2X1 U12504 ( .A(n14020), .B(n14021), .Y(n14006) );
  NAND2X1 U12505 ( .A(u_muldiv_dividend_q[13]), .B(n44828), .Y(n14021) );
  NAND2X1 U12506 ( .A(u_muldiv_quotient_q[13]), .B(n44822), .Y(n14020) );
  NAND2X1 U12507 ( .A(n14022), .B(n14023), .Y(n14004) );
  NOR2X1 U12508 ( .A(n14024), .B(n14025), .Y(n14022) );
  NAND2X1 U12509 ( .A(n14026), .B(n14027), .Y(u_muldiv_N533) );
  NOR2X1 U12511 ( .A(n14028), .B(n14029), .Y(n14026) );
  AND2X1 U12512 ( .A(n14024), .B(n13846), .Y(n14029) );
  NOR2X1 U12513 ( .A(n14030), .B(n44628), .Y(n14028) );
  XNOR2X1 U12514 ( .A(n14024), .B(n14031), .Y(n14030) );
  NAND2X1 U12515 ( .A(n14023), .B(n871), .Y(n14031) );
  NAND2X1 U12516 ( .A(n14032), .B(n14033), .Y(n14024) );
  NAND2X1 U12517 ( .A(u_muldiv_dividend_q[12]), .B(n44828), .Y(n14033) );
  NAND2X1 U12518 ( .A(u_muldiv_quotient_q[12]), .B(n44822), .Y(n14032) );
  NAND2X1 U12519 ( .A(n14034), .B(n14035), .Y(u_muldiv_N532) );
  NOR2X1 U12521 ( .A(n14036), .B(n14037), .Y(n14034) );
  NOR2X1 U12522 ( .A(n871), .B(n709), .Y(n14037) );
  NOR2X1 U12523 ( .A(n14038), .B(n44628), .Y(n14036) );
  XNOR2X1 U12524 ( .A(n14023), .B(n871), .Y(n14038) );
  NAND2X1 U12525 ( .A(n14039), .B(n14040), .Y(n14025) );
  NAND2X1 U12526 ( .A(u_muldiv_dividend_q[11]), .B(n44828), .Y(n14040) );
  NAND2X1 U12527 ( .A(u_muldiv_quotient_q[11]), .B(n44822), .Y(n14039) );
  NOR2X1 U12528 ( .A(n14041), .B(n14042), .Y(n14023) );
  OR2X1 U12529 ( .A(n14043), .B(n14044), .Y(n14041) );
  NAND2X1 U12530 ( .A(n14045), .B(n14046), .Y(u_muldiv_N531) );
  NOR2X1 U12532 ( .A(n14047), .B(n14048), .Y(n14045) );
  NOR2X1 U12533 ( .A(n870), .B(n709), .Y(n14048) );
  NOR2X1 U12534 ( .A(n14049), .B(n44628), .Y(n14047) );
  XNOR2X1 U12535 ( .A(n870), .B(n14050), .Y(n14049) );
  NOR2X1 U12536 ( .A(n14044), .B(n14042), .Y(n14050) );
  NAND2X1 U12537 ( .A(n14051), .B(n14052), .Y(n14043) );
  NAND2X1 U12538 ( .A(u_muldiv_dividend_q[10]), .B(n44829), .Y(n14052) );
  NAND2X1 U12539 ( .A(u_muldiv_quotient_q[10]), .B(n44823), .Y(n14051) );
  NAND2X1 U12540 ( .A(n14053), .B(n14054), .Y(u_muldiv_N530) );
  NOR2X1 U12542 ( .A(n14055), .B(n14056), .Y(n14053) );
  AND2X1 U12543 ( .A(n14044), .B(n13846), .Y(n14056) );
  NOR2X1 U12544 ( .A(n14057), .B(n44628), .Y(n14055) );
  XNOR2X1 U12545 ( .A(n14042), .B(n14044), .Y(n14057) );
  NAND2X1 U12546 ( .A(n14058), .B(n14059), .Y(n14044) );
  NAND2X1 U12547 ( .A(u_muldiv_dividend_q[9]), .B(n44829), .Y(n14059) );
  NAND2X1 U12548 ( .A(u_muldiv_quotient_q[9]), .B(n44823), .Y(n14058) );
  NAND2X1 U12549 ( .A(n14060), .B(n14061), .Y(n14042) );
  NOR2X1 U12550 ( .A(n14062), .B(n14063), .Y(n14060) );
  NAND2X1 U12551 ( .A(n14064), .B(n14065), .Y(u_muldiv_N529) );
  NOR2X1 U12553 ( .A(n14066), .B(n14067), .Y(n14064) );
  AND2X1 U12554 ( .A(n14062), .B(n13846), .Y(n14067) );
  NOR2X1 U12555 ( .A(n14068), .B(n44628), .Y(n14066) );
  XNOR2X1 U12556 ( .A(n14062), .B(n14069), .Y(n14068) );
  NAND2X1 U12557 ( .A(n14061), .B(n869), .Y(n14069) );
  NAND2X1 U12558 ( .A(n14070), .B(n14071), .Y(n14062) );
  NAND2X1 U12559 ( .A(u_muldiv_dividend_q[8]), .B(n44829), .Y(n14071) );
  NAND2X1 U12560 ( .A(u_muldiv_quotient_q[8]), .B(n44820), .Y(n14070) );
  NAND2X1 U12561 ( .A(n14072), .B(n14073), .Y(u_muldiv_N528) );
  NOR2X1 U12563 ( .A(n14074), .B(n14075), .Y(n14072) );
  NOR2X1 U12564 ( .A(n869), .B(n709), .Y(n14075) );
  NOR2X1 U12565 ( .A(n14076), .B(n44628), .Y(n14074) );
  XNOR2X1 U12566 ( .A(n14061), .B(n869), .Y(n14076) );
  NAND2X1 U12567 ( .A(n14077), .B(n14078), .Y(n14063) );
  NAND2X1 U12568 ( .A(u_muldiv_dividend_q[7]), .B(n44830), .Y(n14078) );
  NAND2X1 U12569 ( .A(u_muldiv_quotient_q[7]), .B(n44820), .Y(n14077) );
  NOR2X1 U12570 ( .A(n14079), .B(n14080), .Y(n14061) );
  OR2X1 U12571 ( .A(n14081), .B(n14082), .Y(n14079) );
  NAND2X1 U12572 ( .A(n14083), .B(n14084), .Y(u_muldiv_N527) );
  NOR2X1 U12574 ( .A(n14085), .B(n14086), .Y(n14083) );
  NOR2X1 U12575 ( .A(n868), .B(n709), .Y(n14086) );
  NOR2X1 U12576 ( .A(n14087), .B(n44628), .Y(n14085) );
  XNOR2X1 U12577 ( .A(n868), .B(n14088), .Y(n14087) );
  NOR2X1 U12578 ( .A(n14082), .B(n14080), .Y(n14088) );
  NAND2X1 U12579 ( .A(n14089), .B(n14090), .Y(n14081) );
  NAND2X1 U12580 ( .A(u_muldiv_dividend_q[6]), .B(n44830), .Y(n14090) );
  NAND2X1 U12581 ( .A(u_muldiv_quotient_q[6]), .B(n44820), .Y(n14089) );
  NAND2X1 U12582 ( .A(n14091), .B(n14092), .Y(u_muldiv_N526) );
  NOR2X1 U12584 ( .A(n14093), .B(n14094), .Y(n14091) );
  AND2X1 U12585 ( .A(n14082), .B(n13846), .Y(n14094) );
  NOR2X1 U12586 ( .A(n14095), .B(n44628), .Y(n14093) );
  XNOR2X1 U12587 ( .A(n14080), .B(n14082), .Y(n14095) );
  NAND2X1 U12588 ( .A(n14096), .B(n14097), .Y(n14082) );
  NAND2X1 U12589 ( .A(u_muldiv_dividend_q[5]), .B(n44830), .Y(n14097) );
  NAND2X1 U12590 ( .A(u_muldiv_quotient_q[5]), .B(n44820), .Y(n14096) );
  NAND2X1 U12591 ( .A(n14098), .B(n14099), .Y(n14080) );
  NOR2X1 U12592 ( .A(n14100), .B(n14101), .Y(n14098) );
  NAND2X1 U12593 ( .A(n14102), .B(n14103), .Y(u_muldiv_N525) );
  NOR2X1 U12595 ( .A(n14104), .B(n14105), .Y(n14102) );
  AND2X1 U12596 ( .A(n14100), .B(n13846), .Y(n14105) );
  NOR2X1 U12597 ( .A(n14106), .B(n44628), .Y(n14104) );
  XNOR2X1 U12598 ( .A(n14100), .B(n14107), .Y(n14106) );
  NAND2X1 U12599 ( .A(n14099), .B(n833), .Y(n14107) );
  NAND2X1 U12600 ( .A(n14108), .B(n14109), .Y(n14100) );
  NAND2X1 U12601 ( .A(u_muldiv_dividend_q[4]), .B(n44821), .Y(n14109) );
  NAND2X1 U12602 ( .A(u_muldiv_quotient_q[4]), .B(u_muldiv_div_inst_q), .Y(
        n14108) );
  NAND2X1 U12603 ( .A(n14110), .B(n14111), .Y(u_muldiv_N524) );
  NOR2X1 U12605 ( .A(n14112), .B(n14113), .Y(n14110) );
  NOR2X1 U12606 ( .A(n833), .B(n709), .Y(n14113) );
  NOR2X1 U12607 ( .A(n14114), .B(n44628), .Y(n14112) );
  XNOR2X1 U12608 ( .A(n14099), .B(n833), .Y(n14114) );
  NAND2X1 U12609 ( .A(n14115), .B(n14116), .Y(n14101) );
  NAND2X1 U12610 ( .A(u_muldiv_dividend_q[3]), .B(n44821), .Y(n14116) );
  NAND2X1 U12611 ( .A(u_muldiv_quotient_q[3]), .B(u_muldiv_div_inst_q), .Y(
        n14115) );
  AND2X1 U12612 ( .A(n14117), .B(n712), .Y(n14099) );
  NOR2X1 U12613 ( .A(n14118), .B(n14119), .Y(n14117) );
  NAND2X1 U12614 ( .A(n14120), .B(n14121), .Y(u_muldiv_N523) );
  NOR2X1 U12615 ( .A(n14122), .B(n14123), .Y(n14121) );
  NOR2X1 U12616 ( .A(n14118), .B(n710), .Y(n14123) );
  NOR2X1 U12617 ( .A(n14124), .B(n44628), .Y(n14122) );
  NOR2X1 U12618 ( .A(n14125), .B(n14126), .Y(n14124) );
  NOR2X1 U12619 ( .A(n817), .B(n14118), .Y(n14126) );
  NOR2X1 U12620 ( .A(n14127), .B(n14128), .Y(n14125) );
  NAND2X1 U12621 ( .A(n817), .B(n14118), .Y(n14128) );
  NOR2X1 U12622 ( .A(n14129), .B(n14130), .Y(n14120) );
  AND2X1 U12624 ( .A(n14118), .B(n13846), .Y(n14129) );
  NAND2X1 U12625 ( .A(n14131), .B(n14132), .Y(n14118) );
  NAND2X1 U12626 ( .A(u_muldiv_dividend_q[2]), .B(n37586), .Y(n14132) );
  NAND2X1 U12627 ( .A(u_muldiv_quotient_q[2]), .B(u_muldiv_div_inst_q), .Y(
        n14131) );
  NAND2X1 U12628 ( .A(n14133), .B(n14134), .Y(u_muldiv_N522) );
  NOR2X1 U12630 ( .A(n14135), .B(n14136), .Y(n14133) );
  NOR2X1 U12631 ( .A(n14119), .B(n710), .Y(n14136) );
  NOR2X1 U12632 ( .A(n817), .B(n14138), .Y(n14135) );
  NOR2X1 U12633 ( .A(n14139), .B(n13846), .Y(n14138) );
  NOR2X1 U12634 ( .A(n14127), .B(n44628), .Y(n14139) );
  NAND2X1 U12635 ( .A(n14140), .B(n14141), .Y(n14119) );
  NAND2X1 U12636 ( .A(u_muldiv_dividend_q[1]), .B(n37586), .Y(n14141) );
  NAND2X1 U12637 ( .A(u_muldiv_quotient_q[1]), .B(u_muldiv_div_inst_q), .Y(
        n14140) );
  NAND2X1 U12638 ( .A(n14142), .B(n14143), .Y(u_muldiv_N521) );
  NAND2X1 U12639 ( .A(u_muldiv_mult_result_q[0]), .B(n44632), .Y(n14143) );
  NOR2X1 U12640 ( .A(n14137), .B(n14144), .Y(n14142) );
  NOR2X1 U12641 ( .A(n712), .B(n709), .Y(n14144) );
  NOR2X1 U12642 ( .A(n44631), .B(u_muldiv_invert_res_q), .Y(n13846) );
  NOR2X1 U12643 ( .A(n44628), .B(n712), .Y(n14137) );
  NAND2X1 U12644 ( .A(n14145), .B(n14146), .Y(n14127) );
  NAND2X1 U12645 ( .A(u_muldiv_dividend_q[0]), .B(n37586), .Y(n14146) );
  NAND2X1 U12646 ( .A(u_muldiv_quotient_q[0]), .B(u_muldiv_div_inst_q), .Y(
        n14145) );
  NOR2X1 U12648 ( .A(n14147), .B(n37781), .Y(u_muldiv_N517) );
  NOR2X1 U12649 ( .A(n14147), .B(n37780), .Y(u_muldiv_N516) );
  NOR2X1 U12650 ( .A(n14147), .B(n37779), .Y(u_muldiv_N515) );
  NOR2X1 U12651 ( .A(n14147), .B(n37778), .Y(u_muldiv_N514) );
  NOR2X1 U12652 ( .A(n14147), .B(n37777), .Y(u_muldiv_N513) );
  NOR2X1 U12653 ( .A(u_muldiv_mult_busy_q), .B(n37333), .Y(n14147) );
  NOR2X1 U12654 ( .A(n14165), .B(n44625), .Y(u_muldiv_N359) );
  NOR2X1 U12655 ( .A(u_muldiv_q_mask_q[31]), .B(u_muldiv_quotient_q[31]), .Y(
        n14165) );
  NOR2X1 U12656 ( .A(n14167), .B(n44626), .Y(u_muldiv_N358) );
  NOR2X1 U12657 ( .A(u_muldiv_q_mask_q[30]), .B(u_muldiv_quotient_q[30]), .Y(
        n14167) );
  NOR2X1 U12658 ( .A(n14168), .B(n44625), .Y(u_muldiv_N357) );
  NOR2X1 U12659 ( .A(u_muldiv_q_mask_q[29]), .B(u_muldiv_quotient_q[29]), .Y(
        n14168) );
  NOR2X1 U12660 ( .A(n14169), .B(n44626), .Y(u_muldiv_N356) );
  NOR2X1 U12661 ( .A(u_muldiv_q_mask_q[28]), .B(u_muldiv_quotient_q[28]), .Y(
        n14169) );
  NOR2X1 U12662 ( .A(n14170), .B(n44626), .Y(u_muldiv_N355) );
  NOR2X1 U12663 ( .A(u_muldiv_q_mask_q[27]), .B(u_muldiv_quotient_q[27]), .Y(
        n14170) );
  NOR2X1 U12664 ( .A(n14171), .B(n44626), .Y(u_muldiv_N354) );
  NOR2X1 U12665 ( .A(u_muldiv_q_mask_q[26]), .B(u_muldiv_quotient_q[26]), .Y(
        n14171) );
  NOR2X1 U12666 ( .A(n14172), .B(n44625), .Y(u_muldiv_N353) );
  NOR2X1 U12667 ( .A(u_muldiv_q_mask_q[25]), .B(u_muldiv_quotient_q[25]), .Y(
        n14172) );
  NOR2X1 U12668 ( .A(n14173), .B(n44625), .Y(u_muldiv_N352) );
  NOR2X1 U12669 ( .A(u_muldiv_q_mask_q[24]), .B(u_muldiv_quotient_q[24]), .Y(
        n14173) );
  NOR2X1 U12670 ( .A(n14174), .B(n44625), .Y(u_muldiv_N351) );
  NOR2X1 U12671 ( .A(u_muldiv_q_mask_q[23]), .B(u_muldiv_quotient_q[23]), .Y(
        n14174) );
  NOR2X1 U12672 ( .A(n14175), .B(n44625), .Y(u_muldiv_N350) );
  NOR2X1 U12673 ( .A(u_muldiv_q_mask_q[22]), .B(u_muldiv_quotient_q[22]), .Y(
        n14175) );
  NOR2X1 U12674 ( .A(n14176), .B(n44625), .Y(u_muldiv_N349) );
  NOR2X1 U12675 ( .A(u_muldiv_q_mask_q[21]), .B(u_muldiv_quotient_q[21]), .Y(
        n14176) );
  NOR2X1 U12676 ( .A(n14177), .B(n44626), .Y(u_muldiv_N348) );
  NOR2X1 U12677 ( .A(u_muldiv_q_mask_q[20]), .B(u_muldiv_quotient_q[20]), .Y(
        n14177) );
  NOR2X1 U12678 ( .A(n14178), .B(n44625), .Y(u_muldiv_N347) );
  NOR2X1 U12679 ( .A(u_muldiv_q_mask_q[19]), .B(u_muldiv_quotient_q[19]), .Y(
        n14178) );
  NOR2X1 U12680 ( .A(n14179), .B(n44623), .Y(u_muldiv_N346) );
  NOR2X1 U12681 ( .A(u_muldiv_q_mask_q[18]), .B(u_muldiv_quotient_q[18]), .Y(
        n14179) );
  NAND2X1 U12682 ( .A(n14148), .B(n14180), .Y(u_muldiv_N345) );
  NAND2X1 U12683 ( .A(n44610), .B(u_muldiv_quotient_q[17]), .Y(n14180) );
  NAND2X1 U12684 ( .A(u_muldiv_q_mask_q[17]), .B(n44615), .Y(n14148) );
  NAND2X1 U12685 ( .A(n14149), .B(n14181), .Y(u_muldiv_N344) );
  NAND2X1 U12686 ( .A(n44612), .B(u_muldiv_quotient_q[16]), .Y(n14181) );
  NAND2X1 U12687 ( .A(u_muldiv_q_mask_q[16]), .B(n44616), .Y(n14149) );
  NAND2X1 U12688 ( .A(n14150), .B(n14182), .Y(u_muldiv_N343) );
  NAND2X1 U12689 ( .A(n44614), .B(u_muldiv_quotient_q[15]), .Y(n14182) );
  NAND2X1 U12690 ( .A(u_muldiv_q_mask_q[15]), .B(n44615), .Y(n14150) );
  NAND2X1 U12691 ( .A(n14151), .B(n14183), .Y(u_muldiv_N342) );
  NAND2X1 U12692 ( .A(n44614), .B(u_muldiv_quotient_q[14]), .Y(n14183) );
  NAND2X1 U12693 ( .A(u_muldiv_q_mask_q[14]), .B(n44615), .Y(n14151) );
  NAND2X1 U12694 ( .A(n14152), .B(n14184), .Y(u_muldiv_N341) );
  NAND2X1 U12695 ( .A(n44613), .B(u_muldiv_quotient_q[13]), .Y(n14184) );
  NAND2X1 U12696 ( .A(u_muldiv_q_mask_q[13]), .B(n44615), .Y(n14152) );
  NAND2X1 U12697 ( .A(n14153), .B(n14185), .Y(u_muldiv_N340) );
  NAND2X1 U12698 ( .A(n44613), .B(u_muldiv_quotient_q[12]), .Y(n14185) );
  NAND2X1 U12699 ( .A(u_muldiv_q_mask_q[12]), .B(n44615), .Y(n14153) );
  NAND2X1 U12700 ( .A(n14154), .B(n14186), .Y(u_muldiv_N339) );
  NAND2X1 U12701 ( .A(n44613), .B(u_muldiv_quotient_q[11]), .Y(n14186) );
  NAND2X1 U12702 ( .A(u_muldiv_q_mask_q[11]), .B(n44615), .Y(n14154) );
  NAND2X1 U12703 ( .A(n14155), .B(n14187), .Y(u_muldiv_N338) );
  NAND2X1 U12704 ( .A(n44613), .B(u_muldiv_quotient_q[10]), .Y(n14187) );
  NAND2X1 U12705 ( .A(u_muldiv_q_mask_q[10]), .B(n44615), .Y(n14155) );
  NAND2X1 U12706 ( .A(n14156), .B(n14188), .Y(u_muldiv_N337) );
  NAND2X1 U12707 ( .A(n44613), .B(u_muldiv_quotient_q[9]), .Y(n14188) );
  NAND2X1 U12708 ( .A(u_muldiv_q_mask_q[9]), .B(n44616), .Y(n14156) );
  NAND2X1 U12709 ( .A(n14157), .B(n14189), .Y(u_muldiv_N336) );
  NAND2X1 U12710 ( .A(n44613), .B(u_muldiv_quotient_q[8]), .Y(n14189) );
  NAND2X1 U12711 ( .A(u_muldiv_q_mask_q[8]), .B(n44615), .Y(n14157) );
  NAND2X1 U12712 ( .A(n14158), .B(n14190), .Y(u_muldiv_N335) );
  NAND2X1 U12713 ( .A(n44613), .B(u_muldiv_quotient_q[7]), .Y(n14190) );
  NAND2X1 U12714 ( .A(u_muldiv_q_mask_q[7]), .B(n44615), .Y(n14158) );
  NAND2X1 U12715 ( .A(n14159), .B(n14191), .Y(u_muldiv_N334) );
  NAND2X1 U12716 ( .A(n44612), .B(u_muldiv_quotient_q[6]), .Y(n14191) );
  NAND2X1 U12717 ( .A(u_muldiv_q_mask_q[6]), .B(n44617), .Y(n14159) );
  NAND2X1 U12718 ( .A(n14160), .B(n14192), .Y(u_muldiv_N333) );
  NAND2X1 U12719 ( .A(n44613), .B(u_muldiv_quotient_q[5]), .Y(n14192) );
  NAND2X1 U12720 ( .A(u_muldiv_q_mask_q[5]), .B(n44617), .Y(n14160) );
  NAND2X1 U12721 ( .A(n14161), .B(n14193), .Y(u_muldiv_N332) );
  NAND2X1 U12722 ( .A(n44613), .B(u_muldiv_quotient_q[4]), .Y(n14193) );
  NAND2X1 U12723 ( .A(u_muldiv_q_mask_q[4]), .B(n44617), .Y(n14161) );
  NAND2X1 U12724 ( .A(n14162), .B(n14194), .Y(u_muldiv_N331) );
  NAND2X1 U12725 ( .A(n44613), .B(u_muldiv_quotient_q[3]), .Y(n14194) );
  NAND2X1 U12726 ( .A(u_muldiv_q_mask_q[3]), .B(n44617), .Y(n14162) );
  NAND2X1 U12727 ( .A(n14163), .B(n14195), .Y(u_muldiv_N330) );
  NAND2X1 U12728 ( .A(n44613), .B(u_muldiv_quotient_q[2]), .Y(n14195) );
  NAND2X1 U12729 ( .A(u_muldiv_q_mask_q[2]), .B(n44616), .Y(n14163) );
  NAND2X1 U12730 ( .A(n14164), .B(n14196), .Y(u_muldiv_N329) );
  NAND2X1 U12731 ( .A(n44613), .B(u_muldiv_quotient_q[1]), .Y(n14196) );
  NAND2X1 U12732 ( .A(u_muldiv_q_mask_q[1]), .B(n44616), .Y(n14164) );
  NOR2X1 U12733 ( .A(n14197), .B(n44626), .Y(u_muldiv_N328) );
  NOR2X1 U12734 ( .A(u_muldiv_q_mask_q[0]), .B(u_muldiv_quotient_q[0]), .Y(
        n14197) );
  NAND2X1 U12738 ( .A(n14202), .B(n14203), .Y(u_muldiv_N326) );
  NAND2X1 U12739 ( .A(u_muldiv_divisor_q[62]), .B(n44618), .Y(n14203) );
  NAND2X1 U12746 ( .A(n14210), .B(n14211), .Y(u_muldiv_N325) );
  NAND2X1 U12747 ( .A(u_muldiv_divisor_q[61]), .B(n44618), .Y(n14211) );
  NAND2X1 U12754 ( .A(n14218), .B(n14219), .Y(u_muldiv_N324) );
  NAND2X1 U12755 ( .A(u_muldiv_divisor_q[60]), .B(n44618), .Y(n14219) );
  NAND2X1 U12763 ( .A(n14227), .B(n14228), .Y(u_muldiv_N323) );
  NAND2X1 U12764 ( .A(u_muldiv_divisor_q[59]), .B(n44616), .Y(n14228) );
  NAND2X1 U12771 ( .A(n14234), .B(n14235), .Y(u_muldiv_N322) );
  NAND2X1 U12772 ( .A(u_muldiv_divisor_q[58]), .B(n44618), .Y(n14235) );
  NAND2X1 U12780 ( .A(n14243), .B(n14244), .Y(u_muldiv_N321) );
  NAND2X1 U12781 ( .A(u_muldiv_divisor_q[57]), .B(n44618), .Y(n14244) );
  NAND2X1 U12788 ( .A(n14250), .B(n14251), .Y(u_muldiv_N320) );
  NAND2X1 U12789 ( .A(u_muldiv_divisor_q[56]), .B(n44614), .Y(n14251) );
  NAND2X1 U12796 ( .A(n14258), .B(n14259), .Y(u_muldiv_N319) );
  NAND2X1 U12797 ( .A(u_muldiv_divisor_q[55]), .B(n44618), .Y(n14259) );
  NAND2X1 U12804 ( .A(n14266), .B(n14267), .Y(u_muldiv_N318) );
  NAND2X1 U12805 ( .A(u_muldiv_divisor_q[54]), .B(n44617), .Y(n14267) );
  NAND2X1 U12813 ( .A(n14275), .B(n14276), .Y(u_muldiv_N317) );
  NAND2X1 U12814 ( .A(u_muldiv_divisor_q[53]), .B(n44618), .Y(n14276) );
  NAND2X1 U12821 ( .A(n14282), .B(n14283), .Y(u_muldiv_N316) );
  NAND2X1 U12822 ( .A(u_muldiv_divisor_q[52]), .B(n44618), .Y(n14283) );
  NAND2X1 U12830 ( .A(n14291), .B(n14292), .Y(u_muldiv_N315) );
  NAND2X1 U12831 ( .A(u_muldiv_divisor_q[51]), .B(n44617), .Y(n14292) );
  NAND2X1 U12838 ( .A(n14298), .B(n14299), .Y(u_muldiv_N314) );
  NAND2X1 U12839 ( .A(u_muldiv_divisor_q[50]), .B(n44617), .Y(n14299) );
  NAND2X1 U12847 ( .A(n14307), .B(n14308), .Y(u_muldiv_N313) );
  NAND2X1 U12848 ( .A(u_muldiv_divisor_q[49]), .B(n44617), .Y(n14308) );
  NAND2X1 U12855 ( .A(n14314), .B(n14315), .Y(u_muldiv_N312) );
  NAND2X1 U12856 ( .A(u_muldiv_divisor_q[48]), .B(n44617), .Y(n14315) );
  NAND2X1 U12864 ( .A(n14323), .B(n14324), .Y(u_muldiv_N311) );
  NAND2X1 U12865 ( .A(u_muldiv_divisor_q[47]), .B(n44617), .Y(n14324) );
  NAND2X1 U12872 ( .A(n14330), .B(n14331), .Y(u_muldiv_N310) );
  NAND2X1 U12873 ( .A(u_muldiv_divisor_q[46]), .B(n44617), .Y(n14331) );
  NAND2X1 U12881 ( .A(n14339), .B(n14340), .Y(u_muldiv_N309) );
  NAND2X1 U12882 ( .A(u_muldiv_divisor_q[45]), .B(n44617), .Y(n14340) );
  NAND2X1 U12889 ( .A(n14346), .B(n14347), .Y(u_muldiv_N308) );
  NAND2X1 U12890 ( .A(u_muldiv_divisor_q[44]), .B(n44615), .Y(n14347) );
  NAND2X1 U12898 ( .A(n14355), .B(n14356), .Y(u_muldiv_N307) );
  NAND2X1 U12899 ( .A(u_muldiv_divisor_q[43]), .B(n44617), .Y(n14356) );
  NAND2X1 U12906 ( .A(n14362), .B(n14363), .Y(u_muldiv_N306) );
  NAND2X1 U12907 ( .A(u_muldiv_divisor_q[42]), .B(n44616), .Y(n14363) );
  NAND2X1 U12915 ( .A(n14371), .B(n14372), .Y(u_muldiv_N305) );
  NAND2X1 U12916 ( .A(u_muldiv_divisor_q[41]), .B(n44618), .Y(n14372) );
  NAND2X1 U12923 ( .A(n14378), .B(n14379), .Y(u_muldiv_N304) );
  NAND2X1 U12924 ( .A(u_muldiv_divisor_q[40]), .B(n44618), .Y(n14379) );
  NAND2X1 U12932 ( .A(n14387), .B(n14388), .Y(u_muldiv_N303) );
  NAND2X1 U12933 ( .A(u_muldiv_divisor_q[39]), .B(n44618), .Y(n14388) );
  NAND2X1 U12940 ( .A(n14394), .B(n14395), .Y(u_muldiv_N302) );
  NAND2X1 U12941 ( .A(u_muldiv_divisor_q[38]), .B(n44618), .Y(n14395) );
  NAND2X1 U12949 ( .A(n14403), .B(n14404), .Y(u_muldiv_N301) );
  NAND2X1 U12950 ( .A(u_muldiv_divisor_q[37]), .B(n44618), .Y(n14404) );
  NAND2X1 U12957 ( .A(n14410), .B(n14411), .Y(u_muldiv_N300) );
  NAND2X1 U12958 ( .A(u_muldiv_divisor_q[36]), .B(n44616), .Y(n14411) );
  NAND2X1 U12966 ( .A(n14419), .B(n14420), .Y(u_muldiv_N299) );
  NAND2X1 U12967 ( .A(u_muldiv_divisor_q[35]), .B(n44616), .Y(n14420) );
  NAND2X1 U12974 ( .A(n14426), .B(n14427), .Y(u_muldiv_N298) );
  NAND2X1 U12975 ( .A(u_muldiv_divisor_q[34]), .B(n44616), .Y(n14427) );
  NAND2X1 U12984 ( .A(n14436), .B(n14437), .Y(u_muldiv_N297) );
  NAND2X1 U12985 ( .A(u_muldiv_divisor_q[33]), .B(n44616), .Y(n14437) );
  NAND2X1 U12991 ( .A(n14443), .B(n14444), .Y(u_muldiv_N296) );
  NAND2X1 U12992 ( .A(u_muldiv_divisor_q[32]), .B(n44616), .Y(n14444) );
  AND2X1 U13000 ( .A(n44627), .B(u_muldiv_divisor_q[31]), .Y(u_muldiv_N295) );
  NOR2X1 U13001 ( .A(n44619), .B(n37582), .Y(u_muldiv_N294) );
  NOR2X1 U13002 ( .A(n44619), .B(n37583), .Y(u_muldiv_N293) );
  NOR2X1 U13003 ( .A(n44622), .B(n37576), .Y(u_muldiv_N292) );
  NOR2X1 U13004 ( .A(n44623), .B(n37573), .Y(u_muldiv_N291) );
  NOR2X1 U13005 ( .A(n44621), .B(n42553), .Y(u_muldiv_N290) );
  NOR2X1 U13006 ( .A(n44626), .B(n37564), .Y(u_muldiv_N289) );
  NOR2X1 U13007 ( .A(n44623), .B(n37559), .Y(u_muldiv_N288) );
  NOR2X1 U13008 ( .A(n44620), .B(n37557), .Y(u_muldiv_N287) );
  NOR2X1 U13009 ( .A(n44622), .B(n42551), .Y(u_muldiv_N286) );
  NOR2X1 U13010 ( .A(n44621), .B(n37551), .Y(u_muldiv_N285) );
  NOR2X1 U13011 ( .A(n44622), .B(n37543), .Y(u_muldiv_N284) );
  NOR2X1 U13012 ( .A(n44621), .B(n37538), .Y(u_muldiv_N283) );
  NOR2X1 U13013 ( .A(n44620), .B(n42549), .Y(u_muldiv_N282) );
  NOR2X1 U13014 ( .A(n44620), .B(n37453), .Y(u_muldiv_N281) );
  NOR2X1 U13015 ( .A(n44620), .B(n37452), .Y(u_muldiv_N280) );
  NOR2X1 U13016 ( .A(n44620), .B(n37447), .Y(u_muldiv_N279) );
  NOR2X1 U13017 ( .A(n44620), .B(n42547), .Y(u_muldiv_N278) );
  NOR2X1 U13018 ( .A(n44621), .B(n37443), .Y(u_muldiv_N277) );
  NOR2X1 U13019 ( .A(n44621), .B(n37442), .Y(u_muldiv_N276) );
  NOR2X1 U13020 ( .A(n44621), .B(n37440), .Y(u_muldiv_N275) );
  NOR2X1 U13021 ( .A(n44622), .B(n42555), .Y(u_muldiv_N274) );
  NOR2X1 U13022 ( .A(n44621), .B(n37432), .Y(u_muldiv_N273) );
  NOR2X1 U13023 ( .A(n44622), .B(n37429), .Y(u_muldiv_N272) );
  NOR2X1 U13024 ( .A(n44623), .B(n37427), .Y(u_muldiv_N271) );
  NOR2X1 U13025 ( .A(n44622), .B(n37424), .Y(u_muldiv_N270) );
  NOR2X1 U13026 ( .A(n44622), .B(n37422), .Y(u_muldiv_N269) );
  NOR2X1 U13027 ( .A(n44623), .B(n37421), .Y(u_muldiv_N268) );
  NOR2X1 U13028 ( .A(n44623), .B(n37438), .Y(u_muldiv_N267) );
  NOR2X1 U13029 ( .A(n44624), .B(n37435), .Y(u_muldiv_N266) );
  NOR2X1 U13030 ( .A(n44623), .B(n37419), .Y(u_muldiv_N265) );
  NAND2X1 U13036 ( .A(n44612), .B(n14457), .Y(n14449) );
  XNOR2X1 U13037 ( .A(n14458), .B(n14459), .Y(n14457) );
  NOR2X1 U13038 ( .A(n14460), .B(n708), .Y(n14459) );
  NOR2X1 U13039 ( .A(n713), .B(n14461), .Y(n14460) );
  XNOR2X1 U13040 ( .A(u_muldiv_divisor_q[31]), .B(u_muldiv_dividend_q[31]), 
        .Y(n14458) );
  NAND2X1 U13041 ( .A(n14462), .B(n14463), .Y(u_muldiv_N262) );
  NAND2X1 U13042 ( .A(n44612), .B(n14464), .Y(n14463) );
  NAND2X1 U13043 ( .A(n14465), .B(n14466), .Y(n14464) );
  NAND2X1 U13044 ( .A(n14467), .B(n713), .Y(n14466) );
  XNOR2X1 U13045 ( .A(u_muldiv_divisor_q[30]), .B(u_muldiv_dividend_q[30]), 
        .Y(n14467) );
  NAND2X1 U13046 ( .A(n14469), .B(n14468), .Y(n14465) );
  NAND2X1 U13047 ( .A(n14470), .B(n14471), .Y(n14468) );
  NAND2X1 U13048 ( .A(n14472), .B(n37583), .Y(n14471) );
  NAND2X1 U13049 ( .A(n714), .B(n1630), .Y(n14472) );
  NAND2X1 U13050 ( .A(u_muldiv_dividend_q[29]), .B(n14473), .Y(n14470) );
  OR2X1 U13051 ( .A(n14461), .B(n708), .Y(n14469) );
  NAND2X1 U13059 ( .A(n14481), .B(n14482), .Y(u_muldiv_N261) );
  NAND2X1 U13060 ( .A(n44612), .B(n14483), .Y(n14482) );
  XNOR2X1 U13061 ( .A(n14484), .B(n714), .Y(n14483) );
  NAND2X1 U13062 ( .A(n14485), .B(n14486), .Y(n14473) );
  NAND2X1 U13063 ( .A(n14487), .B(n37576), .Y(n14486) );
  NAND2X1 U13064 ( .A(n715), .B(n805), .Y(n14487) );
  NAND2X1 U13065 ( .A(u_muldiv_dividend_q[28]), .B(n14488), .Y(n14485) );
  XNOR2X1 U13066 ( .A(u_muldiv_divisor_q[29]), .B(u_muldiv_dividend_q[29]), 
        .Y(n14484) );
  NAND2X1 U13074 ( .A(n14495), .B(n14496), .Y(u_muldiv_N260) );
  NAND2X1 U13075 ( .A(n44612), .B(n14497), .Y(n14496) );
  XNOR2X1 U13076 ( .A(n14498), .B(n715), .Y(n14497) );
  NAND2X1 U13077 ( .A(n14499), .B(n14500), .Y(n14488) );
  NAND2X1 U13078 ( .A(n14501), .B(n37573), .Y(n14500) );
  NAND2X1 U13079 ( .A(n716), .B(n1561), .Y(n14501) );
  NAND2X1 U13080 ( .A(u_muldiv_dividend_q[27]), .B(n14502), .Y(n14499) );
  XNOR2X1 U13081 ( .A(u_muldiv_divisor_q[28]), .B(u_muldiv_dividend_q[28]), 
        .Y(n14498) );
  NAND2X1 U13089 ( .A(n14509), .B(n14510), .Y(u_muldiv_N259) );
  NAND2X1 U13090 ( .A(n44612), .B(n14511), .Y(n14510) );
  XNOR2X1 U13091 ( .A(n14512), .B(n716), .Y(n14511) );
  NAND2X1 U13092 ( .A(n14513), .B(n14514), .Y(n14502) );
  NAND2X1 U13093 ( .A(n14515), .B(n42553), .Y(n14514) );
  NAND2X1 U13094 ( .A(n717), .B(n1511), .Y(n14515) );
  NAND2X1 U13095 ( .A(u_muldiv_dividend_q[26]), .B(n14516), .Y(n14513) );
  XNOR2X1 U13096 ( .A(u_muldiv_divisor_q[27]), .B(u_muldiv_dividend_q[27]), 
        .Y(n14512) );
  NAND2X1 U13104 ( .A(n14523), .B(n14524), .Y(u_muldiv_N258) );
  NAND2X1 U13105 ( .A(n44612), .B(n14525), .Y(n14524) );
  XNOR2X1 U13106 ( .A(n14526), .B(n717), .Y(n14525) );
  NAND2X1 U13107 ( .A(n14527), .B(n14528), .Y(n14516) );
  NAND2X1 U13108 ( .A(n14529), .B(n37564), .Y(n14528) );
  OR2X1 U13109 ( .A(n14530), .B(u_muldiv_dividend_q[25]), .Y(n14529) );
  NAND2X1 U13110 ( .A(u_muldiv_dividend_q[25]), .B(n14530), .Y(n14527) );
  XNOR2X1 U13111 ( .A(u_muldiv_divisor_q[26]), .B(u_muldiv_dividend_q[26]), 
        .Y(n14526) );
  NAND2X1 U13119 ( .A(n14537), .B(n14538), .Y(u_muldiv_N257) );
  NAND2X1 U13120 ( .A(n44612), .B(n14539), .Y(n14538) );
  XOR2X1 U13121 ( .A(n14540), .B(n14530), .Y(n14539) );
  NAND2X1 U13122 ( .A(n14541), .B(n14542), .Y(n14530) );
  NAND2X1 U13123 ( .A(n14543), .B(n37559), .Y(n14542) );
  NAND2X1 U13124 ( .A(n718), .B(n1582), .Y(n14543) );
  NAND2X1 U13125 ( .A(u_muldiv_dividend_q[24]), .B(n14544), .Y(n14541) );
  XNOR2X1 U13126 ( .A(u_muldiv_divisor_q[25]), .B(u_muldiv_dividend_q[25]), 
        .Y(n14540) );
  NAND2X1 U13134 ( .A(n14551), .B(n14552), .Y(u_muldiv_N256) );
  NAND2X1 U13135 ( .A(n44612), .B(n14553), .Y(n14552) );
  XNOR2X1 U13136 ( .A(n14554), .B(n718), .Y(n14553) );
  NAND2X1 U13137 ( .A(n14555), .B(n14556), .Y(n14544) );
  NAND2X1 U13138 ( .A(n14557), .B(n37557), .Y(n14556) );
  NAND2X1 U13139 ( .A(n719), .B(n1459), .Y(n14557) );
  NAND2X1 U13140 ( .A(u_muldiv_dividend_q[23]), .B(n14558), .Y(n14555) );
  XNOR2X1 U13141 ( .A(u_muldiv_divisor_q[24]), .B(u_muldiv_dividend_q[24]), 
        .Y(n14554) );
  NAND2X1 U13149 ( .A(n14565), .B(n14566), .Y(u_muldiv_N255) );
  NAND2X1 U13150 ( .A(n44612), .B(n14567), .Y(n14566) );
  XNOR2X1 U13151 ( .A(n14568), .B(n719), .Y(n14567) );
  NAND2X1 U13152 ( .A(n14569), .B(n14570), .Y(n14558) );
  NAND2X1 U13153 ( .A(n14571), .B(n42551), .Y(n14570) );
  NAND2X1 U13154 ( .A(n720), .B(n1471), .Y(n14571) );
  NAND2X1 U13155 ( .A(u_muldiv_dividend_q[22]), .B(n14572), .Y(n14569) );
  XNOR2X1 U13156 ( .A(u_muldiv_divisor_q[23]), .B(u_muldiv_dividend_q[23]), 
        .Y(n14568) );
  NAND2X1 U13164 ( .A(n14579), .B(n14580), .Y(u_muldiv_N254) );
  NAND2X1 U13165 ( .A(n44611), .B(n14581), .Y(n14580) );
  XNOR2X1 U13166 ( .A(n14582), .B(n720), .Y(n14581) );
  NAND2X1 U13167 ( .A(n14583), .B(n14584), .Y(n14572) );
  NAND2X1 U13168 ( .A(n14585), .B(n37551), .Y(n14584) );
  OR2X1 U13169 ( .A(n14586), .B(u_muldiv_dividend_q[21]), .Y(n14585) );
  NAND2X1 U13170 ( .A(u_muldiv_dividend_q[21]), .B(n14586), .Y(n14583) );
  XNOR2X1 U13171 ( .A(u_muldiv_divisor_q[22]), .B(u_muldiv_dividend_q[22]), 
        .Y(n14582) );
  NAND2X1 U13179 ( .A(n14593), .B(n14594), .Y(u_muldiv_N253) );
  NAND2X1 U13180 ( .A(n44611), .B(n14595), .Y(n14594) );
  XOR2X1 U13181 ( .A(n14596), .B(n14586), .Y(n14595) );
  NAND2X1 U13182 ( .A(n14597), .B(n14598), .Y(n14586) );
  NAND2X1 U13183 ( .A(n14599), .B(n37543), .Y(n14598) );
  NAND2X1 U13184 ( .A(n721), .B(n1439), .Y(n14599) );
  NAND2X1 U13185 ( .A(u_muldiv_dividend_q[20]), .B(n14600), .Y(n14597) );
  XNOR2X1 U13186 ( .A(u_muldiv_divisor_q[21]), .B(u_muldiv_dividend_q[21]), 
        .Y(n14596) );
  NAND2X1 U13194 ( .A(n14607), .B(n14608), .Y(u_muldiv_N252) );
  NAND2X1 U13195 ( .A(n44611), .B(n14609), .Y(n14608) );
  XNOR2X1 U13196 ( .A(n14610), .B(n721), .Y(n14609) );
  NAND2X1 U13197 ( .A(n14611), .B(n14612), .Y(n14600) );
  NAND2X1 U13198 ( .A(n14613), .B(n37538), .Y(n14612) );
  NAND2X1 U13199 ( .A(n722), .B(n1409), .Y(n14613) );
  NAND2X1 U13200 ( .A(u_muldiv_dividend_q[19]), .B(n14614), .Y(n14611) );
  XNOR2X1 U13201 ( .A(u_muldiv_divisor_q[20]), .B(u_muldiv_dividend_q[20]), 
        .Y(n14610) );
  NAND2X1 U13209 ( .A(n14621), .B(n14622), .Y(u_muldiv_N251) );
  NAND2X1 U13210 ( .A(n44611), .B(n14623), .Y(n14622) );
  XNOR2X1 U13211 ( .A(n14624), .B(n722), .Y(n14623) );
  NAND2X1 U13212 ( .A(n14625), .B(n14626), .Y(n14614) );
  NAND2X1 U13213 ( .A(n14627), .B(n42549), .Y(n14626) );
  NAND2X1 U13214 ( .A(n723), .B(n37461), .Y(n14627) );
  NAND2X1 U13215 ( .A(u_muldiv_dividend_q[18]), .B(n14628), .Y(n14625) );
  XNOR2X1 U13216 ( .A(u_muldiv_divisor_q[19]), .B(u_muldiv_dividend_q[19]), 
        .Y(n14624) );
  NAND2X1 U13224 ( .A(n14635), .B(n14636), .Y(u_muldiv_N250) );
  NAND2X1 U13225 ( .A(n44611), .B(n14637), .Y(n14636) );
  XNOR2X1 U13226 ( .A(n14638), .B(n723), .Y(n14637) );
  NAND2X1 U13227 ( .A(n14639), .B(n14640), .Y(n14628) );
  NAND2X1 U13228 ( .A(n14641), .B(n37453), .Y(n14640) );
  OR2X1 U13229 ( .A(n14642), .B(u_muldiv_dividend_q[17]), .Y(n14641) );
  NAND2X1 U13230 ( .A(u_muldiv_dividend_q[17]), .B(n14642), .Y(n14639) );
  XNOR2X1 U13231 ( .A(u_muldiv_divisor_q[18]), .B(u_muldiv_dividend_q[18]), 
        .Y(n14638) );
  NAND2X1 U13239 ( .A(n14649), .B(n14650), .Y(u_muldiv_N249) );
  NAND2X1 U13240 ( .A(n44611), .B(n14651), .Y(n14650) );
  XOR2X1 U13241 ( .A(n14652), .B(n14642), .Y(n14651) );
  NAND2X1 U13242 ( .A(n14653), .B(n14654), .Y(n14642) );
  NAND2X1 U13243 ( .A(n14655), .B(n37452), .Y(n14654) );
  NAND2X1 U13244 ( .A(n724), .B(n37451), .Y(n14655) );
  NAND2X1 U13245 ( .A(u_muldiv_dividend_q[16]), .B(n14656), .Y(n14653) );
  XNOR2X1 U13246 ( .A(u_muldiv_divisor_q[17]), .B(u_muldiv_dividend_q[17]), 
        .Y(n14652) );
  NAND2X1 U13254 ( .A(n14663), .B(n14664), .Y(u_muldiv_N248) );
  NAND2X1 U13255 ( .A(n44611), .B(n14665), .Y(n14664) );
  XNOR2X1 U13256 ( .A(n14666), .B(n724), .Y(n14665) );
  NAND2X1 U13257 ( .A(n14667), .B(n14668), .Y(n14656) );
  NAND2X1 U13258 ( .A(n14669), .B(n37447), .Y(n14668) );
  NAND2X1 U13259 ( .A(n725), .B(n37446), .Y(n14669) );
  NAND2X1 U13260 ( .A(u_muldiv_dividend_q[15]), .B(n14670), .Y(n14667) );
  XNOR2X1 U13261 ( .A(u_muldiv_divisor_q[16]), .B(u_muldiv_dividend_q[16]), 
        .Y(n14666) );
  NAND2X1 U13269 ( .A(n14677), .B(n14678), .Y(u_muldiv_N247) );
  NAND2X1 U13270 ( .A(n44611), .B(n14679), .Y(n14678) );
  XNOR2X1 U13271 ( .A(n14680), .B(n725), .Y(n14679) );
  NAND2X1 U13272 ( .A(n14681), .B(n14682), .Y(n14670) );
  NAND2X1 U13273 ( .A(n14683), .B(n42547), .Y(n14682) );
  NAND2X1 U13274 ( .A(n726), .B(n37445), .Y(n14683) );
  NAND2X1 U13275 ( .A(u_muldiv_dividend_q[14]), .B(n14684), .Y(n14681) );
  XNOR2X1 U13276 ( .A(u_muldiv_divisor_q[15]), .B(u_muldiv_dividend_q[15]), 
        .Y(n14680) );
  NAND2X1 U13284 ( .A(n14691), .B(n14692), .Y(u_muldiv_N246) );
  NAND2X1 U13285 ( .A(n44611), .B(n14693), .Y(n14692) );
  XNOR2X1 U13286 ( .A(n14694), .B(n726), .Y(n14693) );
  NAND2X1 U13287 ( .A(n14695), .B(n14696), .Y(n14684) );
  NAND2X1 U13288 ( .A(n14697), .B(n37443), .Y(n14696) );
  OR2X1 U13289 ( .A(n14698), .B(u_muldiv_dividend_q[13]), .Y(n14697) );
  NAND2X1 U13290 ( .A(u_muldiv_dividend_q[13]), .B(n14698), .Y(n14695) );
  XNOR2X1 U13291 ( .A(u_muldiv_divisor_q[14]), .B(u_muldiv_dividend_q[14]), 
        .Y(n14694) );
  NAND2X1 U13299 ( .A(n14705), .B(n14706), .Y(u_muldiv_N245) );
  NAND2X1 U13300 ( .A(n44611), .B(n14707), .Y(n14706) );
  XOR2X1 U13301 ( .A(n14708), .B(n14698), .Y(n14707) );
  NAND2X1 U13302 ( .A(n14709), .B(n14710), .Y(n14698) );
  NAND2X1 U13303 ( .A(n14711), .B(n37442), .Y(n14710) );
  NAND2X1 U13304 ( .A(n727), .B(n37441), .Y(n14711) );
  NAND2X1 U13305 ( .A(u_muldiv_dividend_q[12]), .B(n14712), .Y(n14709) );
  XNOR2X1 U13306 ( .A(u_muldiv_divisor_q[13]), .B(u_muldiv_dividend_q[13]), 
        .Y(n14708) );
  NAND2X1 U13314 ( .A(n14719), .B(n14720), .Y(u_muldiv_N244) );
  NAND2X1 U13315 ( .A(n44611), .B(n14721), .Y(n14720) );
  XNOR2X1 U13316 ( .A(n14722), .B(n727), .Y(n14721) );
  NAND2X1 U13317 ( .A(n14723), .B(n14724), .Y(n14712) );
  NAND2X1 U13318 ( .A(n14725), .B(n37440), .Y(n14724) );
  NAND2X1 U13319 ( .A(n728), .B(n37439), .Y(n14725) );
  NAND2X1 U13320 ( .A(u_muldiv_dividend_q[11]), .B(n14726), .Y(n14723) );
  XNOR2X1 U13321 ( .A(u_muldiv_divisor_q[12]), .B(u_muldiv_dividend_q[12]), 
        .Y(n14722) );
  NAND2X1 U13329 ( .A(n14733), .B(n14734), .Y(u_muldiv_N243) );
  NAND2X1 U13330 ( .A(n44611), .B(n14735), .Y(n14734) );
  XNOR2X1 U13331 ( .A(n14736), .B(n728), .Y(n14735) );
  NAND2X1 U13332 ( .A(n14737), .B(n14738), .Y(n14726) );
  NAND2X1 U13333 ( .A(n14739), .B(n42555), .Y(n14738) );
  NAND2X1 U13334 ( .A(n729), .B(n37437), .Y(n14739) );
  NAND2X1 U13335 ( .A(u_muldiv_dividend_q[10]), .B(n14740), .Y(n14737) );
  XNOR2X1 U13336 ( .A(u_muldiv_divisor_q[11]), .B(u_muldiv_dividend_q[11]), 
        .Y(n14736) );
  NAND2X1 U13344 ( .A(n14747), .B(n14748), .Y(u_muldiv_N242) );
  NAND2X1 U13345 ( .A(n44610), .B(n14749), .Y(n14748) );
  XNOR2X1 U13346 ( .A(n14750), .B(n729), .Y(n14749) );
  NAND2X1 U13347 ( .A(n14751), .B(n14752), .Y(n14740) );
  NAND2X1 U13348 ( .A(n14753), .B(n37432), .Y(n14752) );
  OR2X1 U13349 ( .A(n14754), .B(u_muldiv_dividend_q[9]), .Y(n14753) );
  NAND2X1 U13350 ( .A(u_muldiv_dividend_q[9]), .B(n14754), .Y(n14751) );
  XNOR2X1 U13351 ( .A(u_muldiv_divisor_q[10]), .B(u_muldiv_dividend_q[10]), 
        .Y(n14750) );
  NAND2X1 U13359 ( .A(n14761), .B(n14762), .Y(u_muldiv_N241) );
  NAND2X1 U13360 ( .A(n44610), .B(n14763), .Y(n14762) );
  XOR2X1 U13361 ( .A(n14764), .B(n14754), .Y(n14763) );
  NAND2X1 U13362 ( .A(n14765), .B(n14766), .Y(n14754) );
  NAND2X1 U13363 ( .A(n14767), .B(n37429), .Y(n14766) );
  NAND2X1 U13364 ( .A(n730), .B(n37428), .Y(n14767) );
  NAND2X1 U13365 ( .A(u_muldiv_dividend_q[8]), .B(n14768), .Y(n14765) );
  XNOR2X1 U13366 ( .A(u_muldiv_divisor_q[9]), .B(u_muldiv_dividend_q[9]), .Y(
        n14764) );
  NAND2X1 U13374 ( .A(n14775), .B(n14776), .Y(u_muldiv_N240) );
  NAND2X1 U13375 ( .A(n44610), .B(n14777), .Y(n14776) );
  XNOR2X1 U13376 ( .A(n14778), .B(n730), .Y(n14777) );
  NAND2X1 U13377 ( .A(n14779), .B(n14780), .Y(n14768) );
  NAND2X1 U13378 ( .A(n14781), .B(n37427), .Y(n14780) );
  NAND2X1 U13379 ( .A(n731), .B(n37426), .Y(n14781) );
  NAND2X1 U13380 ( .A(u_muldiv_dividend_q[7]), .B(n14782), .Y(n14779) );
  XNOR2X1 U13381 ( .A(u_muldiv_divisor_q[8]), .B(u_muldiv_dividend_q[8]), .Y(
        n14778) );
  NAND2X1 U13389 ( .A(n14789), .B(n14790), .Y(u_muldiv_N239) );
  NAND2X1 U13390 ( .A(n44610), .B(n14791), .Y(n14790) );
  XNOR2X1 U13391 ( .A(n14792), .B(n731), .Y(n14791) );
  NAND2X1 U13392 ( .A(n14793), .B(n14794), .Y(n14782) );
  NAND2X1 U13393 ( .A(n14795), .B(n37424), .Y(n14794) );
  NAND2X1 U13394 ( .A(n732), .B(n37423), .Y(n14795) );
  NAND2X1 U13395 ( .A(u_muldiv_dividend_q[6]), .B(n14796), .Y(n14793) );
  XNOR2X1 U13396 ( .A(u_muldiv_divisor_q[7]), .B(u_muldiv_dividend_q[7]), .Y(
        n14792) );
  NAND2X1 U13404 ( .A(n14803), .B(n14804), .Y(u_muldiv_N238) );
  NAND2X1 U13405 ( .A(n44610), .B(n14805), .Y(n14804) );
  XNOR2X1 U13406 ( .A(n14806), .B(n732), .Y(n14805) );
  NAND2X1 U13407 ( .A(n14807), .B(n14808), .Y(n14796) );
  NAND2X1 U13408 ( .A(n14809), .B(n37422), .Y(n14808) );
  OR2X1 U13409 ( .A(n14810), .B(u_muldiv_dividend_q[5]), .Y(n14809) );
  NAND2X1 U13410 ( .A(u_muldiv_dividend_q[5]), .B(n14810), .Y(n14807) );
  XNOR2X1 U13411 ( .A(u_muldiv_divisor_q[6]), .B(u_muldiv_dividend_q[6]), .Y(
        n14806) );
  NAND2X1 U13419 ( .A(n14817), .B(n14818), .Y(u_muldiv_N237) );
  NAND2X1 U13420 ( .A(n44610), .B(n14819), .Y(n14818) );
  XOR2X1 U13421 ( .A(n14820), .B(n14810), .Y(n14819) );
  NAND2X1 U13422 ( .A(n14821), .B(n14822), .Y(n14810) );
  NAND2X1 U13423 ( .A(n14823), .B(n37421), .Y(n14822) );
  NAND2X1 U13424 ( .A(n14824), .B(n37420), .Y(n14823) );
  OR2X1 U13425 ( .A(n37420), .B(n14824), .Y(n14821) );
  XNOR2X1 U13426 ( .A(u_muldiv_divisor_q[5]), .B(u_muldiv_dividend_q[5]), .Y(
        n14820) );
  NAND2X1 U13434 ( .A(n14831), .B(n14832), .Y(u_muldiv_N236) );
  NAND2X1 U13435 ( .A(n44610), .B(n14833), .Y(n14832) );
  XNOR2X1 U13436 ( .A(n14834), .B(n14824), .Y(n14833) );
  NOR2X1 U13437 ( .A(n14835), .B(n14836), .Y(n14824) );
  AND2X1 U13438 ( .A(n14837), .B(n14838), .Y(n14836) );
  NAND2X1 U13439 ( .A(u_muldiv_divisor_q[3]), .B(n37326), .Y(n14837) );
  XNOR2X1 U13440 ( .A(u_muldiv_divisor_q[4]), .B(u_muldiv_dividend_q[4]), .Y(
        n14834) );
  NAND2X1 U13448 ( .A(n14845), .B(n14846), .Y(u_muldiv_N235) );
  NAND2X1 U13449 ( .A(n44610), .B(n14847), .Y(n14846) );
  NAND2X1 U13450 ( .A(n14848), .B(n14849), .Y(n14847) );
  NAND2X1 U13451 ( .A(n14835), .B(n14838), .Y(n14849) );
  NOR2X1 U13452 ( .A(n14850), .B(n14851), .Y(n14848) );
  NOR2X1 U13453 ( .A(n37438), .B(n14852), .Y(n14851) );
  XNOR2X1 U13454 ( .A(u_muldiv_dividend_q[3]), .B(n14838), .Y(n14852) );
  NOR2X1 U13455 ( .A(n14838), .B(n14853), .Y(n14850) );
  NAND2X1 U13456 ( .A(n37326), .B(n37438), .Y(n14853) );
  OR2X1 U13457 ( .A(n14854), .B(n14855), .Y(n14838) );
  AND2X1 U13458 ( .A(n14856), .B(n14857), .Y(n14855) );
  NAND2X1 U13459 ( .A(u_muldiv_divisor_q[2]), .B(n37325), .Y(n14856) );
  NAND2X1 U13467 ( .A(n14864), .B(n14865), .Y(u_muldiv_N234) );
  NAND2X1 U13468 ( .A(n44610), .B(n14866), .Y(n14865) );
  NAND2X1 U13469 ( .A(n14867), .B(n14868), .Y(n14866) );
  NAND2X1 U13470 ( .A(n14854), .B(n14857), .Y(n14868) );
  NOR2X1 U13471 ( .A(n14869), .B(n14870), .Y(n14867) );
  NOR2X1 U13472 ( .A(n37435), .B(n14871), .Y(n14870) );
  XNOR2X1 U13473 ( .A(u_muldiv_dividend_q[2]), .B(n14857), .Y(n14871) );
  NOR2X1 U13474 ( .A(n14857), .B(n14872), .Y(n14869) );
  NAND2X1 U13475 ( .A(n37325), .B(n37435), .Y(n14872) );
  NAND2X1 U13483 ( .A(n14878), .B(n14879), .Y(u_muldiv_N233) );
  NAND2X1 U13484 ( .A(n44610), .B(n14880), .Y(n14879) );
  XNOR2X1 U13485 ( .A(n14881), .B(n14882), .Y(n14880) );
  XNOR2X1 U13486 ( .A(n37419), .B(u_muldiv_dividend_q[1]), .Y(n14882) );
  NAND2X1 U13494 ( .A(n44610), .B(n14891), .Y(n14890) );
  NAND2X1 U13495 ( .A(n14881), .B(n14892), .Y(n14891) );
  NAND2X1 U13496 ( .A(u_muldiv_dividend_q[0]), .B(n37418), .Y(n14892) );
  NOR2X1 U13503 ( .A(n37587), .B(n73548), .Y(u_mmu_N250) );
  NOR2X1 U13504 ( .A(n37587), .B(n73549), .Y(u_mmu_N249) );
  NOR2X1 U13535 ( .A(n37587), .B(n432), .Y(u_mmu_N238) );
  NOR2X1 U13536 ( .A(n37587), .B(n436), .Y(u_mmu_N237) );
  NOR2X1 U13537 ( .A(n37587), .B(n437), .Y(u_mmu_N236) );
  NOR2X1 U13538 ( .A(n37587), .B(n438), .Y(u_mmu_N235) );
  NOR2X1 U13867 ( .A(n15220), .B(n15221), .Y(u_lsu_N231) );
  NAND2X1 U13868 ( .A(n73542), .B(n73394), .Y(n15221) );
  NOR2X1 U13999 ( .A(n15319), .B(n15320), .Y(n15318) );
  NAND2X1 U14081 ( .A(n15402), .B(n15403), .Y(n15401) );
  NAND2X1 U14082 ( .A(n73511), .B(n15404), .Y(n15403) );
  NOR2X1 U14083 ( .A(n15405), .B(n15406), .Y(n15402) );
  NOR2X1 U14084 ( .A(n15407), .B(n15408), .Y(n15406) );
  NOR2X1 U14085 ( .A(n15409), .B(n15410), .Y(n15405) );
  NAND2X1 U14086 ( .A(n15411), .B(n15412), .Y(n15400) );
  NAND2X1 U14087 ( .A(n15413), .B(n15414), .Y(n15412) );
  NAND2X1 U14088 ( .A(n15415), .B(n15416), .Y(n15413) );
  NOR2X1 U14089 ( .A(n15417), .B(n15418), .Y(n15415) );
  NOR2X1 U14090 ( .A(n42211), .B(n15420), .Y(n15418) );
  NOR2X1 U14091 ( .A(n73481), .B(n15421), .Y(n15417) );
  NOR2X1 U14092 ( .A(n980), .B(n15422), .Y(n15421) );
  NOR2X1 U14093 ( .A(n50), .B(n15423), .Y(n15411) );
  NOR2X1 U14094 ( .A(n15424), .B(n15414), .Y(n15423) );
  NOR2X1 U14095 ( .A(n15425), .B(n15426), .Y(n15424) );
  NOR2X1 U14096 ( .A(n73481), .B(n42211), .Y(n15426) );
  AND2X1 U14101 ( .A(n15422), .B(n73481), .Y(n15425) );
  NAND2X1 U14106 ( .A(n15438), .B(n15439), .Y(n15437) );
  NAND2X1 U14107 ( .A(n42942), .B(n15441), .Y(n15439) );
  NAND2X1 U14108 ( .A(n15442), .B(n15443), .Y(n15438) );
  NAND2X1 U14109 ( .A(n15444), .B(n15445), .Y(n15436) );
  NAND2X1 U14110 ( .A(n73510), .B(n15447), .Y(n15445) );
  NOR2X1 U14111 ( .A(n15448), .B(n15449), .Y(n15444) );
  NOR2X1 U14112 ( .A(n15450), .B(n43010), .Y(n15449) );
  NOR2X1 U14113 ( .A(n42454), .B(n15453), .Y(n15448) );
  NOR2X1 U14118 ( .A(n15460), .B(n15461), .Y(n15458) );
  NOR2X1 U14119 ( .A(n15462), .B(n42946), .Y(n15461) );
  NOR2X1 U14120 ( .A(n15464), .B(n15465), .Y(n15460) );
  NAND2X1 U14121 ( .A(n15466), .B(n15467), .Y(n15456) );
  NOR2X1 U14122 ( .A(n50), .B(n15468), .Y(n15467) );
  NOR2X1 U14123 ( .A(n15469), .B(n15447), .Y(n15468) );
  NOR2X1 U14124 ( .A(n15470), .B(n15471), .Y(n15469) );
  NOR2X1 U14125 ( .A(n73493), .B(n42305), .Y(n15471) );
  AND2X1 U14126 ( .A(n15473), .B(n73493), .Y(n15470) );
  NOR2X1 U14127 ( .A(n15474), .B(n15475), .Y(n15466) );
  NOR2X1 U14128 ( .A(n42305), .B(n15476), .Y(n15475) );
  NOR2X1 U14133 ( .A(n73494), .B(n15482), .Y(n15474) );
  NOR2X1 U14134 ( .A(n15483), .B(n42971), .Y(n15482) );
  NOR2X1 U14135 ( .A(n73493), .B(n15484), .Y(n15483) );
  NOR2X1 U14136 ( .A(n980), .B(n15473), .Y(n15484) );
  NAND2X1 U14141 ( .A(n15489), .B(n15490), .Y(n15488) );
  OR2X1 U14142 ( .A(n40678), .B(n15492), .Y(n15490) );
  NOR2X1 U14143 ( .A(n15493), .B(n15494), .Y(n15489) );
  NOR2X1 U14144 ( .A(n15495), .B(n15496), .Y(n15494) );
  NOR2X1 U14145 ( .A(n15497), .B(n15498), .Y(n15493) );
  NAND2X1 U14146 ( .A(n15499), .B(n15500), .Y(n15487) );
  NAND2X1 U14147 ( .A(n37341), .B(n15501), .Y(n15500) );
  NOR2X1 U14148 ( .A(n15502), .B(n15503), .Y(n15499) );
  NOR2X1 U14149 ( .A(n15504), .B(n15505), .Y(n15503) );
  NOR2X1 U14150 ( .A(n226), .B(n43007), .Y(n15502) );
  NAND2X1 U14153 ( .A(n15510), .B(n15511), .Y(n15509) );
  NOR2X1 U14154 ( .A(n15512), .B(n15513), .Y(n15511) );
  NOR2X1 U14155 ( .A(n15514), .B(n43011), .Y(n15513) );
  NOR2X1 U14156 ( .A(n15515), .B(n43008), .Y(n15512) );
  NOR2X1 U14157 ( .A(n15516), .B(n15517), .Y(n15510) );
  NOR2X1 U14158 ( .A(n227), .B(n15408), .Y(n15517) );
  NOR2X1 U14159 ( .A(n256), .B(n15491), .Y(n15516) );
  NAND2X1 U14160 ( .A(n15518), .B(n15519), .Y(n15508) );
  NOR2X1 U14161 ( .A(n50), .B(n15520), .Y(n15519) );
  NOR2X1 U14162 ( .A(n15521), .B(n15441), .Y(n15520) );
  NOR2X1 U14163 ( .A(n15522), .B(n15523), .Y(n15521) );
  AND2X1 U14164 ( .A(n15524), .B(n15525), .Y(n15523) );
  NOR2X1 U14165 ( .A(n15526), .B(n15524), .Y(n15522) );
  NOR2X1 U14166 ( .A(n15527), .B(n15528), .Y(n15518) );
  NOR2X1 U14167 ( .A(n15529), .B(n15530), .Y(n15528) );
  NOR2X1 U14168 ( .A(n73484), .B(n15531), .Y(n15527) );
  NOR2X1 U14169 ( .A(n361), .B(n15532), .Y(n15531) );
  NAND2X1 U14170 ( .A(n15533), .B(n15534), .Y(n15532) );
  NAND2X1 U14171 ( .A(n15535), .B(n15524), .Y(n15534) );
  NAND2X1 U14172 ( .A(n15526), .B(n42970), .Y(n15535) );
  NAND2X1 U14176 ( .A(n73483), .B(n15525), .Y(n15533) );
  NAND2X1 U14182 ( .A(n15546), .B(n15547), .Y(n15545) );
  NOR2X1 U14183 ( .A(n15548), .B(n15549), .Y(n15547) );
  NOR2X1 U14184 ( .A(n73482), .B(n42986), .Y(n15549) );
  NOR2X1 U14185 ( .A(n73490), .B(n363), .Y(n15548) );
  NOR2X1 U14186 ( .A(n15550), .B(n15551), .Y(n15546) );
  NOR2X1 U14187 ( .A(n73494), .B(n360), .Y(n15551) );
  NOR2X1 U14188 ( .A(n73480), .B(n42984), .Y(n15550) );
  NAND2X1 U14189 ( .A(n15552), .B(n15553), .Y(n15544) );
  NOR2X1 U14190 ( .A(n15554), .B(n15555), .Y(n15553) );
  NOR2X1 U14191 ( .A(n15556), .B(n15496), .Y(n15555) );
  NOR2X1 U14192 ( .A(n378), .B(n15463), .Y(n15554) );
  NOR2X1 U14193 ( .A(n15557), .B(n15558), .Y(n15552) );
  NOR2X1 U14194 ( .A(n73488), .B(n362), .Y(n15558) );
  NOR2X1 U14195 ( .A(n73486), .B(n364), .Y(n15557) );
  NAND2X1 U14198 ( .A(n15563), .B(n15564), .Y(n15562) );
  NOR2X1 U14199 ( .A(n15565), .B(n15566), .Y(n15564) );
  NOR2X1 U14200 ( .A(n343), .B(n15567), .Y(n15566) );
  NOR2X1 U14201 ( .A(n73485), .B(n15569), .Y(n15565) );
  NOR2X1 U14202 ( .A(n37560), .B(n15571), .Y(n15569) );
  NAND2X1 U14203 ( .A(n15572), .B(n15573), .Y(n15571) );
  NAND2X1 U14204 ( .A(n15574), .B(n15443), .Y(n15573) );
  OR2X1 U14205 ( .A(n15575), .B(n980), .Y(n15574) );
  NAND2X1 U14206 ( .A(n73486), .B(n15568), .Y(n15572) );
  NOR2X1 U14211 ( .A(n15581), .B(n15582), .Y(n15563) );
  NOR2X1 U14212 ( .A(n15583), .B(n15505), .Y(n15582) );
  NOR2X1 U14213 ( .A(n15584), .B(n15498), .Y(n15581) );
  NAND2X1 U14214 ( .A(n15585), .B(n15586), .Y(n15561) );
  NOR2X1 U14215 ( .A(n49), .B(n15587), .Y(n15586) );
  NOR2X1 U14216 ( .A(n15443), .B(n15588), .Y(n15587) );
  NAND2X1 U14217 ( .A(n73485), .B(n15575), .Y(n15588) );
  NOR2X1 U14221 ( .A(n15591), .B(n15592), .Y(n15585) );
  NOR2X1 U14222 ( .A(n43009), .B(n15593), .Y(n15592) );
  NOR2X1 U14223 ( .A(n15594), .B(n15595), .Y(n15591) );
  NAND2X1 U14225 ( .A(n15598), .B(n15599), .Y(n15597) );
  NAND2X1 U14226 ( .A(n15600), .B(n15414), .Y(n15599) );
  NOR2X1 U14227 ( .A(n15601), .B(n15602), .Y(n15598) );
  NOR2X1 U14228 ( .A(n73494), .B(n42986), .Y(n15602) );
  NOR2X1 U14229 ( .A(n255), .B(n15491), .Y(n15601) );
  NAND2X1 U14230 ( .A(n15603), .B(n15604), .Y(n15596) );
  NOR2X1 U14231 ( .A(n15605), .B(n15606), .Y(n15604) );
  NOR2X1 U14232 ( .A(n73397), .B(n42946), .Y(n15606) );
  NOR2X1 U14233 ( .A(n15607), .B(n15496), .Y(n15605) );
  NOR2X1 U14234 ( .A(n15608), .B(n15609), .Y(n15603) );
  NOR2X1 U14235 ( .A(n216), .B(n43007), .Y(n15609) );
  NOR2X1 U14236 ( .A(n15610), .B(n15465), .Y(n15608) );
  NAND2X1 U14239 ( .A(n15615), .B(n15616), .Y(n15614) );
  NOR2X1 U14240 ( .A(n15617), .B(n15618), .Y(n15616) );
  NOR2X1 U14241 ( .A(n257), .B(n15496), .Y(n15618) );
  NOR2X1 U14242 ( .A(n15619), .B(n43008), .Y(n15617) );
  NOR2X1 U14243 ( .A(n15620), .B(n15621), .Y(n15615) );
  NOR2X1 U14244 ( .A(n55), .B(n15529), .Y(n15621) );
  NOR2X1 U14245 ( .A(n15407), .B(n40678), .Y(n15620) );
  NAND2X1 U14246 ( .A(n15622), .B(n15623), .Y(n15613) );
  NOR2X1 U14247 ( .A(n15624), .B(n15625), .Y(n15623) );
  NAND2X1 U14248 ( .A(n15626), .B(n15627), .Y(n15625) );
  NAND2X1 U14249 ( .A(n73488), .B(n15628), .Y(n15626) );
  NAND2X1 U14250 ( .A(n15629), .B(n15630), .Y(n15628) );
  NAND2X1 U14251 ( .A(n73487), .B(n15631), .Y(n15630) );
  NAND2X1 U14252 ( .A(n15632), .B(n15633), .Y(n15629) );
  NOR2X1 U14253 ( .A(n73488), .B(n15634), .Y(n15624) );
  NOR2X1 U14254 ( .A(n42971), .B(n15635), .Y(n15634) );
  NAND2X1 U14255 ( .A(n15636), .B(n15637), .Y(n15635) );
  NAND2X1 U14256 ( .A(n15638), .B(n15633), .Y(n15637) );
  OR2X1 U14257 ( .A(n15631), .B(n980), .Y(n15638) );
  NAND2X1 U14261 ( .A(n73487), .B(n15632), .Y(n15636) );
  NOR2X1 U14266 ( .A(n15646), .B(n15647), .Y(n15622) );
  NOR2X1 U14267 ( .A(n15648), .B(n43010), .Y(n15647) );
  NOR2X1 U14268 ( .A(n73482), .B(n15649), .Y(n15646) );
  NAND2X1 U14270 ( .A(n15652), .B(n15653), .Y(n15651) );
  NOR2X1 U14271 ( .A(n15654), .B(n15655), .Y(n15653) );
  NOR2X1 U14272 ( .A(n73484), .B(n42986), .Y(n15655) );
  NOR2X1 U14273 ( .A(n73491), .B(n363), .Y(n15654) );
  NOR2X1 U14274 ( .A(n15656), .B(n15657), .Y(n15652) );
  NOR2X1 U14275 ( .A(n73486), .B(n42991), .Y(n15657) );
  NOR2X1 U14276 ( .A(n73494), .B(n42985), .Y(n15656) );
  NAND2X1 U14277 ( .A(n15658), .B(n15659), .Y(n15650) );
  NOR2X1 U14278 ( .A(n15660), .B(n15661), .Y(n15659) );
  NOR2X1 U14279 ( .A(n15450), .B(n15408), .Y(n15661) );
  NOR2X1 U14280 ( .A(n42454), .B(n15463), .Y(n15660) );
  NOR2X1 U14281 ( .A(n15662), .B(n15663), .Y(n15658) );
  NOR2X1 U14282 ( .A(n73495), .B(n42943), .Y(n15663) );
  NOR2X1 U14283 ( .A(n73490), .B(n364), .Y(n15662) );
  NOR2X1 U14290 ( .A(n15673), .B(n15674), .Y(n15668) );
  NOR2X1 U14291 ( .A(n73492), .B(n363), .Y(n15674) );
  NOR2X1 U14292 ( .A(n73491), .B(n42943), .Y(n15673) );
  NAND2X1 U14293 ( .A(n15675), .B(n15676), .Y(n15666) );
  NOR2X1 U14294 ( .A(n49), .B(n15677), .Y(n15676) );
  NOR2X1 U14295 ( .A(n15678), .B(n15679), .Y(n15677) );
  NOR2X1 U14296 ( .A(n15680), .B(n15681), .Y(n15678) );
  AND2X1 U14297 ( .A(n15682), .B(n15683), .Y(n15681) );
  NOR2X1 U14298 ( .A(n15684), .B(n15682), .Y(n15680) );
  NOR2X1 U14299 ( .A(n15685), .B(n15686), .Y(n15675) );
  NOR2X1 U14300 ( .A(n15687), .B(n15505), .Y(n15686) );
  NOR2X1 U14301 ( .A(n73490), .B(n15688), .Y(n15685) );
  NOR2X1 U14302 ( .A(n42972), .B(n15689), .Y(n15688) );
  NAND2X1 U14303 ( .A(n15690), .B(n15691), .Y(n15689) );
  NAND2X1 U14304 ( .A(n15692), .B(n15682), .Y(n15691) );
  NAND2X1 U14305 ( .A(n15684), .B(n42969), .Y(n15692) );
  NAND2X1 U14309 ( .A(n73489), .B(n15683), .Y(n15690) );
  NAND2X1 U14315 ( .A(n15702), .B(n15703), .Y(n15701) );
  NOR2X1 U14316 ( .A(n15704), .B(n15705), .Y(n15703) );
  NOR2X1 U14317 ( .A(n73488), .B(n42990), .Y(n15705) );
  NOR2X1 U14318 ( .A(n15495), .B(n15529), .Y(n15704) );
  NOR2X1 U14319 ( .A(n15706), .B(n15707), .Y(n15702) );
  NOR2X1 U14320 ( .A(n15492), .B(n15496), .Y(n15707) );
  NOR2X1 U14321 ( .A(n226), .B(n15491), .Y(n15706) );
  NAND2X1 U14322 ( .A(n15708), .B(n15709), .Y(n15700) );
  NOR2X1 U14323 ( .A(n15710), .B(n15711), .Y(n15709) );
  NOR2X1 U14324 ( .A(n215), .B(n43007), .Y(n15711) );
  NOR2X1 U14325 ( .A(n73486), .B(n42986), .Y(n15710) );
  NOR2X1 U14326 ( .A(n15712), .B(n15713), .Y(n15708) );
  NOR2X1 U14327 ( .A(n73484), .B(n42984), .Y(n15713) );
  NOR2X1 U14328 ( .A(n15504), .B(n43011), .Y(n15712) );
  NAND2X1 U14331 ( .A(n15718), .B(n15719), .Y(n15717) );
  NOR2X1 U14332 ( .A(n15720), .B(n15721), .Y(n15719) );
  NOR2X1 U14333 ( .A(n73494), .B(n15722), .Y(n15721) );
  NOR2X1 U14334 ( .A(n73482), .B(n15723), .Y(n15720) );
  NOR2X1 U14335 ( .A(n15724), .B(n15725), .Y(n15718) );
  NOR2X1 U14336 ( .A(n15515), .B(n43010), .Y(n15725) );
  AND2X1 U14337 ( .A(n15726), .B(n15727), .Y(n15515) );
  NOR2X1 U14339 ( .A(n73484), .B(n15649), .Y(n15724) );
  NAND2X1 U14340 ( .A(n15729), .B(n15730), .Y(n15716) );
  NOR2X1 U14341 ( .A(n15731), .B(n15732), .Y(n15730) );
  NAND2X1 U14342 ( .A(n15733), .B(n15627), .Y(n15732) );
  NAND2X1 U14343 ( .A(n50), .B(n15734), .Y(n15627) );
  NAND2X1 U14344 ( .A(n15736), .B(n73396), .Y(n15733) );
  NOR2X1 U14345 ( .A(n15737), .B(n15594), .Y(n15736) );
  NOR2X1 U14346 ( .A(n15738), .B(n15739), .Y(n15731) );
  NOR2X1 U14347 ( .A(n15740), .B(n15741), .Y(n15738) );
  AND2X1 U14348 ( .A(n15742), .B(n15743), .Y(n15741) );
  NOR2X1 U14349 ( .A(n15744), .B(n15742), .Y(n15740) );
  NOR2X1 U14350 ( .A(n15745), .B(n15746), .Y(n15729) );
  NOR2X1 U14351 ( .A(n73480), .B(n15747), .Y(n15746) );
  NOR2X1 U14352 ( .A(n73495), .B(n15748), .Y(n15745) );
  NOR2X1 U14353 ( .A(n15749), .B(n15750), .Y(n15748) );
  NAND2X1 U14354 ( .A(n15751), .B(n15752), .Y(n15750) );
  NAND2X1 U14355 ( .A(n15753), .B(n15742), .Y(n15752) );
  NAND2X1 U14356 ( .A(n15744), .B(n42970), .Y(n15753) );
  NAND2X1 U14360 ( .A(n73525), .B(n15743), .Y(n15751) );
  NAND2X1 U14366 ( .A(n15763), .B(n15764), .Y(n15762) );
  NOR2X1 U14367 ( .A(n15765), .B(n15766), .Y(n15764) );
  NOR2X1 U14368 ( .A(n73488), .B(n42986), .Y(n15766) );
  NOR2X1 U14369 ( .A(n15556), .B(n15529), .Y(n15765) );
  NOR2X1 U14370 ( .A(n15767), .B(n15768), .Y(n15763) );
  NOR2X1 U14371 ( .A(n73490), .B(n360), .Y(n15768) );
  NOR2X1 U14372 ( .A(n73486), .B(n42985), .Y(n15767) );
  NAND2X1 U14373 ( .A(n15769), .B(n15770), .Y(n15761) );
  NOR2X1 U14374 ( .A(n15771), .B(n15772), .Y(n15770) );
  NOR2X1 U14375 ( .A(n256), .B(n15496), .Y(n15772) );
  NOR2X1 U14376 ( .A(n15514), .B(n15408), .Y(n15771) );
  NOR2X1 U14377 ( .A(n15773), .B(n15774), .Y(n15769) );
  NOR2X1 U14378 ( .A(n378), .B(n40684), .Y(n15774) );
  NOR2X1 U14379 ( .A(n227), .B(n15491), .Y(n15773) );
  NOR2X1 U14384 ( .A(n15782), .B(n15783), .Y(n15779) );
  NAND2X1 U14387 ( .A(n15788), .B(n15789), .Y(n15777) );
  NOR2X1 U14388 ( .A(n54), .B(n15790), .Y(n15789) );
  NOR2X1 U14389 ( .A(n73438), .B(n15791), .Y(n15790) );
  NOR2X1 U14390 ( .A(n15792), .B(n42972), .Y(n15791) );
  NOR2X1 U14391 ( .A(n73437), .B(n42969), .Y(n15792) );
  NOR2X1 U14392 ( .A(n15793), .B(n15794), .Y(n15788) );
  NOR2X1 U14394 ( .A(n15797), .B(n15798), .Y(n15795) );
  NAND2X1 U14395 ( .A(n15799), .B(n15800), .Y(n15798) );
  NAND2X1 U14396 ( .A(n42958), .B(n15801), .Y(n15800) );
  NAND2X1 U14397 ( .A(n73512), .B(n15802), .Y(n15799) );
  NAND2X1 U14398 ( .A(n15803), .B(n15804), .Y(n15797) );
  NAND2X1 U14399 ( .A(n371), .B(n15728), .Y(n15804) );
  NAND2X1 U14400 ( .A(n368), .B(n15805), .Y(n15803) );
  NOR2X1 U14403 ( .A(n15808), .B(n15809), .Y(n15807) );
  AND2X1 U14404 ( .A(n15810), .B(n15811), .Y(n15809) );
  NOR2X1 U14405 ( .A(n73439), .B(n15812), .Y(n15808) );
  NOR2X1 U14406 ( .A(n15811), .B(n15810), .Y(n15812) );
  NOR2X1 U14410 ( .A(n15818), .B(n15819), .Y(n15815) );
  NOR2X1 U14411 ( .A(n73442), .B(n362), .Y(n15819) );
  NOR2X1 U14412 ( .A(n73439), .B(n364), .Y(n15818) );
  NAND2X1 U14413 ( .A(n15820), .B(n15821), .Y(n15813) );
  NOR2X1 U14414 ( .A(n15822), .B(n15823), .Y(n15821) );
  NOR2X1 U14415 ( .A(n378), .B(n15824), .Y(n15823) );
  NOR2X1 U14417 ( .A(n15826), .B(n15827), .Y(n15820) );
  NOR2X1 U14418 ( .A(n73446), .B(n15672), .Y(n15827) );
  NOR2X1 U14419 ( .A(n15828), .B(n15829), .Y(n15826) );
  NOR2X1 U14424 ( .A(n15837), .B(n15838), .Y(n15834) );
  AND2X1 U14427 ( .A(n15839), .B(n15840), .Y(n15784) );
  NOR2X1 U14428 ( .A(n15841), .B(n15842), .Y(n15840) );
  NAND2X1 U14429 ( .A(n15843), .B(n15844), .Y(n15842) );
  NAND2X1 U14430 ( .A(n371), .B(n15845), .Y(n15844) );
  NAND2X1 U14431 ( .A(n368), .B(n15846), .Y(n15843) );
  NOR2X1 U14432 ( .A(n73464), .B(n42959), .Y(n15841) );
  NOR2X1 U14433 ( .A(n15848), .B(n15849), .Y(n15839) );
  NOR2X1 U14434 ( .A(n73456), .B(n42945), .Y(n15849) );
  NOR2X1 U14435 ( .A(n73448), .B(n42946), .Y(n15848) );
  NAND2X1 U14436 ( .A(n15850), .B(n15851), .Y(n15832) );
  NOR2X1 U14437 ( .A(n15852), .B(n15853), .Y(n15851) );
  NOR2X1 U14438 ( .A(n73439), .B(n15854), .Y(n15853) );
  NOR2X1 U14439 ( .A(n361), .B(n15855), .Y(n15854) );
  NAND2X1 U14440 ( .A(n15856), .B(n15857), .Y(n15855) );
  NAND2X1 U14441 ( .A(n15858), .B(n15810), .Y(n15857) );
  NAND2X1 U14442 ( .A(n42189), .B(n42969), .Y(n15858) );
  NAND2X1 U14443 ( .A(n73440), .B(n15860), .Y(n15856) );
  NOR2X1 U14444 ( .A(n15861), .B(n15862), .Y(n15852) );
  NOR2X1 U14445 ( .A(n15863), .B(n15864), .Y(n15861) );
  AND2X1 U14446 ( .A(n15810), .B(n15860), .Y(n15864) );
  NOR2X1 U14451 ( .A(n42189), .B(n15810), .Y(n15863) );
  NAND2X1 U14454 ( .A(n15871), .B(n15872), .Y(n15811) );
  NAND2X1 U14455 ( .A(n15873), .B(n15874), .Y(n15872) );
  OR2X1 U14456 ( .A(n15875), .B(n15876), .Y(n15873) );
  NAND2X1 U14457 ( .A(n15876), .B(n15875), .Y(n15871) );
  NOR2X1 U14459 ( .A(n15877), .B(n15878), .Y(n15850) );
  NOR2X1 U14461 ( .A(n73454), .B(n15880), .Y(n15877) );
  NAND2X1 U14463 ( .A(n15883), .B(n15884), .Y(n15882) );
  NOR2X1 U14464 ( .A(n15885), .B(n15886), .Y(n15883) );
  NOR2X1 U14465 ( .A(n73438), .B(n42991), .Y(n15886) );
  NOR2X1 U14466 ( .A(n73523), .B(n15887), .Y(n15885) );
  NAND2X1 U14467 ( .A(n15888), .B(n15889), .Y(n15881) );
  NOR2X1 U14468 ( .A(n15890), .B(n15891), .Y(n15889) );
  NOR2X1 U14469 ( .A(n15610), .B(n15829), .Y(n15891) );
  NOR2X1 U14470 ( .A(n73397), .B(n15824), .Y(n15890) );
  NOR2X1 U14471 ( .A(n15892), .B(n15893), .Y(n15888) );
  NOR2X1 U14472 ( .A(n73446), .B(n363), .Y(n15893) );
  NOR2X1 U14473 ( .A(n73442), .B(n364), .Y(n15892) );
  NAND2X1 U14476 ( .A(n15898), .B(n15899), .Y(n15897) );
  NOR2X1 U14477 ( .A(n15900), .B(n15901), .Y(n15899) );
  NOR2X1 U14478 ( .A(n15584), .B(n43008), .Y(n15901) );
  NOR2X1 U14479 ( .A(n42450), .B(n42458), .Y(n15584) );
  NOR2X1 U14480 ( .A(n73494), .B(n15723), .Y(n15900) );
  NOR2X1 U14481 ( .A(n15904), .B(n15905), .Y(n15898) );
  NOR2X1 U14482 ( .A(n73492), .B(n40674), .Y(n15905) );
  NOR2X1 U14483 ( .A(n15583), .B(n43011), .Y(n15904) );
  AND2X1 U14484 ( .A(n15906), .B(n15907), .Y(n15583) );
  NOR2X1 U14485 ( .A(n42457), .B(n15909), .Y(n15907) );
  NOR2X1 U14487 ( .A(n42322), .B(n42326), .Y(n15906) );
  NAND2X1 U14488 ( .A(n15912), .B(n15913), .Y(n15896) );
  NOR2X1 U14489 ( .A(n15914), .B(n15915), .Y(n15913) );
  NOR2X1 U14490 ( .A(n15916), .B(n15734), .Y(n15915) );
  NOR2X1 U14491 ( .A(n15917), .B(n15918), .Y(n15916) );
  AND2X1 U14492 ( .A(n15919), .B(n15920), .Y(n15918) );
  NOR2X1 U14493 ( .A(n15921), .B(n15919), .Y(n15917) );
  NOR2X1 U14494 ( .A(n43006), .B(n15593), .Y(n15914) );
  NOR2X1 U14496 ( .A(n15922), .B(n15923), .Y(n15912) );
  NOR2X1 U14497 ( .A(n73482), .B(n15747), .Y(n15923) );
  NOR2X1 U14498 ( .A(n73433), .B(n15924), .Y(n15922) );
  NOR2X1 U14499 ( .A(n15925), .B(n15926), .Y(n15924) );
  NAND2X1 U14500 ( .A(n15927), .B(n15928), .Y(n15926) );
  NAND2X1 U14501 ( .A(n15929), .B(n15919), .Y(n15928) );
  NAND2X1 U14502 ( .A(n15921), .B(n42970), .Y(n15929) );
  NAND2X1 U14506 ( .A(n73491), .B(n15920), .Y(n15927) );
  NOR2X1 U14511 ( .A(n48), .B(n15594), .Y(n15925) );
  NAND2X1 U14513 ( .A(n15939), .B(n15940), .Y(n15938) );
  NOR2X1 U14514 ( .A(n15941), .B(n15942), .Y(n15940) );
  NOR2X1 U14515 ( .A(n73488), .B(n358), .Y(n15942) );
  NOR2X1 U14516 ( .A(n73490), .B(n42988), .Y(n15941) );
  NOR2X1 U14517 ( .A(n15943), .B(n15944), .Y(n15939) );
  NOR2X1 U14518 ( .A(n73495), .B(n42990), .Y(n15944) );
  NOR2X1 U14519 ( .A(n15416), .B(n73491), .Y(n15943) );
  NOR2X1 U14522 ( .A(n15607), .B(n15529), .Y(n15948) );
  NOR2X1 U14524 ( .A(n15949), .B(n15950), .Y(n15945) );
  NOR2X1 U14525 ( .A(n255), .B(n15496), .Y(n15950) );
  NOR2X1 U14526 ( .A(n216), .B(n15491), .Y(n15949) );
  NAND2X1 U14529 ( .A(n15955), .B(n15956), .Y(n15954) );
  NOR2X1 U14530 ( .A(n15957), .B(n15958), .Y(n15956) );
  AND2X1 U14531 ( .A(n73511), .B(n37556), .Y(n15958) );
  AND2X1 U14533 ( .A(n15961), .B(n15962), .Y(n15879) );
  NOR2X1 U14534 ( .A(n15963), .B(n15964), .Y(n15962) );
  NOR2X1 U14535 ( .A(n73478), .B(n15965), .Y(n15964) );
  NOR2X1 U14536 ( .A(n73484), .B(n15966), .Y(n15963) );
  NOR2X1 U14537 ( .A(n15967), .B(n15968), .Y(n15961) );
  NOR2X1 U14538 ( .A(n73462), .B(n42944), .Y(n15968) );
  NOR2X1 U14539 ( .A(n73470), .B(n42960), .Y(n15967) );
  NOR2X1 U14540 ( .A(n15969), .B(n15970), .Y(n15955) );
  NOR2X1 U14544 ( .A(n15973), .B(n15974), .Y(n15972) );
  NAND2X1 U14545 ( .A(n15975), .B(n15976), .Y(n15974) );
  NAND2X1 U14546 ( .A(n371), .B(n15414), .Y(n15976) );
  NAND2X1 U14547 ( .A(n368), .B(n15977), .Y(n15975) );
  NOR2X1 U14548 ( .A(n73466), .B(n42959), .Y(n15973) );
  NOR2X1 U14549 ( .A(n15978), .B(n15979), .Y(n15971) );
  NOR2X1 U14550 ( .A(n73458), .B(n15453), .Y(n15979) );
  NOR2X1 U14551 ( .A(n73450), .B(n15463), .Y(n15978) );
  NAND2X1 U14552 ( .A(n15980), .B(n15981), .Y(n15953) );
  NOR2X1 U14553 ( .A(n15982), .B(n15983), .Y(n15981) );
  NOR2X1 U14554 ( .A(n73442), .B(n15984), .Y(n15983) );
  NOR2X1 U14555 ( .A(n42971), .B(n15985), .Y(n15984) );
  NAND2X1 U14556 ( .A(n15986), .B(n15987), .Y(n15985) );
  NAND2X1 U14557 ( .A(n15988), .B(n15875), .Y(n15987) );
  NAND2X1 U14558 ( .A(n42193), .B(n42969), .Y(n15988) );
  NAND2X1 U14559 ( .A(n73441), .B(n15990), .Y(n15986) );
  NOR2X1 U14560 ( .A(n15991), .B(n15874), .Y(n15982) );
  NOR2X1 U14561 ( .A(n15992), .B(n15993), .Y(n15991) );
  AND2X1 U14562 ( .A(n15875), .B(n15990), .Y(n15993) );
  NOR2X1 U14567 ( .A(n42193), .B(n15875), .Y(n15992) );
  NAND2X1 U14570 ( .A(n16000), .B(n16001), .Y(n15876) );
  NAND2X1 U14571 ( .A(n16002), .B(n16003), .Y(n16001) );
  OR2X1 U14572 ( .A(n16004), .B(n16005), .Y(n16002) );
  NAND2X1 U14573 ( .A(n16005), .B(n16004), .Y(n16000) );
  NOR2X1 U14575 ( .A(n16006), .B(n16007), .Y(n15980) );
  NOR2X1 U14576 ( .A(n73456), .B(n15880), .Y(n16007) );
  NOR2X1 U14578 ( .A(n16009), .B(n16010), .Y(n16008) );
  NAND2X1 U14579 ( .A(n16011), .B(n16012), .Y(n16010) );
  NAND2X1 U14580 ( .A(n371), .B(n15443), .Y(n16012) );
  NAND2X1 U14581 ( .A(n368), .B(n15845), .Y(n16011) );
  NAND2X1 U14583 ( .A(n16015), .B(n16016), .Y(n16014) );
  NOR2X1 U14584 ( .A(n16017), .B(n16018), .Y(n16016) );
  NOR2X1 U14585 ( .A(n73438), .B(n42987), .Y(n16018) );
  NOR2X1 U14586 ( .A(n15887), .B(n42984), .Y(n16017) );
  NOR2X1 U14587 ( .A(n16019), .B(n53), .Y(n16015) );
  NOR2X1 U14588 ( .A(n73439), .B(n360), .Y(n16019) );
  NAND2X1 U14589 ( .A(n16020), .B(n16021), .Y(n16013) );
  NOR2X1 U14590 ( .A(n16022), .B(n16023), .Y(n16021) );
  NOR2X1 U14591 ( .A(n340), .B(n15829), .Y(n16023) );
  NOR2X1 U14592 ( .A(n42454), .B(n15824), .Y(n16022) );
  NOR2X1 U14593 ( .A(n16024), .B(n16025), .Y(n16020) );
  NOR2X1 U14594 ( .A(n73448), .B(n40669), .Y(n16025) );
  NOR2X1 U14595 ( .A(n73446), .B(n362), .Y(n16024) );
  NAND2X1 U14598 ( .A(n16030), .B(n16031), .Y(n16029) );
  NOR2X1 U14599 ( .A(n16032), .B(n16033), .Y(n16031) );
  NAND2X1 U14603 ( .A(n16036), .B(n16037), .Y(n15836) );
  NOR2X1 U14604 ( .A(n16038), .B(n16039), .Y(n16037) );
  NAND2X1 U14605 ( .A(n16040), .B(n16041), .Y(n16039) );
  NAND2X1 U14606 ( .A(n371), .B(n15447), .Y(n16041) );
  NAND2X1 U14607 ( .A(n368), .B(n16042), .Y(n16040) );
  NOR2X1 U14608 ( .A(n73468), .B(n42960), .Y(n16038) );
  NOR2X1 U14609 ( .A(n16043), .B(n16044), .Y(n16036) );
  NAND2X1 U14610 ( .A(n16045), .B(n16046), .Y(n16044) );
  NAND2X1 U14611 ( .A(n73511), .B(n16047), .Y(n16046) );
  NAND2X1 U14612 ( .A(n73512), .B(n16048), .Y(n16045) );
  NOR2X1 U14613 ( .A(n73444), .B(n15465), .Y(n16043) );
  NOR2X1 U14614 ( .A(n16049), .B(n16050), .Y(n16030) );
  NOR2X1 U14615 ( .A(n16051), .B(n42945), .Y(n16050) );
  NOR2X1 U14616 ( .A(n15462), .B(n15829), .Y(n16049) );
  NAND2X1 U14617 ( .A(n16052), .B(n16053), .Y(n16028) );
  NOR2X1 U14618 ( .A(n16054), .B(n16055), .Y(n16053) );
  NAND2X1 U14619 ( .A(n16056), .B(n16057), .Y(n16055) );
  NAND2X1 U14620 ( .A(n73444), .B(n16058), .Y(n16057) );
  NAND2X1 U14621 ( .A(n16059), .B(n16060), .Y(n16058) );
  NAND2X1 U14622 ( .A(n73443), .B(n16061), .Y(n16060) );
  NAND2X1 U14623 ( .A(n16062), .B(n16004), .Y(n16059) );
  NAND2X1 U14624 ( .A(n16063), .B(n16003), .Y(n16056) );
  NAND2X1 U14625 ( .A(n16064), .B(n16065), .Y(n16063) );
  NAND2X1 U14626 ( .A(n73443), .B(n16062), .Y(n16065) );
  NOR2X1 U14631 ( .A(n981), .B(n16070), .Y(n16064) );
  NOR2X1 U14632 ( .A(n73443), .B(n16071), .Y(n16070) );
  NOR2X1 U14633 ( .A(n980), .B(n16061), .Y(n16071) );
  NAND2X1 U14636 ( .A(n16074), .B(n16075), .Y(n16005) );
  NAND2X1 U14637 ( .A(n16076), .B(n16077), .Y(n16075) );
  OR2X1 U14638 ( .A(n16078), .B(n16079), .Y(n16076) );
  NAND2X1 U14639 ( .A(n16079), .B(n16078), .Y(n16074) );
  NOR2X1 U14641 ( .A(n73458), .B(n15880), .Y(n16054) );
  NOR2X1 U14642 ( .A(n16081), .B(n16082), .Y(n16052) );
  AND2X1 U14643 ( .A(n73511), .B(n37552), .Y(n16082) );
  NOR2X1 U14644 ( .A(n73456), .B(n16084), .Y(n16081) );
  NAND2X1 U14646 ( .A(n16087), .B(n16088), .Y(n16086) );
  NOR2X1 U14647 ( .A(n16089), .B(n16090), .Y(n16088) );
  NOR2X1 U14648 ( .A(n73450), .B(n40669), .Y(n16090) );
  NOR2X1 U14649 ( .A(n73448), .B(n42943), .Y(n16089) );
  NOR2X1 U14650 ( .A(n16091), .B(n53), .Y(n16087) );
  NOR2X1 U14651 ( .A(n16092), .B(n16093), .Y(n15884) );
  NOR2X1 U14652 ( .A(n15887), .B(n73433), .Y(n16093) );
  NOR2X1 U14653 ( .A(n15495), .B(n15498), .Y(n16091) );
  NAND2X1 U14654 ( .A(n16094), .B(n16095), .Y(n16085) );
  NOR2X1 U14655 ( .A(n16096), .B(n16097), .Y(n16095) );
  NOR2X1 U14656 ( .A(n16098), .B(n15965), .Y(n16097) );
  NOR2X1 U14657 ( .A(n15464), .B(n15966), .Y(n16096) );
  NOR2X1 U14658 ( .A(n16099), .B(n16100), .Y(n16094) );
  NOR2X1 U14659 ( .A(n73446), .B(n40674), .Y(n16100) );
  NOR2X1 U14660 ( .A(n16101), .B(n42960), .Y(n16099) );
  NAND2X1 U14663 ( .A(n16106), .B(n16107), .Y(n16105) );
  NOR2X1 U14664 ( .A(n16108), .B(n16109), .Y(n16107) );
  NAND2X1 U14665 ( .A(n16110), .B(n16111), .Y(n16109) );
  NAND2X1 U14666 ( .A(n42452), .B(n73511), .Y(n16111) );
  NAND2X1 U14667 ( .A(n369), .B(n16113), .Y(n16110) );
  NOR2X1 U14668 ( .A(n15828), .B(n15966), .Y(n16108) );
  NOR2X1 U14669 ( .A(n16114), .B(n16115), .Y(n16106) );
  NOR2X1 U14670 ( .A(n16116), .B(n42960), .Y(n16115) );
  NOR2X1 U14671 ( .A(n16117), .B(n42944), .Y(n16114) );
  NAND2X1 U14672 ( .A(n16118), .B(n16119), .Y(n16104) );
  NOR2X1 U14673 ( .A(n16120), .B(n16121), .Y(n16119) );
  NAND2X1 U14674 ( .A(n16122), .B(n16123), .Y(n16121) );
  NAND2X1 U14675 ( .A(n73446), .B(n16124), .Y(n16123) );
  NAND2X1 U14676 ( .A(n16125), .B(n16126), .Y(n16124) );
  NAND2X1 U14677 ( .A(n73445), .B(n16127), .Y(n16126) );
  NAND2X1 U14678 ( .A(n16128), .B(n16078), .Y(n16125) );
  NAND2X1 U14679 ( .A(n16129), .B(n16077), .Y(n16122) );
  NAND2X1 U14680 ( .A(n16130), .B(n15416), .Y(n16129) );
  NOR2X1 U14681 ( .A(n16131), .B(n16132), .Y(n16130) );
  AND2X1 U14682 ( .A(n16128), .B(n73445), .Y(n16132) );
  NOR2X1 U14687 ( .A(n73445), .B(n16137), .Y(n16131) );
  NOR2X1 U14688 ( .A(n980), .B(n16127), .Y(n16137) );
  NAND2X1 U14691 ( .A(n16140), .B(n16141), .Y(n16079) );
  NAND2X1 U14692 ( .A(n16142), .B(n16143), .Y(n16141) );
  OR2X1 U14693 ( .A(n16144), .B(n16145), .Y(n16142) );
  NAND2X1 U14694 ( .A(n16145), .B(n16144), .Y(n16140) );
  NOR2X1 U14696 ( .A(n73460), .B(n15880), .Y(n16120) );
  NOR2X1 U14697 ( .A(n16146), .B(n16147), .Y(n16118) );
  NOR2X1 U14698 ( .A(n73462), .B(n16148), .Y(n16147) );
  NOR2X1 U14699 ( .A(n73458), .B(n16084), .Y(n16146) );
  NAND2X1 U14701 ( .A(n16151), .B(n16152), .Y(n16150) );
  NOR2X1 U14702 ( .A(n16153), .B(n16154), .Y(n16152) );
  NAND2X1 U14703 ( .A(n16155), .B(n16156), .Y(n16154) );
  NAND2X1 U14704 ( .A(n15442), .B(n16047), .Y(n16156) );
  NAND2X1 U14705 ( .A(n37539), .B(n15874), .Y(n16155) );
  NOR2X1 U14706 ( .A(n73439), .B(n42985), .Y(n16153) );
  NOR2X1 U14707 ( .A(n16158), .B(n16092), .Y(n16151) );
  NOR2X1 U14708 ( .A(n73444), .B(n42991), .Y(n16158) );
  NAND2X1 U14709 ( .A(n16159), .B(n16160), .Y(n16149) );
  NOR2X1 U14710 ( .A(n16161), .B(n16162), .Y(n16160) );
  NAND2X1 U14711 ( .A(n16163), .B(n16164), .Y(n16162) );
  NAND2X1 U14712 ( .A(n368), .B(n16165), .Y(n16164) );
  OR2X1 U14713 ( .A(n43008), .B(n16166), .Y(n16163) );
  NOR2X1 U14714 ( .A(n73454), .B(n15672), .Y(n16161) );
  NOR2X1 U14715 ( .A(n16167), .B(n16168), .Y(n16159) );
  NOR2X1 U14716 ( .A(n73450), .B(n362), .Y(n16168) );
  NOR2X1 U14717 ( .A(n73448), .B(n364), .Y(n16167) );
  NAND2X1 U14720 ( .A(n16173), .B(n16174), .Y(n16172) );
  NOR2X1 U14721 ( .A(n16175), .B(n16176), .Y(n16174) );
  NAND2X1 U14722 ( .A(n16177), .B(n16178), .Y(n16176) );
  NAND2X1 U14724 ( .A(n16179), .B(n16180), .Y(n16009) );
  NAND2X1 U14725 ( .A(n42958), .B(n15846), .Y(n16180) );
  NAND2X1 U14726 ( .A(n73512), .B(n16181), .Y(n16179) );
  NAND2X1 U14727 ( .A(n369), .B(n16182), .Y(n16177) );
  NOR2X1 U14728 ( .A(n15610), .B(n15966), .Y(n16175) );
  NOR2X1 U14729 ( .A(n16183), .B(n16184), .Y(n16173) );
  NOR2X1 U14730 ( .A(n16185), .B(n15453), .Y(n16184) );
  NOR2X1 U14731 ( .A(n16186), .B(n15505), .Y(n16183) );
  NAND2X1 U14732 ( .A(n16187), .B(n16188), .Y(n16171) );
  NOR2X1 U14733 ( .A(n16189), .B(n16190), .Y(n16188) );
  NAND2X1 U14734 ( .A(n16191), .B(n16192), .Y(n16190) );
  NAND2X1 U14735 ( .A(n42312), .B(n73511), .Y(n16192) );
  NAND2X1 U14736 ( .A(n73448), .B(n16194), .Y(n16191) );
  NAND2X1 U14737 ( .A(n16195), .B(n16196), .Y(n16194) );
  NAND2X1 U14738 ( .A(n73447), .B(n16197), .Y(n16196) );
  NAND2X1 U14739 ( .A(n16198), .B(n16144), .Y(n16195) );
  NOR2X1 U14740 ( .A(n73448), .B(n16199), .Y(n16189) );
  NOR2X1 U14741 ( .A(n42972), .B(n16200), .Y(n16199) );
  NAND2X1 U14742 ( .A(n16201), .B(n16202), .Y(n16200) );
  NAND2X1 U14743 ( .A(n16203), .B(n16144), .Y(n16202) );
  OR2X1 U14744 ( .A(n16197), .B(n980), .Y(n16203) );
  NAND2X1 U14748 ( .A(n73447), .B(n16198), .Y(n16201) );
  NAND2X1 U14753 ( .A(n16210), .B(n16211), .Y(n16145) );
  NAND2X1 U14754 ( .A(n16212), .B(n16213), .Y(n16211) );
  OR2X1 U14755 ( .A(n16214), .B(n16215), .Y(n16212) );
  NAND2X1 U14756 ( .A(n16215), .B(n16214), .Y(n16210) );
  NOR2X1 U14757 ( .A(n16216), .B(n16217), .Y(n16187) );
  NOR2X1 U14758 ( .A(n73460), .B(n16084), .Y(n16217) );
  NOR2X1 U14759 ( .A(n73462), .B(n15880), .Y(n16216) );
  NAND2X1 U14761 ( .A(n16220), .B(n16221), .Y(n16219) );
  NOR2X1 U14762 ( .A(n16222), .B(n16223), .Y(n16221) );
  NAND2X1 U14763 ( .A(n16224), .B(n16225), .Y(n16223) );
  NAND2X1 U14764 ( .A(n15442), .B(n15802), .Y(n16225) );
  NAND2X1 U14765 ( .A(n37539), .B(n16003), .Y(n16224) );
  NOR2X1 U14766 ( .A(n73442), .B(n358), .Y(n16222) );
  NOR2X1 U14767 ( .A(n16226), .B(n16092), .Y(n16220) );
  NOR2X1 U14768 ( .A(n73446), .B(n42990), .Y(n16226) );
  NAND2X1 U14769 ( .A(n16227), .B(n16228), .Y(n16218) );
  NOR2X1 U14770 ( .A(n16229), .B(n16230), .Y(n16228) );
  NAND2X1 U14771 ( .A(n16231), .B(n16232), .Y(n16230) );
  NAND2X1 U14772 ( .A(n368), .B(n16233), .Y(n16232) );
  NAND2X1 U14773 ( .A(n42958), .B(n16234), .Y(n16231) );
  NOR2X1 U14774 ( .A(n73456), .B(n15672), .Y(n16229) );
  NOR2X1 U14775 ( .A(n16235), .B(n16236), .Y(n16227) );
  NOR2X1 U14776 ( .A(n73452), .B(n42943), .Y(n16236) );
  NOR2X1 U14777 ( .A(n73450), .B(n364), .Y(n16235) );
  NAND2X1 U14780 ( .A(n16242), .B(n16243), .Y(n16241) );
  NOR2X1 U14781 ( .A(n16244), .B(n16245), .Y(n16243) );
  NAND2X1 U14782 ( .A(n16246), .B(n16247), .Y(n16245) );
  OR2X1 U14783 ( .A(n16148), .B(n73466), .Y(n16247) );
  NAND2X1 U14784 ( .A(n42958), .B(n16248), .Y(n16246) );
  NOR2X1 U14785 ( .A(n42454), .B(n15829), .Y(n16244) );
  NOR2X1 U14786 ( .A(n16249), .B(n16250), .Y(n16242) );
  NOR2X1 U14787 ( .A(n16251), .B(n42945), .Y(n16250) );
  NOR2X1 U14788 ( .A(n340), .B(n15966), .Y(n16249) );
  NAND2X1 U14789 ( .A(n16252), .B(n16253), .Y(n16240) );
  NOR2X1 U14790 ( .A(n16254), .B(n16255), .Y(n16253) );
  NAND2X1 U14791 ( .A(n16256), .B(n16257), .Y(n16255) );
  NAND2X1 U14792 ( .A(n42314), .B(n73511), .Y(n16257) );
  NAND2X1 U14793 ( .A(n73450), .B(n16259), .Y(n16256) );
  NAND2X1 U14794 ( .A(n16260), .B(n16261), .Y(n16259) );
  NAND2X1 U14795 ( .A(n73449), .B(n16262), .Y(n16261) );
  NAND2X1 U14796 ( .A(n16263), .B(n16214), .Y(n16260) );
  NOR2X1 U14797 ( .A(n73450), .B(n16264), .Y(n16254) );
  NOR2X1 U14798 ( .A(n361), .B(n16265), .Y(n16264) );
  NAND2X1 U14799 ( .A(n16266), .B(n16267), .Y(n16265) );
  NAND2X1 U14800 ( .A(n16268), .B(n16214), .Y(n16267) );
  OR2X1 U14801 ( .A(n16262), .B(n980), .Y(n16268) );
  NAND2X1 U14805 ( .A(n73449), .B(n16263), .Y(n16266) );
  NAND2X1 U14810 ( .A(n16275), .B(n16276), .Y(n16215) );
  NAND2X1 U14811 ( .A(n16277), .B(n16047), .Y(n16276) );
  OR2X1 U14812 ( .A(n16278), .B(n16279), .Y(n16277) );
  NAND2X1 U14813 ( .A(n16279), .B(n16278), .Y(n16275) );
  NOR2X1 U14814 ( .A(n16280), .B(n16281), .Y(n16252) );
  NOR2X1 U14815 ( .A(n73462), .B(n16084), .Y(n16281) );
  NOR2X1 U14817 ( .A(n73464), .B(n15880), .Y(n16280) );
  NAND2X1 U14820 ( .A(n16284), .B(n16285), .Y(n16283) );
  NOR2X1 U14821 ( .A(n16286), .B(n16287), .Y(n16285) );
  NAND2X1 U14822 ( .A(n16288), .B(n16289), .Y(n16287) );
  NAND2X1 U14823 ( .A(n15442), .B(n16290), .Y(n16289) );
  NAND2X1 U14824 ( .A(n37539), .B(n16077), .Y(n16288) );
  NOR2X1 U14825 ( .A(n73444), .B(n42984), .Y(n16286) );
  NOR2X1 U14826 ( .A(n16291), .B(n16092), .Y(n16284) );
  NOR2X1 U14827 ( .A(n73448), .B(n42990), .Y(n16291) );
  NAND2X1 U14828 ( .A(n16292), .B(n16293), .Y(n16282) );
  NOR2X1 U14829 ( .A(n16294), .B(n16295), .Y(n16293) );
  NAND2X1 U14830 ( .A(n16296), .B(n16297), .Y(n16295) );
  NAND2X1 U14831 ( .A(n368), .B(n16298), .Y(n16297) );
  NAND2X1 U14832 ( .A(n73570), .B(n16299), .Y(n16296) );
  NOR2X1 U14833 ( .A(n73458), .B(n15672), .Y(n16294) );
  NOR2X1 U14834 ( .A(n16300), .B(n16301), .Y(n16292) );
  NOR2X1 U14835 ( .A(n73454), .B(n362), .Y(n16301) );
  NOR2X1 U14836 ( .A(n73452), .B(n364), .Y(n16300) );
  NAND2X1 U14839 ( .A(n16306), .B(n16307), .Y(n16305) );
  NOR2X1 U14840 ( .A(n16308), .B(n16309), .Y(n16307) );
  NOR2X1 U14841 ( .A(n15462), .B(n15966), .Y(n16309) );
  NOR2X1 U14842 ( .A(n16051), .B(n42946), .Y(n16308) );
  NOR2X1 U14843 ( .A(n16310), .B(n16311), .Y(n16306) );
  NOR2X1 U14844 ( .A(n16101), .B(n42944), .Y(n16311) );
  NOR2X1 U14845 ( .A(n16312), .B(n15965), .Y(n16310) );
  NAND2X1 U14846 ( .A(n16313), .B(n16314), .Y(n16304) );
  NOR2X1 U14847 ( .A(n16315), .B(n16316), .Y(n16314) );
  NAND2X1 U14848 ( .A(n16317), .B(n16318), .Y(n16316) );
  NAND2X1 U14849 ( .A(n73452), .B(n16319), .Y(n16318) );
  NAND2X1 U14850 ( .A(n16320), .B(n16321), .Y(n16319) );
  NAND2X1 U14851 ( .A(n73451), .B(n16322), .Y(n16321) );
  NAND2X1 U14852 ( .A(n16323), .B(n16278), .Y(n16320) );
  NAND2X1 U14853 ( .A(n16324), .B(n16047), .Y(n16317) );
  NAND2X1 U14854 ( .A(n16325), .B(n15416), .Y(n16324) );
  NOR2X1 U14855 ( .A(n16326), .B(n16327), .Y(n16325) );
  AND2X1 U14856 ( .A(n16323), .B(n73451), .Y(n16327) );
  NOR2X1 U14861 ( .A(n73451), .B(n16332), .Y(n16326) );
  NOR2X1 U14862 ( .A(n980), .B(n16322), .Y(n16332) );
  NAND2X1 U14865 ( .A(n16335), .B(n16336), .Y(n16279) );
  NAND2X1 U14866 ( .A(n16337), .B(n15802), .Y(n16336) );
  OR2X1 U14867 ( .A(n16338), .B(n16339), .Y(n16337) );
  NAND2X1 U14868 ( .A(n16339), .B(n16338), .Y(n16335) );
  NOR2X1 U14870 ( .A(n73468), .B(n16148), .Y(n16315) );
  NOR2X1 U14871 ( .A(n16340), .B(n16341), .Y(n16313) );
  NOR2X1 U14874 ( .A(n16343), .B(n42959), .Y(n16340) );
  NAND2X1 U14876 ( .A(n16346), .B(n16347), .Y(n16345) );
  NOR2X1 U14877 ( .A(n16348), .B(n16349), .Y(n16347) );
  NOR2X1 U14878 ( .A(n15495), .B(n43008), .Y(n16349) );
  NOR2X1 U14879 ( .A(n73446), .B(n42985), .Y(n16348) );
  NOR2X1 U14880 ( .A(n16350), .B(n16092), .Y(n16346) );
  NAND2X1 U14881 ( .A(n16351), .B(n16352), .Y(n16092) );
  NAND2X1 U14882 ( .A(n73524), .B(n54), .Y(n16352) );
  NOR2X1 U14883 ( .A(n73450), .B(n42991), .Y(n16350) );
  NAND2X1 U14884 ( .A(n16353), .B(n16354), .Y(n16344) );
  NOR2X1 U14885 ( .A(n16355), .B(n16356), .Y(n16354) );
  NAND2X1 U14886 ( .A(n16357), .B(n16358), .Y(n16356) );
  NAND2X1 U14887 ( .A(n73395), .B(n16048), .Y(n16358) );
  NAND2X1 U14888 ( .A(n73510), .B(n15802), .Y(n16357) );
  NOR2X1 U14889 ( .A(n73456), .B(n42943), .Y(n16355) );
  NOR2X1 U14890 ( .A(n16359), .B(n16360), .Y(n16353) );
  NOR2X1 U14891 ( .A(n73448), .B(n42988), .Y(n16360) );
  NOR2X1 U14892 ( .A(n73458), .B(n363), .Y(n16359) );
  NAND2X1 U14895 ( .A(n16365), .B(n16366), .Y(n16364) );
  NOR2X1 U14896 ( .A(n16367), .B(n16368), .Y(n16366) );
  NOR2X1 U14897 ( .A(n300), .B(n42960), .Y(n16368) );
  NOR2X1 U14898 ( .A(n15828), .B(n15965), .Y(n16367) );
  NOR2X1 U14899 ( .A(n16369), .B(n16370), .Y(n16365) );
  NOR2X1 U14900 ( .A(n73462), .B(n15672), .Y(n16370) );
  NOR2X1 U14901 ( .A(n16166), .B(n43010), .Y(n16369) );
  NAND2X1 U14902 ( .A(n16371), .B(n16372), .Y(n16363) );
  NOR2X1 U14903 ( .A(n16373), .B(n16374), .Y(n16372) );
  NAND2X1 U14904 ( .A(n16375), .B(n16376), .Y(n16374) );
  NAND2X1 U14905 ( .A(n73454), .B(n16377), .Y(n16376) );
  NAND2X1 U14906 ( .A(n16378), .B(n16379), .Y(n16377) );
  NAND2X1 U14907 ( .A(n73453), .B(n16380), .Y(n16379) );
  NAND2X1 U14908 ( .A(n16381), .B(n16338), .Y(n16378) );
  NAND2X1 U14909 ( .A(n16382), .B(n15802), .Y(n16375) );
  NAND2X1 U14910 ( .A(n16383), .B(n15416), .Y(n16382) );
  NOR2X1 U14911 ( .A(n16384), .B(n16385), .Y(n16383) );
  AND2X1 U14912 ( .A(n16381), .B(n73453), .Y(n16385) );
  NOR2X1 U14917 ( .A(n73453), .B(n16390), .Y(n16384) );
  NOR2X1 U14918 ( .A(n980), .B(n16380), .Y(n16390) );
  NAND2X1 U14921 ( .A(n16393), .B(n16394), .Y(n16339) );
  NAND2X1 U14922 ( .A(n16395), .B(n16290), .Y(n16394) );
  OR2X1 U14923 ( .A(n16396), .B(n16397), .Y(n16395) );
  NAND2X1 U14924 ( .A(n16397), .B(n16396), .Y(n16393) );
  NOR2X1 U14926 ( .A(n378), .B(n15966), .Y(n16373) );
  NOR2X1 U14927 ( .A(n16398), .B(n16399), .Y(n16371) );
  NOR2X1 U14928 ( .A(n16116), .B(n15453), .Y(n16399) );
  NOR2X1 U14929 ( .A(n16117), .B(n15463), .Y(n16398) );
  NAND2X1 U14931 ( .A(n16402), .B(n16403), .Y(n16401) );
  NOR2X1 U14932 ( .A(n16404), .B(n16405), .Y(n16403) );
  NOR2X1 U14933 ( .A(n73448), .B(n358), .Y(n16405) );
  NOR2X1 U14934 ( .A(n73450), .B(n42987), .Y(n16404) );
  NOR2X1 U14935 ( .A(n16406), .B(n16407), .Y(n16402) );
  NOR2X1 U14936 ( .A(n73452), .B(n42990), .Y(n16406) );
  NAND2X1 U14937 ( .A(n16408), .B(n16409), .Y(n16400) );
  NOR2X1 U14938 ( .A(n16410), .B(n16411), .Y(n16409) );
  NOR2X1 U14939 ( .A(n73456), .B(n40674), .Y(n16411) );
  NOR2X1 U14940 ( .A(n15556), .B(n15505), .Y(n16410) );
  NOR2X1 U14941 ( .A(n16412), .B(n16413), .Y(n16408) );
  NOR2X1 U14942 ( .A(n73460), .B(n40669), .Y(n16413) );
  NOR2X1 U14943 ( .A(n73458), .B(n42943), .Y(n16412) );
  NAND2X1 U14946 ( .A(n16418), .B(n16419), .Y(n16417) );
  NOR2X1 U14947 ( .A(n16420), .B(n16421), .Y(n16419) );
  NOR2X1 U14948 ( .A(n15610), .B(n15965), .Y(n16421) );
  NOR2X1 U14949 ( .A(n16185), .B(n42946), .Y(n16420) );
  NOR2X1 U14950 ( .A(n16422), .B(n16423), .Y(n16418) );
  NOR2X1 U14951 ( .A(n309), .B(n42945), .Y(n16423) );
  NOR2X1 U14952 ( .A(n180), .B(n15847), .Y(n16422) );
  NAND2X1 U14953 ( .A(n16424), .B(n16425), .Y(n16416) );
  NOR2X1 U14954 ( .A(n16426), .B(n16427), .Y(n16425) );
  NAND2X1 U14955 ( .A(n16428), .B(n16429), .Y(n16427) );
  NAND2X1 U14956 ( .A(n73456), .B(n16430), .Y(n16429) );
  NAND2X1 U14957 ( .A(n16431), .B(n16432), .Y(n16430) );
  NAND2X1 U14958 ( .A(n73455), .B(n16433), .Y(n16432) );
  NAND2X1 U14959 ( .A(n16434), .B(n16396), .Y(n16431) );
  NAND2X1 U14960 ( .A(n16435), .B(n16290), .Y(n16428) );
  NAND2X1 U14961 ( .A(n16436), .B(n15416), .Y(n16435) );
  NOR2X1 U14962 ( .A(n16437), .B(n16438), .Y(n16436) );
  AND2X1 U14963 ( .A(n16434), .B(n73455), .Y(n16438) );
  NOR2X1 U14968 ( .A(n73455), .B(n16443), .Y(n16437) );
  NOR2X1 U14969 ( .A(n980), .B(n16433), .Y(n16443) );
  NAND2X1 U14972 ( .A(n16446), .B(n16447), .Y(n16397) );
  NAND2X1 U14973 ( .A(n16448), .B(n16449), .Y(n16447) );
  OR2X1 U14974 ( .A(n16450), .B(n16451), .Y(n16448) );
  NAND2X1 U14975 ( .A(n16451), .B(n16450), .Y(n16446) );
  NOR2X1 U14977 ( .A(n73472), .B(n16148), .Y(n16426) );
  NOR2X1 U14979 ( .A(n16452), .B(n16453), .Y(n16424) );
  NOR2X1 U14980 ( .A(n16186), .B(n43011), .Y(n16453) );
  NOR2X1 U14981 ( .A(n73397), .B(n15966), .Y(n16452) );
  NAND2X1 U14983 ( .A(n16456), .B(n16457), .Y(n16455) );
  NOR2X1 U14984 ( .A(n16458), .B(n16459), .Y(n16457) );
  NOR2X1 U14985 ( .A(n73450), .B(n42984), .Y(n16459) );
  NOR2X1 U14986 ( .A(n73452), .B(n42988), .Y(n16458) );
  NOR2X1 U14987 ( .A(n16460), .B(n16407), .Y(n16456) );
  NOR2X1 U14988 ( .A(n73454), .B(n42991), .Y(n16460) );
  NAND2X1 U14989 ( .A(n16461), .B(n16462), .Y(n16454) );
  NOR2X1 U14990 ( .A(n16463), .B(n16464), .Y(n16462) );
  NAND2X1 U14991 ( .A(n16465), .B(n16466), .Y(n16464) );
  NAND2X1 U14992 ( .A(n73395), .B(n16181), .Y(n16466) );
  NAND2X1 U14993 ( .A(n73510), .B(n16449), .Y(n16465) );
  NOR2X1 U14994 ( .A(n73460), .B(n42943), .Y(n16463) );
  NOR2X1 U14995 ( .A(n16467), .B(n16468), .Y(n16461) );
  NOR2X1 U14996 ( .A(n15607), .B(n43008), .Y(n16468) );
  NOR2X1 U14997 ( .A(n73462), .B(n363), .Y(n16467) );
  NAND2X1 U15000 ( .A(n16473), .B(n16474), .Y(n16472) );
  NOR2X1 U15001 ( .A(n16475), .B(n16476), .Y(n16474) );
  NOR2X1 U15002 ( .A(n257), .B(n15505), .Y(n16476) );
  NOR2X1 U15003 ( .A(n340), .B(n15965), .Y(n16475) );
  NOR2X1 U15004 ( .A(n16477), .B(n16478), .Y(n16473) );
  NOR2X1 U15005 ( .A(n179), .B(n42960), .Y(n16478) );
  NOR2X1 U15006 ( .A(n55), .B(n43010), .Y(n16477) );
  NAND2X1 U15007 ( .A(n16479), .B(n16480), .Y(n16471) );
  NOR2X1 U15008 ( .A(n16481), .B(n16482), .Y(n16480) );
  NAND2X1 U15009 ( .A(n16483), .B(n16484), .Y(n16482) );
  NAND2X1 U15010 ( .A(n73458), .B(n16485), .Y(n16484) );
  NAND2X1 U15011 ( .A(n16486), .B(n16487), .Y(n16485) );
  NAND2X1 U15012 ( .A(n73457), .B(n16488), .Y(n16487) );
  NAND2X1 U15013 ( .A(n16489), .B(n16450), .Y(n16486) );
  NAND2X1 U15014 ( .A(n16490), .B(n16449), .Y(n16483) );
  NAND2X1 U15015 ( .A(n16491), .B(n15416), .Y(n16490) );
  NOR2X1 U15016 ( .A(n16492), .B(n16493), .Y(n16491) );
  AND2X1 U15017 ( .A(n16489), .B(n73457), .Y(n16493) );
  NOR2X1 U15022 ( .A(n73457), .B(n16498), .Y(n16492) );
  NOR2X1 U15023 ( .A(n980), .B(n16488), .Y(n16498) );
  NAND2X1 U15026 ( .A(n16501), .B(n16502), .Y(n16451) );
  NAND2X1 U15027 ( .A(n16503), .B(n16048), .Y(n16502) );
  OR2X1 U15028 ( .A(n16504), .B(n16505), .Y(n16503) );
  NAND2X1 U15029 ( .A(n16505), .B(n16504), .Y(n16501) );
  AND2X1 U15031 ( .A(n16248), .B(n73512), .Y(n16481) );
  NAND2X1 U15032 ( .A(n16506), .B(n16507), .Y(n16248) );
  NOR2X1 U15033 ( .A(n16508), .B(n16509), .Y(n16479) );
  NOR2X1 U15034 ( .A(n16251), .B(n15463), .Y(n16509) );
  NOR2X1 U15035 ( .A(n42454), .B(n15966), .Y(n16508) );
  NAND2X1 U15037 ( .A(n16512), .B(n16513), .Y(n16511) );
  NOR2X1 U15038 ( .A(n16514), .B(n16515), .Y(n16513) );
  NOR2X1 U15039 ( .A(n73452), .B(n42985), .Y(n16515) );
  NOR2X1 U15040 ( .A(n73454), .B(n42987), .Y(n16514) );
  NOR2X1 U15041 ( .A(n16516), .B(n16407), .Y(n16512) );
  NOR2X1 U15042 ( .A(n73456), .B(n42991), .Y(n16516) );
  NAND2X1 U15043 ( .A(n16517), .B(n16518), .Y(n16510) );
  NOR2X1 U15044 ( .A(n16519), .B(n16520), .Y(n16518) );
  NOR2X1 U15045 ( .A(n73460), .B(n40674), .Y(n16520) );
  NOR2X1 U15046 ( .A(n73466), .B(n15672), .Y(n16519) );
  NOR2X1 U15047 ( .A(n16521), .B(n16522), .Y(n16517) );
  NOR2X1 U15048 ( .A(n73464), .B(n40669), .Y(n16522) );
  NOR2X1 U15049 ( .A(n73462), .B(n362), .Y(n16521) );
  NAND2X1 U15052 ( .A(n16527), .B(n16528), .Y(n16526) );
  NOR2X1 U15053 ( .A(n16529), .B(n16530), .Y(n16528) );
  NOR2X1 U15054 ( .A(n15462), .B(n15965), .Y(n16530) );
  NOR2X1 U15057 ( .A(n16532), .B(n16533), .Y(n16527) );
  NOR2X1 U15058 ( .A(n16101), .B(n42946), .Y(n16533) );
  NOR2X1 U15059 ( .A(n16312), .B(n15847), .Y(n16532) );
  NAND2X1 U15060 ( .A(n16534), .B(n16535), .Y(n16525) );
  NOR2X1 U15061 ( .A(n16536), .B(n16537), .Y(n16535) );
  NOR2X1 U15062 ( .A(n73460), .B(n16538), .Y(n16537) );
  NOR2X1 U15063 ( .A(n42971), .B(n16539), .Y(n16538) );
  NAND2X1 U15064 ( .A(n16540), .B(n16541), .Y(n16539) );
  NAND2X1 U15065 ( .A(n16542), .B(n16504), .Y(n16541) );
  NAND2X1 U15066 ( .A(n42197), .B(n42970), .Y(n16542) );
  NAND2X1 U15067 ( .A(n73459), .B(n16544), .Y(n16540) );
  NOR2X1 U15068 ( .A(n16545), .B(n16048), .Y(n16536) );
  NOR2X1 U15069 ( .A(n16546), .B(n16547), .Y(n16545) );
  AND2X1 U15070 ( .A(n16504), .B(n16544), .Y(n16547) );
  NOR2X1 U15075 ( .A(n42197), .B(n16504), .Y(n16546) );
  NAND2X1 U15078 ( .A(n16554), .B(n16555), .Y(n16505) );
  NAND2X1 U15079 ( .A(n16556), .B(n15801), .Y(n16555) );
  OR2X1 U15080 ( .A(n16557), .B(n16558), .Y(n16556) );
  NAND2X1 U15081 ( .A(n16558), .B(n16557), .Y(n16554) );
  NOR2X1 U15083 ( .A(n16559), .B(n16560), .Y(n16534) );
  NOR2X1 U15084 ( .A(n16051), .B(n40684), .Y(n16560) );
  AND2X1 U15085 ( .A(n16561), .B(n16562), .Y(n16051) );
  NOR2X1 U15087 ( .A(n42313), .B(n42320), .Y(n16561) );
  NOR2X1 U15088 ( .A(n16343), .B(n42944), .Y(n16559) );
  AND2X1 U15089 ( .A(n16098), .B(n16566), .Y(n16343) );
  NAND2X1 U15091 ( .A(n16569), .B(n52), .Y(n16568) );
  NAND2X1 U15092 ( .A(n16351), .B(n16570), .Y(n16407) );
  NAND2X1 U15093 ( .A(n16571), .B(n54), .Y(n16570) );
  NOR2X1 U15094 ( .A(n73525), .B(n73433), .Y(n16571) );
  NOR2X1 U15095 ( .A(n16572), .B(n16573), .Y(n16569) );
  NOR2X1 U15096 ( .A(n73458), .B(n42990), .Y(n16573) );
  NOR2X1 U15097 ( .A(n15492), .B(n43008), .Y(n16572) );
  NAND2X1 U15098 ( .A(n16574), .B(n16575), .Y(n16567) );
  NOR2X1 U15099 ( .A(n16576), .B(n16577), .Y(n16575) );
  NOR2X1 U15100 ( .A(n73456), .B(n42988), .Y(n16577) );
  NOR2X1 U15101 ( .A(n73468), .B(n15672), .Y(n16576) );
  NOR2X1 U15102 ( .A(n16578), .B(n16579), .Y(n16574) );
  NOR2X1 U15103 ( .A(n15495), .B(n43011), .Y(n16579) );
  NOR2X1 U15104 ( .A(n73454), .B(n358), .Y(n16578) );
  NAND2X1 U15107 ( .A(n16584), .B(n16585), .Y(n16583) );
  OR2X1 U15108 ( .A(n15649), .B(n73488), .Y(n16585) );
  NOR2X1 U15109 ( .A(n16586), .B(n16587), .Y(n16584) );
  NOR2X1 U15110 ( .A(n73486), .B(n15722), .Y(n16587) );
  NOR2X1 U15111 ( .A(n73484), .B(n15723), .Y(n16586) );
  NAND2X1 U15113 ( .A(n16588), .B(n16589), .Y(n16582) );
  NOR2X1 U15114 ( .A(n16590), .B(n16591), .Y(n16589) );
  NOR2X1 U15115 ( .A(n16592), .B(n16593), .Y(n16591) );
  NOR2X1 U15116 ( .A(n16594), .B(n16595), .Y(n16592) );
  AND2X1 U15117 ( .A(n16596), .B(n16597), .Y(n16595) );
  NOR2X1 U15118 ( .A(n16598), .B(n16596), .Y(n16594) );
  NOR2X1 U15120 ( .A(n16600), .B(n16601), .Y(n16599) );
  NOR2X1 U15121 ( .A(n73492), .B(n15498), .Y(n16601) );
  NOR2X1 U15122 ( .A(n73482), .B(n43010), .Y(n16600) );
  NOR2X1 U15123 ( .A(n16602), .B(n16603), .Y(n16588) );
  NOR2X1 U15124 ( .A(n73494), .B(n15747), .Y(n16603) );
  NOR2X1 U15125 ( .A(n73523), .B(n16604), .Y(n16602) );
  NOR2X1 U15126 ( .A(n37560), .B(n16605), .Y(n16604) );
  NAND2X1 U15127 ( .A(n16606), .B(n16607), .Y(n16605) );
  NAND2X1 U15128 ( .A(n16608), .B(n16596), .Y(n16607) );
  NAND2X1 U15129 ( .A(n16598), .B(n42969), .Y(n16608) );
  NAND2X1 U15133 ( .A(n73492), .B(n16597), .Y(n16606) );
  NAND2X1 U15140 ( .A(n16618), .B(n16619), .Y(n16617) );
  NAND2X1 U15141 ( .A(n42989), .B(n15919), .Y(n16619) );
  NOR2X1 U15142 ( .A(n16621), .B(n16622), .Y(n16618) );
  NOR2X1 U15143 ( .A(n73490), .B(n42984), .Y(n16622) );
  NOR2X1 U15144 ( .A(n73495), .B(n42987), .Y(n16621) );
  NAND2X1 U15145 ( .A(n16623), .B(n16624), .Y(n16616) );
  NOR2X1 U15146 ( .A(n16625), .B(n16626), .Y(n16624) );
  NOR2X1 U15147 ( .A(n15407), .B(n15496), .Y(n16626) );
  NOR2X1 U15148 ( .A(n15409), .B(n15594), .Y(n16625) );
  AND2X1 U15149 ( .A(n16627), .B(n16628), .Y(n15409) );
  NOR2X1 U15150 ( .A(n16629), .B(n16630), .Y(n16628) );
  NOR2X1 U15151 ( .A(n55), .B(n15737), .Y(n16630) );
  NOR2X1 U15152 ( .A(n15648), .B(n16631), .Y(n16629) );
  AND2X1 U15153 ( .A(n16632), .B(n16507), .Y(n15648) );
  NOR2X1 U15155 ( .A(n16633), .B(n16634), .Y(n16627) );
  NOR2X1 U15156 ( .A(n15619), .B(n16635), .Y(n16634) );
  AND2X1 U15157 ( .A(n16636), .B(n16637), .Y(n15619) );
  NOR2X1 U15159 ( .A(n42448), .B(n42456), .Y(n16636) );
  AND2X1 U15160 ( .A(n16640), .B(n16342), .Y(n16633) );
  NOR2X1 U15161 ( .A(n16641), .B(n16642), .Y(n16623) );
  NOR2X1 U15162 ( .A(n15450), .B(n15491), .Y(n16642) );
  NOR2X1 U15163 ( .A(n42454), .B(n15465), .Y(n16641) );
  NAND2X1 U15166 ( .A(n16647), .B(n16648), .Y(n16646) );
  NAND2X1 U15167 ( .A(n73512), .B(n16165), .Y(n16648) );
  NOR2X1 U15168 ( .A(n16649), .B(n16650), .Y(n16647) );
  NOR2X1 U15169 ( .A(n378), .B(n15965), .Y(n16650) );
  NOR2X1 U15170 ( .A(n16116), .B(n15463), .Y(n16649) );
  AND2X1 U15171 ( .A(n16651), .B(n16652), .Y(n16116) );
  NOR2X1 U15172 ( .A(n16653), .B(n42324), .Y(n16652) );
  NOR2X1 U15174 ( .A(n42311), .B(n16656), .Y(n16651) );
  NAND2X1 U15176 ( .A(n16657), .B(n16658), .Y(n16645) );
  NOR2X1 U15177 ( .A(n51), .B(n16659), .Y(n16658) );
  NOR2X1 U15178 ( .A(n16660), .B(n15801), .Y(n16659) );
  NOR2X1 U15179 ( .A(n16661), .B(n16662), .Y(n16660) );
  AND2X1 U15180 ( .A(n16557), .B(n16663), .Y(n16662) );
  NOR2X1 U15181 ( .A(n42198), .B(n16557), .Y(n16661) );
  NOR2X1 U15182 ( .A(n16665), .B(n16666), .Y(n16657) );
  NOR2X1 U15183 ( .A(n16117), .B(n40684), .Y(n16666) );
  AND2X1 U15184 ( .A(n16667), .B(n16668), .Y(n16117) );
  NOR2X1 U15185 ( .A(n16669), .B(n42317), .Y(n16667) );
  NOR2X1 U15187 ( .A(n73462), .B(n16671), .Y(n16665) );
  NOR2X1 U15188 ( .A(n42972), .B(n16672), .Y(n16671) );
  NAND2X1 U15189 ( .A(n16673), .B(n16674), .Y(n16672) );
  NAND2X1 U15190 ( .A(n16675), .B(n16557), .Y(n16674) );
  NAND2X1 U15191 ( .A(n42198), .B(n42970), .Y(n16675) );
  NAND2X1 U15195 ( .A(n73461), .B(n16663), .Y(n16673) );
  NAND2X1 U15200 ( .A(n16682), .B(n16683), .Y(n16558) );
  NAND2X1 U15201 ( .A(n16684), .B(n16181), .Y(n16683) );
  OR2X1 U15202 ( .A(n16685), .B(n16686), .Y(n16684) );
  NAND2X1 U15203 ( .A(n16686), .B(n16685), .Y(n16682) );
  NAND2X1 U15205 ( .A(n16689), .B(n16690), .Y(n16688) );
  NAND2X1 U15206 ( .A(n42989), .B(n16048), .Y(n16690) );
  NOR2X1 U15207 ( .A(n16691), .B(n16692), .Y(n16689) );
  NOR2X1 U15208 ( .A(n73456), .B(n42985), .Y(n16692) );
  NOR2X1 U15209 ( .A(n73458), .B(n42988), .Y(n16691) );
  NAND2X1 U15210 ( .A(n16693), .B(n16694), .Y(n16687) );
  NOR2X1 U15211 ( .A(n16695), .B(n16696), .Y(n16694) );
  NOR2X1 U15212 ( .A(n15828), .B(n42960), .Y(n16696) );
  NOR2X1 U15213 ( .A(n16166), .B(n43007), .Y(n16695) );
  NOR2X1 U15214 ( .A(n16697), .B(n16698), .Y(n16693) );
  NOR2X1 U15215 ( .A(n15556), .B(n43011), .Y(n16698) );
  NOR2X1 U15216 ( .A(n256), .B(n15505), .Y(n16697) );
  NAND2X1 U15219 ( .A(n16703), .B(n16704), .Y(n16702) );
  NOR2X1 U15220 ( .A(n16705), .B(n16706), .Y(n16704) );
  NOR2X1 U15221 ( .A(n73397), .B(n15965), .Y(n16706) );
  NOR2X1 U15222 ( .A(n16185), .B(n40684), .Y(n16705) );
  AND2X1 U15223 ( .A(n16707), .B(n16708), .Y(n16185) );
  NOR2X1 U15225 ( .A(n16709), .B(n16710), .Y(n16707) );
  NOR2X1 U15228 ( .A(n16711), .B(n16712), .Y(n16703) );
  NOR2X1 U15229 ( .A(n309), .B(n42946), .Y(n16712) );
  NOR2X1 U15230 ( .A(n180), .B(n15453), .Y(n16711) );
  NAND2X1 U15231 ( .A(n16713), .B(n16714), .Y(n16701) );
  NOR2X1 U15232 ( .A(n51), .B(n16715), .Y(n16714) );
  NOR2X1 U15233 ( .A(n16716), .B(n16181), .Y(n16715) );
  NOR2X1 U15234 ( .A(n16717), .B(n16718), .Y(n16716) );
  AND2X1 U15235 ( .A(n16685), .B(n16719), .Y(n16718) );
  NOR2X1 U15236 ( .A(n42199), .B(n16685), .Y(n16717) );
  NOR2X1 U15237 ( .A(n16721), .B(n16722), .Y(n16713) );
  NOR2X1 U15238 ( .A(n16186), .B(n15408), .Y(n16722) );
  AND2X1 U15239 ( .A(n16723), .B(n16724), .Y(n16186) );
  NAND2X1 U15240 ( .A(n54), .B(n16593), .Y(n16724) );
  NOR2X1 U15241 ( .A(n73464), .B(n16725), .Y(n16721) );
  NOR2X1 U15242 ( .A(n361), .B(n16726), .Y(n16725) );
  NAND2X1 U15243 ( .A(n16727), .B(n16728), .Y(n16726) );
  NAND2X1 U15244 ( .A(n16729), .B(n16685), .Y(n16728) );
  NAND2X1 U15245 ( .A(n42199), .B(n42969), .Y(n16729) );
  NAND2X1 U15249 ( .A(n73463), .B(n16719), .Y(n16727) );
  NAND2X1 U15254 ( .A(n16736), .B(n16737), .Y(n16686) );
  NAND2X1 U15255 ( .A(n16738), .B(n16563), .Y(n16737) );
  OR2X1 U15256 ( .A(n16739), .B(n16740), .Y(n16738) );
  NAND2X1 U15257 ( .A(n16740), .B(n16739), .Y(n16736) );
  NAND2X1 U15259 ( .A(n16743), .B(n16744), .Y(n16742) );
  NAND2X1 U15260 ( .A(n42989), .B(n15801), .Y(n16744) );
  NOR2X1 U15261 ( .A(n16745), .B(n16746), .Y(n16743) );
  NOR2X1 U15262 ( .A(n73458), .B(n358), .Y(n16746) );
  NOR2X1 U15263 ( .A(n73460), .B(n42987), .Y(n16745) );
  NAND2X1 U15264 ( .A(n16747), .B(n16748), .Y(n16741) );
  NOR2X1 U15265 ( .A(n16749), .B(n16750), .Y(n16748) );
  NOR2X1 U15266 ( .A(n15610), .B(n15847), .Y(n16750) );
  NOR2X1 U15267 ( .A(n73472), .B(n15672), .Y(n16749) );
  NOR2X1 U15268 ( .A(n16751), .B(n16752), .Y(n16747) );
  NOR2X1 U15269 ( .A(n255), .B(n43008), .Y(n16752) );
  NOR2X1 U15270 ( .A(n15607), .B(n43010), .Y(n16751) );
  NAND2X1 U15273 ( .A(n16757), .B(n16758), .Y(n16756) );
  NOR2X1 U15274 ( .A(n16759), .B(n16760), .Y(n16758) );
  NOR2X1 U15275 ( .A(n257), .B(n43011), .Y(n16760) );
  NOR2X1 U15276 ( .A(n42454), .B(n15965), .Y(n16759) );
  NOR2X1 U15277 ( .A(n16761), .B(n16762), .Y(n16757) );
  NOR2X1 U15278 ( .A(n55), .B(n43007), .Y(n16762) );
  NOR2X1 U15279 ( .A(n15407), .B(n15505), .Y(n16761) );
  NAND2X1 U15280 ( .A(n16763), .B(n16764), .Y(n16755) );
  NOR2X1 U15281 ( .A(n51), .B(n16765), .Y(n16764) );
  NOR2X1 U15282 ( .A(n16766), .B(n16563), .Y(n16765) );
  NOR2X1 U15283 ( .A(n16767), .B(n16768), .Y(n16766) );
  AND2X1 U15284 ( .A(n16739), .B(n16769), .Y(n16768) );
  NOR2X1 U15285 ( .A(n42201), .B(n16739), .Y(n16767) );
  NOR2X1 U15286 ( .A(n16771), .B(n16772), .Y(n16763) );
  NOR2X1 U15287 ( .A(n16251), .B(n40684), .Y(n16772) );
  AND2X1 U15288 ( .A(n16773), .B(n16774), .Y(n16251) );
  NOR2X1 U15290 ( .A(n16776), .B(n42319), .Y(n16773) );
  NOR2X1 U15292 ( .A(n73466), .B(n16778), .Y(n16771) );
  NOR2X1 U15293 ( .A(n42971), .B(n16779), .Y(n16778) );
  NAND2X1 U15294 ( .A(n16780), .B(n16781), .Y(n16779) );
  NAND2X1 U15295 ( .A(n16782), .B(n16739), .Y(n16781) );
  NAND2X1 U15296 ( .A(n42201), .B(n42970), .Y(n16782) );
  NAND2X1 U15300 ( .A(n73465), .B(n16769), .Y(n16780) );
  NAND2X1 U15305 ( .A(n16789), .B(n16790), .Y(n16740) );
  NAND2X1 U15306 ( .A(n16791), .B(n16775), .Y(n16790) );
  OR2X1 U15307 ( .A(n16792), .B(n16793), .Y(n16791) );
  NAND2X1 U15308 ( .A(n16793), .B(n16792), .Y(n16789) );
  NAND2X1 U15310 ( .A(n16796), .B(n16797), .Y(n16795) );
  NAND2X1 U15311 ( .A(n42989), .B(n16181), .Y(n16797) );
  NOR2X1 U15312 ( .A(n16798), .B(n16799), .Y(n16796) );
  NOR2X1 U15313 ( .A(n73460), .B(n42984), .Y(n16799) );
  NOR2X1 U15314 ( .A(n73462), .B(n42988), .Y(n16798) );
  NAND2X1 U15315 ( .A(n16800), .B(n16801), .Y(n16794) );
  NOR2X1 U15316 ( .A(n16802), .B(n16803), .Y(n16801) );
  NOR2X1 U15317 ( .A(n179), .B(n42945), .Y(n16803) );
  NOR2X1 U15318 ( .A(n340), .B(n42959), .Y(n16802) );
  NOR2X1 U15319 ( .A(n16804), .B(n16805), .Y(n16800) );
  NOR2X1 U15320 ( .A(n73474), .B(n15672), .Y(n16805) );
  NOR2X1 U15321 ( .A(n16506), .B(n15463), .Y(n16804) );
  NAND2X1 U15324 ( .A(n16810), .B(n16811), .Y(n16809) );
  NOR2X1 U15325 ( .A(n16812), .B(n16813), .Y(n16811) );
  NOR2X1 U15326 ( .A(n16101), .B(n40684), .Y(n16813) );
  AND2X1 U15327 ( .A(n16814), .B(n16815), .Y(n16101) );
  NOR2X1 U15328 ( .A(n42326), .B(n42321), .Y(n16814) );
  NOR2X1 U15330 ( .A(n16312), .B(n42944), .Y(n16812) );
  AND2X1 U15331 ( .A(n15464), .B(n16817), .Y(n16312) );
  NOR2X1 U15332 ( .A(n16818), .B(n16819), .Y(n16810) );
  NOR2X1 U15333 ( .A(n16098), .B(n42946), .Y(n16819) );
  NOR2X1 U15334 ( .A(n15462), .B(n42959), .Y(n16818) );
  NAND2X1 U15335 ( .A(n16820), .B(n16821), .Y(n16808) );
  NOR2X1 U15336 ( .A(n51), .B(n16822), .Y(n16821) );
  NOR2X1 U15337 ( .A(n16823), .B(n16775), .Y(n16822) );
  NOR2X1 U15338 ( .A(n16824), .B(n16825), .Y(n16823) );
  AND2X1 U15339 ( .A(n16792), .B(n16826), .Y(n16825) );
  NOR2X1 U15340 ( .A(n42299), .B(n16792), .Y(n16824) );
  NOR2X1 U15341 ( .A(n16828), .B(n16829), .Y(n16820) );
  NOR2X1 U15344 ( .A(n73468), .B(n16830), .Y(n16828) );
  NOR2X1 U15345 ( .A(n42972), .B(n16831), .Y(n16830) );
  NAND2X1 U15346 ( .A(n16832), .B(n16833), .Y(n16831) );
  NAND2X1 U15347 ( .A(n16834), .B(n16792), .Y(n16833) );
  NAND2X1 U15348 ( .A(n42299), .B(n42969), .Y(n16834) );
  NAND2X1 U15352 ( .A(n73467), .B(n16826), .Y(n16832) );
  NAND2X1 U15357 ( .A(n16841), .B(n16842), .Y(n16793) );
  NAND2X1 U15358 ( .A(n16843), .B(n15805), .Y(n16842) );
  OR2X1 U15359 ( .A(n16844), .B(n16845), .Y(n16843) );
  NAND2X1 U15360 ( .A(n16845), .B(n16844), .Y(n16841) );
  NAND2X1 U15362 ( .A(n16848), .B(n16849), .Y(n16847) );
  NAND2X1 U15363 ( .A(n42989), .B(n16563), .Y(n16849) );
  NOR2X1 U15364 ( .A(n16850), .B(n16851), .Y(n16848) );
  NOR2X1 U15365 ( .A(n226), .B(n43008), .Y(n16851) );
  NOR2X1 U15366 ( .A(n15492), .B(n43009), .Y(n16850) );
  NAND2X1 U15367 ( .A(n16852), .B(n16853), .Y(n16846) );
  NOR2X1 U15368 ( .A(n16854), .B(n16855), .Y(n16853) );
  NOR2X1 U15369 ( .A(n73464), .B(n42987), .Y(n16855) );
  NOR2X1 U15370 ( .A(n73476), .B(n15672), .Y(n16854) );
  NOR2X1 U15371 ( .A(n16856), .B(n16857), .Y(n16852) );
  NOR2X1 U15372 ( .A(n73462), .B(n42985), .Y(n16857) );
  NOR2X1 U15373 ( .A(n15495), .B(n43007), .Y(n16856) );
  NAND2X1 U15376 ( .A(n16862), .B(n16863), .Y(n16861) );
  NAND2X1 U15377 ( .A(n37341), .B(n16864), .Y(n16863) );
  NOR2X1 U15378 ( .A(n16865), .B(n16866), .Y(n16862) );
  NOR2X1 U15379 ( .A(n16867), .B(n15498), .Y(n16866) );
  NOR2X1 U15380 ( .A(n378), .B(n42959), .Y(n16865) );
  NAND2X1 U15381 ( .A(n16868), .B(n16869), .Y(n16860) );
  NOR2X1 U15382 ( .A(n16870), .B(n16871), .Y(n16869) );
  NOR2X1 U15383 ( .A(n73470), .B(n16872), .Y(n16871) );
  NOR2X1 U15384 ( .A(n361), .B(n16873), .Y(n16872) );
  NAND2X1 U15385 ( .A(n16874), .B(n16875), .Y(n16873) );
  NAND2X1 U15386 ( .A(n16876), .B(n16844), .Y(n16875) );
  NAND2X1 U15387 ( .A(n42202), .B(n42968), .Y(n16876) );
  NAND2X1 U15388 ( .A(n73469), .B(n16878), .Y(n16874) );
  NOR2X1 U15389 ( .A(n16879), .B(n15805), .Y(n16870) );
  NOR2X1 U15390 ( .A(n16880), .B(n16881), .Y(n16879) );
  AND2X1 U15391 ( .A(n16844), .B(n16878), .Y(n16881) );
  NOR2X1 U15396 ( .A(n42202), .B(n16844), .Y(n16880) );
  NAND2X1 U15399 ( .A(n16888), .B(n16889), .Y(n16845) );
  NAND2X1 U15400 ( .A(n16890), .B(n15846), .Y(n16889) );
  OR2X1 U15401 ( .A(n16891), .B(n16892), .Y(n16890) );
  NAND2X1 U15402 ( .A(n16892), .B(n16891), .Y(n16888) );
  NOR2X1 U15404 ( .A(n16893), .B(n16894), .Y(n16868) );
  NOR2X1 U15405 ( .A(n16166), .B(n40678), .Y(n16894) );
  NOR2X1 U15406 ( .A(n54), .B(n73396), .Y(n16166) );
  NOR2X1 U15407 ( .A(n300), .B(n15463), .Y(n16893) );
  NAND2X1 U15408 ( .A(n16895), .B(n16896), .Y(n16165) );
  NOR2X1 U15409 ( .A(n16897), .B(n16898), .Y(n16896) );
  NOR2X1 U15412 ( .A(n42448), .B(n16899), .Y(n16895) );
  NAND2X1 U15416 ( .A(n16902), .B(n16903), .Y(n16901) );
  NOR2X1 U15417 ( .A(n16904), .B(n16905), .Y(n16902) );
  NOR2X1 U15418 ( .A(n73476), .B(n40669), .Y(n16905) );
  NOR2X1 U15419 ( .A(n73474), .B(n42943), .Y(n16904) );
  NAND2X1 U15420 ( .A(n16906), .B(n16907), .Y(n16900) );
  NOR2X1 U15421 ( .A(n16908), .B(n16909), .Y(n16907) );
  NOR2X1 U15422 ( .A(n15828), .B(n15453), .Y(n16909) );
  NOR2X1 U15423 ( .A(n227), .B(n15505), .Y(n16908) );
  NOR2X1 U15424 ( .A(n16911), .B(n16912), .Y(n16906) );
  NOR2X1 U15425 ( .A(n73472), .B(n40674), .Y(n16912) );
  NOR2X1 U15426 ( .A(n15556), .B(n43007), .Y(n16911) );
  NAND2X1 U15429 ( .A(n16917), .B(n16918), .Y(n16916) );
  NAND2X1 U15430 ( .A(n42958), .B(n16182), .Y(n16918) );
  NOR2X1 U15431 ( .A(n16919), .B(n16920), .Y(n16917) );
  NOR2X1 U15432 ( .A(n309), .B(n40684), .Y(n16920) );
  NAND2X1 U15433 ( .A(n16921), .B(n16922), .Y(n16234) );
  NOR2X1 U15435 ( .A(n16923), .B(n42322), .Y(n16921) );
  NOR2X1 U15438 ( .A(n180), .B(n42946), .Y(n16919) );
  NAND2X1 U15439 ( .A(n16924), .B(n16925), .Y(n16233) );
  NOR2X1 U15440 ( .A(n16926), .B(n16927), .Y(n16925) );
  NOR2X1 U15443 ( .A(n42449), .B(n42457), .Y(n16924) );
  NAND2X1 U15445 ( .A(n16929), .B(n16930), .Y(n16915) );
  NAND2X1 U15446 ( .A(n16931), .B(n15846), .Y(n16930) );
  NAND2X1 U15447 ( .A(n16932), .B(n15416), .Y(n16931) );
  NOR2X1 U15448 ( .A(n16933), .B(n16934), .Y(n16932) );
  NOR2X1 U15449 ( .A(n42203), .B(n16891), .Y(n16934) );
  NOR2X1 U15450 ( .A(n73471), .B(n16936), .Y(n16933) );
  NOR2X1 U15451 ( .A(n980), .B(n16937), .Y(n16936) );
  NOR2X1 U15452 ( .A(n16938), .B(n16939), .Y(n16929) );
  NOR2X1 U15453 ( .A(n16940), .B(n15846), .Y(n16939) );
  NOR2X1 U15454 ( .A(n16941), .B(n16942), .Y(n16940) );
  NOR2X1 U15455 ( .A(n73471), .B(n42203), .Y(n16942) );
  AND2X1 U15460 ( .A(n16937), .B(n73471), .Y(n16941) );
  NAND2X1 U15463 ( .A(n16949), .B(n16950), .Y(n16892) );
  NAND2X1 U15464 ( .A(n16951), .B(n15977), .Y(n16950) );
  OR2X1 U15465 ( .A(n16952), .B(n16953), .Y(n16951) );
  NAND2X1 U15466 ( .A(n16953), .B(n16952), .Y(n16949) );
  NOR2X1 U15468 ( .A(n15410), .B(n15595), .Y(n16938) );
  NAND2X1 U15469 ( .A(n73433), .B(n16954), .Y(n15595) );
  NAND2X1 U15471 ( .A(n16903), .B(n16957), .Y(n16956) );
  NAND2X1 U15472 ( .A(n37341), .B(n16958), .Y(n16957) );
  NAND2X1 U15473 ( .A(n16959), .B(n16960), .Y(n16955) );
  NAND2X1 U15474 ( .A(n73570), .B(n16961), .Y(n16960) );
  NOR2X1 U15475 ( .A(n16962), .B(n16963), .Y(n16959) );
  NOR2X1 U15476 ( .A(n15610), .B(n42945), .Y(n16963) );
  NOR2X1 U15477 ( .A(n15607), .B(n43006), .Y(n16962) );
  NAND2X1 U15480 ( .A(n16968), .B(n16969), .Y(n16967) );
  NAND2X1 U15481 ( .A(n73512), .B(n15404), .Y(n16969) );
  NAND2X1 U15482 ( .A(n16970), .B(n16971), .Y(n15404) );
  NOR2X1 U15483 ( .A(n16972), .B(n16973), .Y(n16971) );
  NOR2X1 U15486 ( .A(n16974), .B(n16975), .Y(n16970) );
  NOR2X1 U15489 ( .A(n16976), .B(n16977), .Y(n16968) );
  NOR2X1 U15490 ( .A(n55), .B(n40678), .Y(n16977) );
  NAND2X1 U15491 ( .A(n16978), .B(n16979), .Y(n16299) );
  NOR2X1 U15492 ( .A(n16980), .B(n16981), .Y(n16979) );
  NOR2X1 U15495 ( .A(n16982), .B(n16983), .Y(n16978) );
  NOR2X1 U15498 ( .A(n15407), .B(n43009), .Y(n16976) );
  AND2X1 U15499 ( .A(n16984), .B(n16985), .Y(n15407) );
  NOR2X1 U15500 ( .A(n16986), .B(n16987), .Y(n16985) );
  NOR2X1 U15503 ( .A(n42452), .B(n37556), .Y(n16984) );
  NAND2X1 U15506 ( .A(n16988), .B(n16989), .Y(n16966) );
  OR2X1 U15507 ( .A(n43007), .B(n257), .Y(n16989) );
  NAND2X1 U15508 ( .A(n16990), .B(n16991), .Y(n16640) );
  NOR2X1 U15509 ( .A(n16992), .B(n16993), .Y(n16991) );
  NOR2X1 U15512 ( .A(n16994), .B(n16995), .Y(n16990) );
  NOR2X1 U15515 ( .A(n16996), .B(n16997), .Y(n16988) );
  NOR2X1 U15516 ( .A(n73474), .B(n16998), .Y(n16997) );
  NOR2X1 U15517 ( .A(n42971), .B(n16999), .Y(n16998) );
  NAND2X1 U15518 ( .A(n17000), .B(n17001), .Y(n16999) );
  NAND2X1 U15519 ( .A(n17002), .B(n16952), .Y(n17001) );
  NAND2X1 U15520 ( .A(n42204), .B(n42968), .Y(n17002) );
  NAND2X1 U15521 ( .A(n73473), .B(n17004), .Y(n17000) );
  NOR2X1 U15522 ( .A(n17005), .B(n15977), .Y(n16996) );
  NOR2X1 U15523 ( .A(n17006), .B(n17007), .Y(n17005) );
  AND2X1 U15524 ( .A(n16952), .B(n17004), .Y(n17007) );
  NOR2X1 U15529 ( .A(n42204), .B(n16952), .Y(n17006) );
  NAND2X1 U15532 ( .A(n17014), .B(n17015), .Y(n16953) );
  NAND2X1 U15533 ( .A(n17016), .B(n16042), .Y(n17015) );
  OR2X1 U15534 ( .A(n17017), .B(n17018), .Y(n17016) );
  NAND2X1 U15535 ( .A(n17018), .B(n17017), .Y(n17014) );
  NAND2X1 U15538 ( .A(n17021), .B(n16903), .Y(n17020) );
  NOR2X1 U15539 ( .A(n17022), .B(n17023), .Y(n17021) );
  NOR2X1 U15540 ( .A(n16632), .B(n15498), .Y(n17023) );
  AND2X1 U15541 ( .A(n17024), .B(n17025), .Y(n16632) );
  NOR2X1 U15543 ( .A(n42311), .B(n42319), .Y(n17024) );
  NOR2X1 U15546 ( .A(n16506), .B(n15465), .Y(n17022) );
  AND2X1 U15547 ( .A(n17027), .B(n17028), .Y(n16506) );
  NOR2X1 U15549 ( .A(n17029), .B(n42456), .Y(n17027) );
  NAND2X1 U15552 ( .A(n17030), .B(n17031), .Y(n17019) );
  NAND2X1 U15553 ( .A(n73511), .B(n16298), .Y(n17031) );
  NAND2X1 U15554 ( .A(n17032), .B(n17033), .Y(n16298) );
  NOR2X1 U15555 ( .A(n17034), .B(n17035), .Y(n17033) );
  NOR2X1 U15558 ( .A(n17036), .B(n17037), .Y(n17032) );
  NOR2X1 U15561 ( .A(n17038), .B(n17039), .Y(n17030) );
  NOR2X1 U15562 ( .A(n15450), .B(n43008), .Y(n17039) );
  AND2X1 U15563 ( .A(n17040), .B(n17041), .Y(n15450) );
  NOR2X1 U15564 ( .A(n17042), .B(n42317), .Y(n17041) );
  NOR2X1 U15567 ( .A(n17043), .B(n17044), .Y(n17040) );
  NOR2X1 U15570 ( .A(n42454), .B(n42959), .Y(n17038) );
  NOR2X1 U15580 ( .A(n17054), .B(n17055), .Y(n17052) );
  NOR2X1 U15581 ( .A(n73494), .B(n15672), .Y(n17055) );
  NOR2X1 U15583 ( .A(n16098), .B(n15465), .Y(n17054) );
  AND2X1 U15584 ( .A(n17056), .B(n17057), .Y(n16098) );
  NOR2X1 U15586 ( .A(n17058), .B(n42459), .Y(n17056) );
  NAND2X1 U15588 ( .A(n17060), .B(n17061), .Y(n17050) );
  NOR2X1 U15589 ( .A(n17062), .B(n17063), .Y(n17061) );
  NOR2X1 U15590 ( .A(n73476), .B(n17064), .Y(n17063) );
  NOR2X1 U15591 ( .A(n42972), .B(n17065), .Y(n17064) );
  NAND2X1 U15592 ( .A(n17066), .B(n17067), .Y(n17065) );
  NAND2X1 U15593 ( .A(n17068), .B(n17017), .Y(n17067) );
  NAND2X1 U15594 ( .A(n42300), .B(n42968), .Y(n17068) );
  NAND2X1 U15595 ( .A(n73475), .B(n17070), .Y(n17066) );
  NOR2X1 U15596 ( .A(n17071), .B(n16042), .Y(n17062) );
  NOR2X1 U15597 ( .A(n17072), .B(n17073), .Y(n17071) );
  AND2X1 U15598 ( .A(n17017), .B(n17070), .Y(n17073) );
  NOR2X1 U15603 ( .A(n42300), .B(n17017), .Y(n17072) );
  NAND2X1 U15606 ( .A(n17080), .B(n17081), .Y(n17018) );
  NAND2X1 U15607 ( .A(n17082), .B(n15728), .Y(n17081) );
  OR2X1 U15608 ( .A(n318), .B(n17083), .Y(n17082) );
  NAND2X1 U15609 ( .A(n17083), .B(n318), .Y(n17080) );
  NOR2X1 U15611 ( .A(n17084), .B(n17085), .Y(n17060) );
  NOR2X1 U15612 ( .A(n15462), .B(n42944), .Y(n17085) );
  AND2X1 U15613 ( .A(n17086), .B(n17087), .Y(n15462) );
  NOR2X1 U15614 ( .A(n17088), .B(n17089), .Y(n17087) );
  NOR2X1 U15617 ( .A(n17090), .B(n17091), .Y(n17086) );
  NOR2X1 U15620 ( .A(n15464), .B(n15463), .Y(n17084) );
  AND2X1 U15621 ( .A(n17092), .B(n17093), .Y(n15464) );
  NOR2X1 U15623 ( .A(n42450), .B(n17095), .Y(n17092) );
  NAND2X1 U15626 ( .A(n17099), .B(n16903), .Y(n17097) );
  NOR2X1 U15627 ( .A(n17101), .B(n17103), .Y(n17099) );
  NOR2X1 U15628 ( .A(n15495), .B(n15491), .Y(n17103) );
  NOR2X1 U15629 ( .A(n215), .B(n15505), .Y(n17101) );
  NAND2X1 U15630 ( .A(n17104), .B(n17105), .Y(n17096) );
  NAND2X1 U15631 ( .A(n37341), .B(n17106), .Y(n17105) );
  NOR2X1 U15632 ( .A(n17107), .B(n17108), .Y(n17104) );
  NOR2X1 U15633 ( .A(n17109), .B(n15498), .Y(n17108) );
  NOR2X1 U15634 ( .A(n15492), .B(n43006), .Y(n17107) );
  NAND2X1 U15637 ( .A(n17114), .B(n17115), .Y(n17113) );
  NAND2X1 U15638 ( .A(n37341), .B(n16910), .Y(n17115) );
  NAND2X1 U15639 ( .A(n17116), .B(n17117), .Y(n16910) );
  NOR2X1 U15640 ( .A(n17118), .B(n42314), .Y(n17117) );
  NOR2X1 U15643 ( .A(n17119), .B(n17120), .Y(n17116) );
  NOR2X1 U15646 ( .A(n17121), .B(n17122), .Y(n17114) );
  NOR2X1 U15647 ( .A(n256), .B(n43006), .Y(n17122) );
  NAND2X1 U15648 ( .A(n17123), .B(n17124), .Y(n16864) );
  NOR2X1 U15649 ( .A(n17125), .B(n17126), .Y(n17124) );
  NOR2X1 U15652 ( .A(n17127), .B(n17128), .Y(n17123) );
  NOR2X1 U15655 ( .A(n15726), .B(n15498), .Y(n17121) );
  AND2X1 U15656 ( .A(n17129), .B(n17130), .Y(n15726) );
  NOR2X1 U15658 ( .A(n17131), .B(n42324), .Y(n17129) );
  NAND2X1 U15661 ( .A(n17132), .B(n17133), .Y(n17112) );
  NOR2X1 U15662 ( .A(n17134), .B(n17135), .Y(n17133) );
  NOR2X1 U15663 ( .A(n73478), .B(n17136), .Y(n17135) );
  NOR2X1 U15664 ( .A(n361), .B(n17137), .Y(n17136) );
  NAND2X1 U15665 ( .A(n17138), .B(n17139), .Y(n17137) );
  NAND2X1 U15666 ( .A(n17140), .B(n318), .Y(n17139) );
  NAND2X1 U15667 ( .A(n42301), .B(n42968), .Y(n17140) );
  NAND2X1 U15668 ( .A(n73477), .B(n17143), .Y(n17138) );
  NOR2X1 U15669 ( .A(n17144), .B(n15728), .Y(n17134) );
  NOR2X1 U15670 ( .A(n17145), .B(n17146), .Y(n17144) );
  AND2X1 U15671 ( .A(n318), .B(n17143), .Y(n17146) );
  NOR2X1 U15676 ( .A(n42301), .B(n318), .Y(n17145) );
  NAND2X1 U15679 ( .A(n17153), .B(n17154), .Y(n17083) );
  NAND2X1 U15680 ( .A(n17155), .B(n15845), .Y(n17154) );
  OR2X1 U15681 ( .A(n330), .B(n17156), .Y(n17155) );
  NAND2X1 U15682 ( .A(n17156), .B(n330), .Y(n17153) );
  NOR2X1 U15684 ( .A(n17157), .B(n17158), .Y(n17132) );
  NOR2X1 U15685 ( .A(n15514), .B(n43008), .Y(n17158) );
  AND2X1 U15686 ( .A(n16867), .B(n17159), .Y(n15514) );
  AND2X1 U15688 ( .A(n17160), .B(n16668), .Y(n16867) );
  NOR2X1 U15693 ( .A(n15496), .B(n15530), .Y(n17157) );
  NAND2X1 U15696 ( .A(n17166), .B(n16903), .Y(n17165) );
  AND2X1 U15697 ( .A(n17167), .B(n15735), .Y(n16903) );
  NAND2X1 U15698 ( .A(n51), .B(n15734), .Y(n17167) );
  NOR2X1 U15699 ( .A(n17168), .B(n17169), .Y(n17166) );
  NOR2X1 U15700 ( .A(n73494), .B(n40669), .Y(n17169) );
  NOR2X1 U15701 ( .A(n73482), .B(n362), .Y(n17168) );
  NAND2X1 U15702 ( .A(n17170), .B(n17171), .Y(n17164) );
  NOR2X1 U15703 ( .A(n17172), .B(n17173), .Y(n17171) );
  NOR2X1 U15704 ( .A(n15828), .B(n42946), .Y(n17173) );
  AND2X1 U15705 ( .A(n17174), .B(n17175), .Y(n15828) );
  NOR2X1 U15706 ( .A(n17176), .B(n17177), .Y(n17175) );
  NOR2X1 U15709 ( .A(n17178), .B(n17179), .Y(n17174) );
  NOR2X1 U15712 ( .A(n378), .B(n42945), .Y(n17172) );
  NAND2X1 U15713 ( .A(n17180), .B(n17181), .Y(n16113) );
  NOR2X1 U15714 ( .A(n17182), .B(n17183), .Y(n17181) );
  NOR2X1 U15720 ( .A(n17186), .B(n17187), .Y(n17170) );
  NOR2X1 U15721 ( .A(n73480), .B(n40674), .Y(n17187) );
  NOR2X1 U15722 ( .A(n15556), .B(n40678), .Y(n17186) );
  AND2X1 U15723 ( .A(n17188), .B(n17189), .Y(n15556) );
  NOR2X1 U15724 ( .A(n17190), .B(n17191), .Y(n17189) );
  NOR2X1 U15727 ( .A(n17192), .B(n17193), .Y(n17188) );
  NAND2X1 U15732 ( .A(n17198), .B(n17199), .Y(n17197) );
  NOR2X1 U15733 ( .A(n17200), .B(n17201), .Y(n17199) );
  NOR2X1 U15734 ( .A(n73482), .B(n40674), .Y(n17201) );
  NOR2X1 U15736 ( .A(n42303), .B(n17203), .Y(n17200) );
  NOR2X1 U15737 ( .A(n17204), .B(n17205), .Y(n17198) );
  NOR2X1 U15738 ( .A(n73484), .B(n40669), .Y(n17205) );
  NOR2X1 U15740 ( .A(n73494), .B(n42943), .Y(n17204) );
  NAND2X1 U15742 ( .A(n17206), .B(n17207), .Y(n17196) );
  NOR2X1 U15743 ( .A(n17316), .B(n17317), .Y(n17207) );
  NAND2X1 U15744 ( .A(n17318), .B(n15735), .Y(n17317) );
  NAND2X1 U15745 ( .A(n51), .B(n15742), .Y(n15735) );
  NAND2X1 U15746 ( .A(n17319), .B(n73572), .Y(n17318) );
  NOR2X1 U15747 ( .A(n73433), .B(n48), .Y(n17319) );
  NAND2X1 U15748 ( .A(n17320), .B(n17321), .Y(n16954) );
  NAND2X1 U15749 ( .A(n51), .B(n16593), .Y(n17321) );
  NAND2X1 U15750 ( .A(n54), .B(n15682), .Y(n16351) );
  NOR2X1 U15752 ( .A(n73513), .B(n73438), .Y(n17322) );
  NOR2X1 U15753 ( .A(n17324), .B(n17325), .Y(n17320) );
  NOR2X1 U15754 ( .A(n73489), .B(n16723), .Y(n17325) );
  AND2X1 U15755 ( .A(n17326), .B(n17327), .Y(n16723) );
  NOR2X1 U15758 ( .A(n17328), .B(n15682), .Y(n17324) );
  NOR2X1 U15764 ( .A(n17332), .B(n15845), .Y(n17316) );
  NOR2X1 U15765 ( .A(n17333), .B(n17334), .Y(n17332) );
  NOR2X1 U15766 ( .A(n73479), .B(n42303), .Y(n17334) );
  AND2X1 U15771 ( .A(n17340), .B(n73479), .Y(n17333) );
  NOR2X1 U15772 ( .A(n17341), .B(n17342), .Y(n17206) );
  NOR2X1 U15773 ( .A(n73472), .B(n15649), .Y(n17342) );
  NOR2X1 U15774 ( .A(n73480), .B(n17343), .Y(n17341) );
  NOR2X1 U15775 ( .A(n17344), .B(n42971), .Y(n17343) );
  NOR2X1 U15776 ( .A(n73479), .B(n17345), .Y(n17344) );
  NOR2X1 U15777 ( .A(n980), .B(n17340), .Y(n17345) );
  NAND2X1 U15780 ( .A(n17348), .B(n17349), .Y(n17156) );
  NAND2X1 U15781 ( .A(n17350), .B(n15414), .Y(n17349) );
  OR2X1 U15782 ( .A(n15433), .B(n15420), .Y(n17350) );
  NAND2X1 U15783 ( .A(n15433), .B(n15420), .Y(n17348) );
  NAND2X1 U15784 ( .A(n17351), .B(n17352), .Y(n15433) );
  NAND2X1 U15785 ( .A(n17353), .B(n15447), .Y(n17352) );
  OR2X1 U15786 ( .A(n17354), .B(n15481), .Y(n17353) );
  NAND2X1 U15787 ( .A(n15481), .B(n17354), .Y(n17351) );
  NAND2X1 U15788 ( .A(n17355), .B(n17356), .Y(n15481) );
  NAND2X1 U15789 ( .A(n17357), .B(n15441), .Y(n17356) );
  OR2X1 U15790 ( .A(n15524), .B(n15539), .Y(n17357) );
  NAND2X1 U15791 ( .A(n15539), .B(n15524), .Y(n17355) );
  NAND2X1 U15792 ( .A(n17358), .B(n17359), .Y(n15539) );
  NAND2X1 U15793 ( .A(n17360), .B(n15443), .Y(n17359) );
  OR2X1 U15794 ( .A(n17361), .B(n15580), .Y(n17360) );
  NAND2X1 U15795 ( .A(n15580), .B(n17361), .Y(n17358) );
  NAND2X1 U15796 ( .A(n17362), .B(n17363), .Y(n15580) );
  NAND2X1 U15797 ( .A(n17364), .B(n17094), .Y(n17363) );
  OR2X1 U15798 ( .A(n15633), .B(n15641), .Y(n17364) );
  NAND2X1 U15799 ( .A(n15641), .B(n15633), .Y(n17362) );
  NAND2X1 U15800 ( .A(n17365), .B(n17366), .Y(n15641) );
  NAND2X1 U15801 ( .A(n17367), .B(n15682), .Y(n17366) );
  OR2X1 U15802 ( .A(n15679), .B(n15695), .Y(n17367) );
  NAND2X1 U15803 ( .A(n15695), .B(n15679), .Y(n17365) );
  NAND2X1 U15804 ( .A(n17368), .B(n17369), .Y(n15695) );
  NAND2X1 U15805 ( .A(n17370), .B(n15742), .Y(n17369) );
  OR2X1 U15806 ( .A(n15739), .B(n15756), .Y(n17370) );
  NAND2X1 U15807 ( .A(n15756), .B(n15739), .Y(n17368) );
  NAND2X1 U15808 ( .A(n17371), .B(n17372), .Y(n15756) );
  NAND2X1 U15809 ( .A(n17373), .B(n15734), .Y(n17372) );
  OR2X1 U15810 ( .A(n15919), .B(n15932), .Y(n17373) );
  NAND2X1 U15811 ( .A(n15932), .B(n15919), .Y(n17371) );
  NAND2X1 U15813 ( .A(n17376), .B(n16593), .Y(n17375) );
  NAND2X1 U15818 ( .A(n17380), .B(n17381), .Y(n17379) );
  NOR2X1 U15819 ( .A(n17382), .B(n17383), .Y(n17381) );
  NOR2X1 U15820 ( .A(n73476), .B(n42988), .Y(n17383) );
  NOR2X1 U15821 ( .A(n255), .B(n43006), .Y(n17382) );
  NAND2X1 U15822 ( .A(n17384), .B(n17385), .Y(n16958) );
  NOR2X1 U15823 ( .A(n17386), .B(n17387), .Y(n17385) );
  NOR2X1 U15826 ( .A(n37552), .B(n17388), .Y(n17384) );
  NOR2X1 U15829 ( .A(n17389), .B(n17390), .Y(n17380) );
  NOR2X1 U15830 ( .A(n73478), .B(n360), .Y(n17390) );
  NOR2X1 U15831 ( .A(n73474), .B(n358), .Y(n17389) );
  NAND2X1 U15832 ( .A(n17391), .B(n17392), .Y(n17378) );
  NOR2X1 U15833 ( .A(n17393), .B(n17394), .Y(n17392) );
  NOR2X1 U15834 ( .A(n15610), .B(n42946), .Y(n17394) );
  AND2X1 U15836 ( .A(n17395), .B(n17396), .Y(n15610) );
  NOR2X1 U15837 ( .A(n17397), .B(n17398), .Y(n17396) );
  NOR2X1 U15840 ( .A(n17399), .B(n42458), .Y(n17395) );
  NOR2X1 U15843 ( .A(n15607), .B(n40678), .Y(n17393) );
  AND2X1 U15844 ( .A(n17400), .B(n17401), .Y(n15607) );
  NOR2X1 U15845 ( .A(n17402), .B(n17403), .Y(n17401) );
  NOR2X1 U15848 ( .A(n17404), .B(n17405), .Y(n17400) );
  NOR2X1 U15851 ( .A(n17406), .B(n17407), .Y(n17391) );
  NOR2X1 U15852 ( .A(n73397), .B(n42944), .Y(n17407) );
  NOR2X1 U15860 ( .A(n216), .B(n43009), .Y(n17406) );
  NAND2X1 U15861 ( .A(n17413), .B(n17414), .Y(n16961) );
  NOR2X1 U15862 ( .A(n42313), .B(n17415), .Y(n17414) );
  NOR2X1 U15865 ( .A(n17416), .B(n17417), .Y(n17413) );
  NOR2X1 U15872 ( .A(n15687), .B(n43009), .Y(n17425) );
  AND2X1 U15874 ( .A(n15497), .B(n16817), .Y(n15687) );
  AND2X1 U15876 ( .A(n17426), .B(n17427), .Y(n15497) );
  NOR2X1 U15878 ( .A(n42449), .B(n42459), .Y(n17426) );
  OR2X1 U15895 ( .A(n17446), .B(n73438), .Y(n17444) );
  NAND2X1 U15897 ( .A(n17447), .B(n17448), .Y(n17446) );
  NAND2X1 U15898 ( .A(n73439), .B(n17449), .Y(n17448) );
  NAND2X1 U15899 ( .A(n73440), .B(n17450), .Y(n17449) );
  OR2X1 U15900 ( .A(n17450), .B(n73440), .Y(n17447) );
  NAND2X1 U15901 ( .A(n17451), .B(n17452), .Y(n17450) );
  NAND2X1 U15902 ( .A(n17453), .B(n17454), .Y(n17452) );
  NAND2X1 U15903 ( .A(n73442), .B(n15875), .Y(n17454) );
  NOR2X1 U15904 ( .A(n17455), .B(n17456), .Y(n17453) );
  AND2X1 U15905 ( .A(n16004), .B(n17457), .Y(n17456) );
  NOR2X1 U15906 ( .A(n17458), .B(n16003), .Y(n17455) );
  NOR2X1 U15907 ( .A(n16004), .B(n17457), .Y(n17458) );
  NAND2X1 U15908 ( .A(n17459), .B(n17460), .Y(n17457) );
  NAND2X1 U15909 ( .A(n73446), .B(n17461), .Y(n17460) );
  OR2X1 U15910 ( .A(n17462), .B(n16078), .Y(n17461) );
  NAND2X1 U15911 ( .A(n17462), .B(n16078), .Y(n17459) );
  NAND2X1 U15912 ( .A(n17463), .B(n17464), .Y(n17462) );
  NAND2X1 U15913 ( .A(n73448), .B(n17465), .Y(n17464) );
  NAND2X1 U15914 ( .A(n73447), .B(n17466), .Y(n17465) );
  OR2X1 U15915 ( .A(n17466), .B(n73447), .Y(n17463) );
  NAND2X1 U15916 ( .A(n17467), .B(n17468), .Y(n17466) );
  NAND2X1 U15917 ( .A(n17469), .B(n17470), .Y(n17468) );
  NAND2X1 U15918 ( .A(n73450), .B(n16214), .Y(n17470) );
  NOR2X1 U15919 ( .A(n17471), .B(n17472), .Y(n17469) );
  AND2X1 U15920 ( .A(n16278), .B(n17473), .Y(n17472) );
  NOR2X1 U15921 ( .A(n17474), .B(n16047), .Y(n17471) );
  NOR2X1 U15922 ( .A(n16278), .B(n17473), .Y(n17474) );
  NAND2X1 U15923 ( .A(n17475), .B(n17476), .Y(n17473) );
  NAND2X1 U15924 ( .A(n73454), .B(n17477), .Y(n17476) );
  OR2X1 U15925 ( .A(n17478), .B(n16338), .Y(n17477) );
  NAND2X1 U15926 ( .A(n17478), .B(n16338), .Y(n17475) );
  NAND2X1 U15927 ( .A(n17479), .B(n17480), .Y(n17478) );
  NAND2X1 U15928 ( .A(n73456), .B(n17481), .Y(n17480) );
  NAND2X1 U15929 ( .A(n73455), .B(n17482), .Y(n17481) );
  OR2X1 U15930 ( .A(n17482), .B(n73455), .Y(n17479) );
  NAND2X1 U15931 ( .A(n17483), .B(n17484), .Y(n17482) );
  NAND2X1 U15932 ( .A(n17485), .B(n17486), .Y(n17484) );
  NAND2X1 U15933 ( .A(n73458), .B(n16450), .Y(n17486) );
  NOR2X1 U15934 ( .A(n17487), .B(n17488), .Y(n17485) );
  AND2X1 U15935 ( .A(n16504), .B(n17489), .Y(n17488) );
  NOR2X1 U15936 ( .A(n17490), .B(n16048), .Y(n17487) );
  NOR2X1 U15937 ( .A(n16504), .B(n17489), .Y(n17490) );
  NAND2X1 U15938 ( .A(n17491), .B(n17492), .Y(n17489) );
  NAND2X1 U15939 ( .A(n73462), .B(n17493), .Y(n17492) );
  OR2X1 U15940 ( .A(n17494), .B(n16557), .Y(n17493) );
  NAND2X1 U15941 ( .A(n17494), .B(n16557), .Y(n17491) );
  NAND2X1 U15942 ( .A(n17495), .B(n17496), .Y(n17494) );
  NAND2X1 U15943 ( .A(n73464), .B(n17497), .Y(n17496) );
  NAND2X1 U15944 ( .A(n73463), .B(n17498), .Y(n17497) );
  OR2X1 U15945 ( .A(n17498), .B(n73463), .Y(n17495) );
  NAND2X1 U15946 ( .A(n17499), .B(n17500), .Y(n17498) );
  NAND2X1 U15947 ( .A(n17501), .B(n17502), .Y(n17500) );
  NAND2X1 U15948 ( .A(n73466), .B(n16739), .Y(n17502) );
  NOR2X1 U15949 ( .A(n17503), .B(n17504), .Y(n17501) );
  AND2X1 U15950 ( .A(n16792), .B(n17505), .Y(n17504) );
  NOR2X1 U15951 ( .A(n17506), .B(n16775), .Y(n17503) );
  NOR2X1 U15952 ( .A(n16792), .B(n17505), .Y(n17506) );
  NAND2X1 U15953 ( .A(n17507), .B(n17508), .Y(n17505) );
  NAND2X1 U15954 ( .A(n73470), .B(n17509), .Y(n17508) );
  OR2X1 U15955 ( .A(n17510), .B(n16844), .Y(n17509) );
  NAND2X1 U15956 ( .A(n17510), .B(n16844), .Y(n17507) );
  NAND2X1 U15957 ( .A(n17511), .B(n17512), .Y(n17510) );
  NAND2X1 U15958 ( .A(n73472), .B(n17513), .Y(n17512) );
  NAND2X1 U15959 ( .A(n73471), .B(n17514), .Y(n17513) );
  OR2X1 U15960 ( .A(n17514), .B(n73471), .Y(n17511) );
  NAND2X1 U15961 ( .A(n17515), .B(n17516), .Y(n17514) );
  NAND2X1 U15962 ( .A(n17517), .B(n17518), .Y(n17516) );
  NAND2X1 U15963 ( .A(n73474), .B(n16952), .Y(n17518) );
  NOR2X1 U15964 ( .A(n17519), .B(n17520), .Y(n17517) );
  NOR2X1 U15965 ( .A(n73475), .B(n17521), .Y(n17520) );
  NOR2X1 U15966 ( .A(n17522), .B(n16042), .Y(n17519) );
  AND2X1 U15967 ( .A(n17521), .B(n73475), .Y(n17522) );
  NAND2X1 U15968 ( .A(n17523), .B(n17524), .Y(n17521) );
  NAND2X1 U15969 ( .A(n17525), .B(n17526), .Y(n17524) );
  NAND2X1 U15970 ( .A(n73478), .B(n318), .Y(n17526) );
  NOR2X1 U15971 ( .A(n17527), .B(n17528), .Y(n17525) );
  NOR2X1 U15972 ( .A(n73479), .B(n15845), .Y(n17528) );
  NOR2X1 U15973 ( .A(n17529), .B(n17530), .Y(n17527) );
  NOR2X1 U15974 ( .A(n17531), .B(n17532), .Y(n17530) );
  NAND2X1 U15975 ( .A(n17533), .B(n17534), .Y(n17532) );
  NAND2X1 U15977 ( .A(n73480), .B(n15420), .Y(n17533) );
  NOR2X1 U15981 ( .A(n17539), .B(n17540), .Y(n17529) );
  NAND2X1 U15982 ( .A(n17541), .B(n17542), .Y(n17540) );
  NAND2X1 U15983 ( .A(n17543), .B(n17544), .Y(n17542) );
  NAND2X1 U15984 ( .A(n17545), .B(n17546), .Y(n17544) );
  NAND2X1 U15985 ( .A(n73484), .B(n15524), .Y(n17546) );
  NOR2X1 U15986 ( .A(n17547), .B(n17548), .Y(n17545) );
  NOR2X1 U15987 ( .A(n73485), .B(n15443), .Y(n17548) );
  NOR2X1 U15988 ( .A(n17549), .B(n17550), .Y(n17547) );
  NOR2X1 U15989 ( .A(n17551), .B(n17552), .Y(n17550) );
  NAND2X1 U15990 ( .A(n17553), .B(n17554), .Y(n17552) );
  NAND2X1 U15991 ( .A(n73488), .B(n15567), .Y(n17554) );
  NAND2X1 U15992 ( .A(n73486), .B(n15633), .Y(n17553) );
  NOR2X1 U15998 ( .A(n17560), .B(n17561), .Y(n17549) );
  NAND2X1 U15999 ( .A(n17562), .B(n17563), .Y(n17561) );
  NAND2X1 U16000 ( .A(n17564), .B(n15682), .Y(n17563) );
  NAND2X1 U16001 ( .A(n15679), .B(n17565), .Y(n17564) );
  OR2X1 U16002 ( .A(n17565), .B(n15679), .Y(n17562) );
  NAND2X1 U16003 ( .A(n17566), .B(n17567), .Y(n17565) );
  NAND2X1 U16004 ( .A(n17568), .B(n17569), .Y(n17567) );
  NAND2X1 U16005 ( .A(n73495), .B(n15742), .Y(n17569) );
  NOR2X1 U16006 ( .A(n17570), .B(n17571), .Y(n17568) );
  AND2X1 U16007 ( .A(n17572), .B(n73491), .Y(n17571) );
  NOR2X1 U16008 ( .A(n73433), .B(n17573), .Y(n17570) );
  NOR2X1 U16009 ( .A(n73491), .B(n17572), .Y(n17573) );
  NAND2X1 U16014 ( .A(n73525), .B(n15739), .Y(n17566) );
  NOR2X1 U16015 ( .A(n73487), .B(n17094), .Y(n17560) );
  NAND2X1 U16016 ( .A(n17577), .B(n17578), .Y(n17543) );
  NOR2X1 U16022 ( .A(n17584), .B(n17585), .Y(n17577) );
  NOR2X1 U16023 ( .A(n73483), .B(n15447), .Y(n17585) );
  AND2X1 U16024 ( .A(n15476), .B(n73484), .Y(n17584) );
  NOR2X1 U16025 ( .A(n73481), .B(n15414), .Y(n17539) );
  NAND2X1 U16026 ( .A(n73477), .B(n15728), .Y(n17523) );
  NAND2X1 U16027 ( .A(n73473), .B(n15977), .Y(n17515) );
  NAND2X1 U16028 ( .A(n73465), .B(n16563), .Y(n17499) );
  NAND2X1 U16029 ( .A(n73457), .B(n16449), .Y(n17483) );
  NAND2X1 U16030 ( .A(n73449), .B(n16213), .Y(n17467) );
  NAND2X1 U16031 ( .A(n73441), .B(n15874), .Y(n17451) );
  AND2X1 U16282 ( .A(n17768), .B(n17769), .Y(n15495) );
  NOR2X1 U16283 ( .A(n17770), .B(n17771), .Y(n17769) );
  NOR2X1 U16296 ( .A(n17781), .B(n17782), .Y(n17768) );
  NAND2X1 U16317 ( .A(n17796), .B(n16080), .Y(n15749) );
  NAND2X1 U16336 ( .A(n73573), .B(n73572), .Y(n15505) );
  NOR2X1 U16342 ( .A(n17810), .B(n17811), .Y(n17809) );
  NOR2X1 U16343 ( .A(n226), .B(n15496), .Y(n17811) );
  NAND2X1 U16344 ( .A(n73432), .B(n73572), .Y(n15496) );
  NAND2X1 U16346 ( .A(n17812), .B(n17813), .Y(n17106) );
  NOR2X1 U16347 ( .A(n17814), .B(n17815), .Y(n17813) );
  NOR2X1 U16360 ( .A(n17824), .B(n42312), .Y(n17812) );
  NOR2X1 U16373 ( .A(n215), .B(n40678), .Y(n17810) );
  NAND2X1 U16374 ( .A(n16342), .B(n73572), .Y(n15491) );
  NAND2X1 U16375 ( .A(n17833), .B(n17834), .Y(n15501) );
  NOR2X1 U16376 ( .A(n17835), .B(n17836), .Y(n17834) );
  NOR2X1 U16389 ( .A(n42320), .B(n17845), .Y(n17833) );
  NOR2X1 U16402 ( .A(n17854), .B(n17855), .Y(n17808) );
  NOR2X1 U16403 ( .A(n15492), .B(n15529), .Y(n17855) );
  NAND2X1 U16404 ( .A(n73524), .B(n16342), .Y(n15529) );
  NOR2X1 U16405 ( .A(n15734), .B(n73489), .Y(n16342) );
  AND2X1 U16406 ( .A(n17856), .B(n17857), .Y(n15492) );
  NOR2X1 U16407 ( .A(n17858), .B(n17859), .Y(n17857) );
  NOR2X1 U16420 ( .A(n17868), .B(n17869), .Y(n17856) );
  NOR2X1 U16433 ( .A(n73492), .B(n42991), .Y(n17854) );
  NOR2X1 U16440 ( .A(n73491), .B(n42987), .Y(n17883) );
  NOR2X1 U16454 ( .A(n17898), .B(n17899), .Y(n17896) );
  NOR2X1 U16456 ( .A(n17900), .B(n1009), .Y(n17898) );
  NOR2X1 U16466 ( .A(n17909), .B(n17910), .Y(n17880) );
  NOR2X1 U16467 ( .A(n73495), .B(n42984), .Y(n17910) );
  NAND2X1 U16469 ( .A(n73572), .B(n73571), .Y(n15498) );
  NAND2X1 U16470 ( .A(n73489), .B(n73433), .Y(n16635) );
  NAND2X1 U16471 ( .A(n73525), .B(n42455), .Y(n15410) );
  NOR2X1 U16475 ( .A(n15504), .B(n43006), .Y(n17909) );
  NAND2X1 U16476 ( .A(n73524), .B(n73573), .Y(n15408) );
  NAND2X1 U16477 ( .A(n73489), .B(n15734), .Y(n16631) );
  NAND2X1 U16504 ( .A(n42434), .B(n17938), .Y(n17937) );
  AND2X1 U16505 ( .A(n17109), .B(n16566), .Y(n15504) );
  AND2X1 U16513 ( .A(n17943), .B(n17944), .Y(n17109) );
  NOR2X1 U16521 ( .A(n17949), .B(n42321), .Y(n17943) );
  NOR2X1 U16604 ( .A(n44803), .B(n37638), .Y(n18000) );
  NOR2X1 U16608 ( .A(n44806), .B(n37609), .Y(n18003) );
  NOR2X1 U16611 ( .A(n44803), .B(n37637), .Y(n18009) );
  NOR2X1 U16615 ( .A(n44806), .B(n37608), .Y(n18011) );
  NOR2X1 U16618 ( .A(n44803), .B(n37636), .Y(n18016) );
  NOR2X1 U16622 ( .A(n44806), .B(n37607), .Y(n18018) );
  NOR2X1 U16625 ( .A(n44803), .B(n37635), .Y(n18023) );
  NOR2X1 U16629 ( .A(n44806), .B(n37606), .Y(n18025) );
  NOR2X1 U16632 ( .A(n44803), .B(n37634), .Y(n18030) );
  NOR2X1 U16636 ( .A(n44806), .B(n37605), .Y(n18032) );
  NOR2X1 U16639 ( .A(n44803), .B(n37662), .Y(n18037) );
  NOR2X1 U16643 ( .A(n44806), .B(n37633), .Y(n18039) );
  NOR2X1 U16646 ( .A(n44803), .B(n37661), .Y(n18044) );
  NOR2X1 U16650 ( .A(n44806), .B(n37632), .Y(n18046) );
  NOR2X1 U16653 ( .A(n44803), .B(n37660), .Y(n18051) );
  NOR2X1 U16657 ( .A(n44806), .B(n37631), .Y(n18053) );
  NOR2X1 U16660 ( .A(n44803), .B(n37659), .Y(n18058) );
  NOR2X1 U16664 ( .A(n44806), .B(n37630), .Y(n18060) );
  NOR2X1 U16667 ( .A(n44803), .B(n37658), .Y(n18065) );
  NOR2X1 U16671 ( .A(n44806), .B(n37629), .Y(n18067) );
  NOR2X1 U16674 ( .A(n44803), .B(n37604), .Y(n18072) );
  NOR2X1 U16678 ( .A(n44806), .B(n37601), .Y(n18074) );
  NOR2X1 U16681 ( .A(n44803), .B(n37603), .Y(n18079) );
  NOR2X1 U16685 ( .A(n44806), .B(n37600), .Y(n18081) );
  NOR2X1 U16688 ( .A(n44797), .B(n37657), .Y(n18086) );
  NOR2X1 U16692 ( .A(n44800), .B(n37628), .Y(n18089) );
  NOR2X1 U16695 ( .A(n44797), .B(n37656), .Y(n18095) );
  NOR2X1 U16699 ( .A(n44800), .B(n37627), .Y(n18097) );
  NOR2X1 U16702 ( .A(n44797), .B(n37655), .Y(n18102) );
  NOR2X1 U16706 ( .A(n44800), .B(n37626), .Y(n18104) );
  NOR2X1 U16709 ( .A(n44797), .B(n37654), .Y(n18109) );
  NOR2X1 U16713 ( .A(n44800), .B(n37625), .Y(n18111) );
  NOR2X1 U16716 ( .A(n44797), .B(n37653), .Y(n18116) );
  NOR2X1 U16720 ( .A(n44800), .B(n37624), .Y(n18118) );
  NOR2X1 U16723 ( .A(n44797), .B(n37652), .Y(n18123) );
  NOR2X1 U16727 ( .A(n44800), .B(n37623), .Y(n18125) );
  NOR2X1 U16730 ( .A(n44797), .B(n37651), .Y(n18130) );
  NOR2X1 U16734 ( .A(n44800), .B(n37622), .Y(n18132) );
  NOR2X1 U16737 ( .A(n44797), .B(n37650), .Y(n18137) );
  NOR2X1 U16741 ( .A(n44800), .B(n37621), .Y(n18139) );
  NOR2X1 U16744 ( .A(n44797), .B(n37649), .Y(n18144) );
  NOR2X1 U16748 ( .A(n44800), .B(n37620), .Y(n18146) );
  NOR2X1 U16751 ( .A(n44797), .B(n37648), .Y(n18151) );
  NOR2X1 U16755 ( .A(n44800), .B(n37619), .Y(n18153) );
  NOR2X1 U16758 ( .A(n44797), .B(n37647), .Y(n18158) );
  NOR2X1 U16762 ( .A(n44800), .B(n37618), .Y(n18160) );
  NOR2X1 U16765 ( .A(n44797), .B(n37602), .Y(n18165) );
  NOR2X1 U16769 ( .A(n44800), .B(n37599), .Y(n18167) );
  NOR2X1 U16772 ( .A(n44798), .B(n37646), .Y(n18172) );
  NOR2X1 U16776 ( .A(n44801), .B(n37617), .Y(n18174) );
  NOR2X1 U16779 ( .A(n44798), .B(n37645), .Y(n18179) );
  NOR2X1 U16783 ( .A(n44801), .B(n37616), .Y(n18181) );
  NOR2X1 U16786 ( .A(n44798), .B(n37644), .Y(n18186) );
  NOR2X1 U16790 ( .A(n44801), .B(n37615), .Y(n18188) );
  NOR2X1 U16793 ( .A(n44798), .B(n37643), .Y(n18193) );
  NOR2X1 U16797 ( .A(n44801), .B(n37614), .Y(n18195) );
  NOR2X1 U16800 ( .A(n44798), .B(n37642), .Y(n18200) );
  NOR2X1 U16804 ( .A(n44801), .B(n37613), .Y(n18202) );
  NOR2X1 U16807 ( .A(n44798), .B(n37641), .Y(n18207) );
  NOR2X1 U16811 ( .A(n44801), .B(n37612), .Y(n18209) );
  NOR2X1 U16814 ( .A(n44798), .B(n37640), .Y(n18214) );
  NOR2X1 U16818 ( .A(n44801), .B(n37611), .Y(n18216) );
  NOR2X1 U16821 ( .A(n44798), .B(n37639), .Y(n18221) );
  NOR2X1 U16825 ( .A(n44801), .B(n37610), .Y(n18223) );
  NOR2X1 U16828 ( .A(n37638), .B(n44798), .Y(n18228) );
  NOR2X1 U16832 ( .A(n37609), .B(n44801), .Y(n18229) );
  NOR2X1 U16835 ( .A(n37637), .B(n44798), .Y(n18234) );
  NOR2X1 U16839 ( .A(n37608), .B(n44801), .Y(n18235) );
  NOR2X1 U16842 ( .A(n37636), .B(n44798), .Y(n18240) );
  NOR2X1 U16846 ( .A(n37607), .B(n44801), .Y(n18241) );
  NOR2X1 U16849 ( .A(n37635), .B(n44798), .Y(n18246) );
  NOR2X1 U16853 ( .A(n37606), .B(n44801), .Y(n18247) );
  NOR2X1 U16856 ( .A(n37634), .B(n44798), .Y(n18252) );
  NOR2X1 U16860 ( .A(n37605), .B(n44801), .Y(n18253) );
  NOR2X1 U16863 ( .A(n37662), .B(n44799), .Y(n18258) );
  NOR2X1 U16867 ( .A(n37633), .B(n44802), .Y(n18259) );
  NOR2X1 U16870 ( .A(n37661), .B(n44799), .Y(n18264) );
  NOR2X1 U16874 ( .A(n37632), .B(n44802), .Y(n18265) );
  NOR2X1 U16877 ( .A(n37660), .B(n44799), .Y(n18270) );
  NOR2X1 U16881 ( .A(n37631), .B(n44802), .Y(n18271) );
  NOR2X1 U16884 ( .A(n37659), .B(n44799), .Y(n18276) );
  NOR2X1 U16888 ( .A(n37630), .B(n44802), .Y(n18277) );
  NOR2X1 U16891 ( .A(n37658), .B(n44799), .Y(n18282) );
  NOR2X1 U16895 ( .A(n37629), .B(n44802), .Y(n18283) );
  NOR2X1 U16898 ( .A(n37604), .B(n44799), .Y(n18288) );
  NOR2X1 U16902 ( .A(n37601), .B(n44802), .Y(n18289) );
  NOR2X1 U16905 ( .A(n37603), .B(n44799), .Y(n18294) );
  NOR2X1 U16910 ( .A(n37600), .B(n44802), .Y(n18297) );
  NOR2X1 U16913 ( .A(n37657), .B(n44595), .Y(n18303) );
  NOR2X1 U16917 ( .A(n37628), .B(n44586), .Y(n18306) );
  NOR2X1 U16920 ( .A(n37656), .B(n44595), .Y(n18313) );
  NOR2X1 U16924 ( .A(n37627), .B(n44586), .Y(n18314) );
  NOR2X1 U16927 ( .A(n37655), .B(n44595), .Y(n18319) );
  NOR2X1 U16931 ( .A(n37626), .B(n44586), .Y(n18320) );
  NOR2X1 U16934 ( .A(n37654), .B(n44595), .Y(n18325) );
  NOR2X1 U16938 ( .A(n37625), .B(n44586), .Y(n18326) );
  NOR2X1 U16941 ( .A(n37653), .B(n44595), .Y(n18331) );
  NOR2X1 U16945 ( .A(n37624), .B(n44586), .Y(n18332) );
  NOR2X1 U16948 ( .A(n37652), .B(n44595), .Y(n18337) );
  NOR2X1 U16952 ( .A(n37623), .B(n44586), .Y(n18338) );
  NOR2X1 U16955 ( .A(n37651), .B(n44595), .Y(n18343) );
  NOR2X1 U16959 ( .A(n37622), .B(n44586), .Y(n18344) );
  NOR2X1 U16962 ( .A(n37650), .B(n44595), .Y(n18349) );
  NOR2X1 U16966 ( .A(n37621), .B(n44586), .Y(n18350) );
  NOR2X1 U16969 ( .A(n37649), .B(n44595), .Y(n18355) );
  NOR2X1 U16973 ( .A(n37620), .B(n44586), .Y(n18356) );
  NOR2X1 U16976 ( .A(n37648), .B(n44595), .Y(n18361) );
  NOR2X1 U16980 ( .A(n37619), .B(n44586), .Y(n18362) );
  NOR2X1 U16983 ( .A(n37647), .B(n44595), .Y(n18367) );
  NOR2X1 U16987 ( .A(n37618), .B(n44586), .Y(n18368) );
  NOR2X1 U16990 ( .A(n37602), .B(n44595), .Y(n18373) );
  NOR2X1 U16994 ( .A(n37599), .B(n44586), .Y(n18374) );
  NOR2X1 U16997 ( .A(n37646), .B(n44596), .Y(n18379) );
  NOR2X1 U17001 ( .A(n37617), .B(n44587), .Y(n18380) );
  NOR2X1 U17004 ( .A(n37645), .B(n44596), .Y(n18385) );
  NOR2X1 U17008 ( .A(n37616), .B(n44587), .Y(n18386) );
  NOR2X1 U17011 ( .A(n37644), .B(n44596), .Y(n18391) );
  NOR2X1 U17015 ( .A(n37615), .B(n44587), .Y(n18392) );
  NOR2X1 U17018 ( .A(n37643), .B(n44596), .Y(n18397) );
  NOR2X1 U17022 ( .A(n37614), .B(n44587), .Y(n18398) );
  NOR2X1 U17025 ( .A(n37642), .B(n44596), .Y(n18403) );
  NOR2X1 U17029 ( .A(n37613), .B(n44587), .Y(n18404) );
  NOR2X1 U17032 ( .A(n37641), .B(n44596), .Y(n18409) );
  NOR2X1 U17036 ( .A(n37612), .B(n44587), .Y(n18410) );
  NOR2X1 U17039 ( .A(n37640), .B(n44596), .Y(n18415) );
  NOR2X1 U17043 ( .A(n37611), .B(n44587), .Y(n18416) );
  NOR2X1 U17046 ( .A(n37639), .B(n44596), .Y(n18421) );
  NOR2X1 U17050 ( .A(n37610), .B(n44587), .Y(n18422) );
  NOR2X1 U17053 ( .A(n37638), .B(n44596), .Y(n18427) );
  NOR2X1 U17057 ( .A(n37609), .B(n44587), .Y(n18428) );
  NOR2X1 U17060 ( .A(n37637), .B(n44596), .Y(n18433) );
  NOR2X1 U17064 ( .A(n37608), .B(n44587), .Y(n18434) );
  NOR2X1 U17067 ( .A(n37636), .B(n44596), .Y(n18439) );
  NOR2X1 U17071 ( .A(n37607), .B(n44587), .Y(n18440) );
  NOR2X1 U17074 ( .A(n37635), .B(n44596), .Y(n18445) );
  NOR2X1 U17078 ( .A(n37606), .B(n44587), .Y(n18446) );
  NOR2X1 U17081 ( .A(n37634), .B(n44597), .Y(n18451) );
  NOR2X1 U17085 ( .A(n37605), .B(n44588), .Y(n18452) );
  NOR2X1 U17088 ( .A(n37662), .B(n44597), .Y(n18457) );
  NOR2X1 U17092 ( .A(n37633), .B(n44588), .Y(n18458) );
  NOR2X1 U17095 ( .A(n37661), .B(n44597), .Y(n18463) );
  NOR2X1 U17099 ( .A(n37632), .B(n44588), .Y(n18464) );
  NOR2X1 U17102 ( .A(n37660), .B(n44597), .Y(n18469) );
  NOR2X1 U17106 ( .A(n37631), .B(n44588), .Y(n18470) );
  NOR2X1 U17109 ( .A(n37659), .B(n44597), .Y(n18475) );
  NOR2X1 U17113 ( .A(n37630), .B(n44588), .Y(n18476) );
  NOR2X1 U17116 ( .A(n37658), .B(n44597), .Y(n18481) );
  NOR2X1 U17120 ( .A(n37629), .B(n44588), .Y(n18482) );
  NOR2X1 U17123 ( .A(n37604), .B(n44597), .Y(n18487) );
  NOR2X1 U17127 ( .A(n37601), .B(n44588), .Y(n18488) );
  NOR2X1 U17130 ( .A(n37603), .B(n44597), .Y(n18493) );
  NAND2X1 U17132 ( .A(n563), .B(n44591), .Y(n18305) );
  NOR2X1 U17135 ( .A(n37600), .B(n44588), .Y(n18494) );
  NOR2X1 U17138 ( .A(n37657), .B(n44785), .Y(n18499) );
  NOR2X1 U17142 ( .A(n37628), .B(n44788), .Y(n18501) );
  NOR2X1 U17145 ( .A(n37656), .B(n44785), .Y(n18507) );
  NOR2X1 U17149 ( .A(n37627), .B(n44788), .Y(n18508) );
  NOR2X1 U17152 ( .A(n37655), .B(n44785), .Y(n18513) );
  NOR2X1 U17156 ( .A(n37626), .B(n44788), .Y(n18514) );
  NOR2X1 U17159 ( .A(n37654), .B(n44785), .Y(n18519) );
  NOR2X1 U17163 ( .A(n37625), .B(n44788), .Y(n18520) );
  NOR2X1 U17166 ( .A(n37653), .B(n44785), .Y(n18525) );
  NOR2X1 U17170 ( .A(n37624), .B(n44788), .Y(n18526) );
  NOR2X1 U17173 ( .A(n37652), .B(n44785), .Y(n18531) );
  NOR2X1 U17177 ( .A(n37623), .B(n44788), .Y(n18532) );
  NOR2X1 U17180 ( .A(n37651), .B(n44785), .Y(n18537) );
  NOR2X1 U17184 ( .A(n37622), .B(n44788), .Y(n18538) );
  NOR2X1 U17187 ( .A(n37650), .B(n44785), .Y(n18543) );
  NOR2X1 U17191 ( .A(n37621), .B(n44788), .Y(n18544) );
  NOR2X1 U17194 ( .A(n37649), .B(n44785), .Y(n18549) );
  NOR2X1 U17198 ( .A(n37620), .B(n44788), .Y(n18550) );
  NOR2X1 U17201 ( .A(n37648), .B(n44785), .Y(n18555) );
  NOR2X1 U17205 ( .A(n37619), .B(n44788), .Y(n18556) );
  NOR2X1 U17208 ( .A(n37647), .B(n44785), .Y(n18561) );
  NOR2X1 U17212 ( .A(n37618), .B(n44788), .Y(n18562) );
  NOR2X1 U17215 ( .A(n37602), .B(n44785), .Y(n18567) );
  NOR2X1 U17219 ( .A(n37599), .B(n44788), .Y(n18568) );
  NOR2X1 U17222 ( .A(n37646), .B(n44786), .Y(n18573) );
  NOR2X1 U17226 ( .A(n37617), .B(n44789), .Y(n18574) );
  NOR2X1 U17229 ( .A(n37645), .B(n44786), .Y(n18579) );
  NOR2X1 U17233 ( .A(n37616), .B(n44789), .Y(n18580) );
  NOR2X1 U17236 ( .A(n37644), .B(n44786), .Y(n18585) );
  NOR2X1 U17240 ( .A(n37615), .B(n44789), .Y(n18586) );
  NOR2X1 U17243 ( .A(n37643), .B(n44786), .Y(n18591) );
  NOR2X1 U17247 ( .A(n37614), .B(n44789), .Y(n18592) );
  NOR2X1 U17250 ( .A(n37642), .B(n44786), .Y(n18597) );
  NOR2X1 U17254 ( .A(n37613), .B(n44789), .Y(n18598) );
  NOR2X1 U17257 ( .A(n37641), .B(n44786), .Y(n18603) );
  NOR2X1 U17261 ( .A(n37612), .B(n44789), .Y(n18604) );
  NOR2X1 U17264 ( .A(n37640), .B(n44786), .Y(n18609) );
  NOR2X1 U17268 ( .A(n37611), .B(n44789), .Y(n18610) );
  NOR2X1 U17271 ( .A(n37639), .B(n44786), .Y(n18615) );
  NOR2X1 U17275 ( .A(n37610), .B(n44789), .Y(n18616) );
  NOR2X1 U17278 ( .A(n37638), .B(n44786), .Y(n18621) );
  NOR2X1 U17282 ( .A(n37609), .B(n44789), .Y(n18622) );
  NOR2X1 U17285 ( .A(n37637), .B(n44786), .Y(n18627) );
  NOR2X1 U17289 ( .A(n37608), .B(n44789), .Y(n18628) );
  NOR2X1 U17292 ( .A(n37636), .B(n44786), .Y(n18633) );
  NOR2X1 U17296 ( .A(n37607), .B(n44789), .Y(n18634) );
  NOR2X1 U17299 ( .A(n37635), .B(n44786), .Y(n18639) );
  NOR2X1 U17303 ( .A(n37606), .B(n44789), .Y(n18640) );
  NOR2X1 U17306 ( .A(n37634), .B(n44787), .Y(n18645) );
  NOR2X1 U17310 ( .A(n37605), .B(n44790), .Y(n18646) );
  NOR2X1 U17313 ( .A(n37662), .B(n44787), .Y(n18651) );
  NOR2X1 U17317 ( .A(n37633), .B(n44790), .Y(n18652) );
  NOR2X1 U17320 ( .A(n37661), .B(n44787), .Y(n18657) );
  NOR2X1 U17324 ( .A(n37632), .B(n44790), .Y(n18658) );
  NOR2X1 U17327 ( .A(n37660), .B(n44787), .Y(n18663) );
  NOR2X1 U17331 ( .A(n37631), .B(n44790), .Y(n18664) );
  NOR2X1 U17334 ( .A(n37659), .B(n44787), .Y(n18669) );
  NOR2X1 U17338 ( .A(n37630), .B(n44790), .Y(n18670) );
  NOR2X1 U17341 ( .A(n37658), .B(n44787), .Y(n18675) );
  NOR2X1 U17345 ( .A(n37629), .B(n44790), .Y(n18676) );
  NOR2X1 U17348 ( .A(n37604), .B(n44787), .Y(n18681) );
  NOR2X1 U17352 ( .A(n37601), .B(n44790), .Y(n18682) );
  NOR2X1 U17355 ( .A(n37603), .B(n44787), .Y(n18687) );
  NOR2X1 U17360 ( .A(n37600), .B(n44790), .Y(n18689) );
  NOR2X1 U17363 ( .A(n37657), .B(n44775), .Y(n18695) );
  NOR2X1 U17367 ( .A(n37628), .B(n44778), .Y(n18697) );
  NOR2X1 U17370 ( .A(n37656), .B(n44775), .Y(n18703) );
  NOR2X1 U17374 ( .A(n37627), .B(n44778), .Y(n18704) );
  NOR2X1 U17377 ( .A(n37655), .B(n44775), .Y(n18709) );
  NOR2X1 U17381 ( .A(n37626), .B(n44778), .Y(n18710) );
  NOR2X1 U17384 ( .A(n37654), .B(n44775), .Y(n18715) );
  NOR2X1 U17388 ( .A(n37625), .B(n44778), .Y(n18716) );
  NOR2X1 U17391 ( .A(n37653), .B(n44775), .Y(n18721) );
  NOR2X1 U17395 ( .A(n37624), .B(n44778), .Y(n18722) );
  NOR2X1 U17398 ( .A(n37652), .B(n44775), .Y(n18727) );
  NOR2X1 U17402 ( .A(n37623), .B(n44778), .Y(n18728) );
  NOR2X1 U17405 ( .A(n37651), .B(n44775), .Y(n18733) );
  NOR2X1 U17409 ( .A(n37622), .B(n44778), .Y(n18734) );
  NOR2X1 U17412 ( .A(n37650), .B(n44775), .Y(n18739) );
  NOR2X1 U17416 ( .A(n37621), .B(n44778), .Y(n18740) );
  NOR2X1 U17419 ( .A(n37649), .B(n44775), .Y(n18745) );
  NOR2X1 U17423 ( .A(n37620), .B(n44778), .Y(n18746) );
  NOR2X1 U17426 ( .A(n37648), .B(n44775), .Y(n18751) );
  NOR2X1 U17430 ( .A(n37619), .B(n44778), .Y(n18752) );
  NOR2X1 U17433 ( .A(n37647), .B(n44775), .Y(n18757) );
  NOR2X1 U17437 ( .A(n37618), .B(n44778), .Y(n18758) );
  NOR2X1 U17440 ( .A(n37602), .B(n44775), .Y(n18763) );
  NOR2X1 U17444 ( .A(n37599), .B(n44778), .Y(n18764) );
  NOR2X1 U17447 ( .A(n37646), .B(n44776), .Y(n18769) );
  NOR2X1 U17451 ( .A(n37617), .B(n44779), .Y(n18770) );
  NOR2X1 U17454 ( .A(n37645), .B(n44776), .Y(n18775) );
  NOR2X1 U17458 ( .A(n37616), .B(n44779), .Y(n18776) );
  NOR2X1 U17461 ( .A(n37644), .B(n44776), .Y(n18781) );
  NOR2X1 U17465 ( .A(n37615), .B(n44779), .Y(n18782) );
  NOR2X1 U17468 ( .A(n37643), .B(n44776), .Y(n18787) );
  NOR2X1 U17472 ( .A(n37614), .B(n44779), .Y(n18788) );
  NOR2X1 U17475 ( .A(n37642), .B(n44776), .Y(n18793) );
  NOR2X1 U17479 ( .A(n37613), .B(n44779), .Y(n18794) );
  NOR2X1 U17482 ( .A(n37641), .B(n44776), .Y(n18799) );
  NOR2X1 U17486 ( .A(n37612), .B(n44779), .Y(n18800) );
  NOR2X1 U17489 ( .A(n37640), .B(n44776), .Y(n18805) );
  NOR2X1 U17493 ( .A(n37611), .B(n44779), .Y(n18806) );
  NOR2X1 U17496 ( .A(n37639), .B(n44776), .Y(n18811) );
  NOR2X1 U17500 ( .A(n37610), .B(n44779), .Y(n18812) );
  NOR2X1 U17503 ( .A(n37638), .B(n44776), .Y(n18817) );
  NOR2X1 U17507 ( .A(n37609), .B(n44779), .Y(n18818) );
  NOR2X1 U17510 ( .A(n37637), .B(n44776), .Y(n18823) );
  NOR2X1 U17514 ( .A(n37608), .B(n44779), .Y(n18824) );
  NOR2X1 U17517 ( .A(n37636), .B(n44776), .Y(n18829) );
  NOR2X1 U17521 ( .A(n37607), .B(n44779), .Y(n18830) );
  NOR2X1 U17524 ( .A(n37635), .B(n44776), .Y(n18835) );
  NOR2X1 U17528 ( .A(n37606), .B(n44779), .Y(n18836) );
  NOR2X1 U17531 ( .A(n37634), .B(n44777), .Y(n18841) );
  NOR2X1 U17535 ( .A(n37605), .B(n44780), .Y(n18842) );
  NOR2X1 U17538 ( .A(n37662), .B(n44777), .Y(n18847) );
  NOR2X1 U17542 ( .A(n37633), .B(n44780), .Y(n18848) );
  NOR2X1 U17545 ( .A(n37661), .B(n44777), .Y(n18853) );
  NOR2X1 U17549 ( .A(n37632), .B(n44780), .Y(n18854) );
  NOR2X1 U17552 ( .A(n37660), .B(n44777), .Y(n18859) );
  NOR2X1 U17556 ( .A(n37631), .B(n44780), .Y(n18860) );
  NOR2X1 U17559 ( .A(n37659), .B(n44777), .Y(n18865) );
  NOR2X1 U17563 ( .A(n37630), .B(n44780), .Y(n18866) );
  NOR2X1 U17566 ( .A(n37658), .B(n44777), .Y(n18871) );
  NOR2X1 U17570 ( .A(n37629), .B(n44780), .Y(n18872) );
  NOR2X1 U17573 ( .A(n37604), .B(n44777), .Y(n18877) );
  NOR2X1 U17577 ( .A(n37601), .B(n44780), .Y(n18878) );
  NOR2X1 U17580 ( .A(n37603), .B(n44777), .Y(n18883) );
  NAND2X1 U17582 ( .A(n555), .B(n44576), .Y(n18696) );
  NOR2X1 U17585 ( .A(n37600), .B(n44780), .Y(n18885) );
  NOR2X1 U17588 ( .A(n37657), .B(n44791), .Y(n18891) );
  NOR2X1 U17592 ( .A(n37628), .B(n44794), .Y(n18893) );
  NOR2X1 U17595 ( .A(n37656), .B(n44791), .Y(n18899) );
  NOR2X1 U17599 ( .A(n37627), .B(n44794), .Y(n18900) );
  NOR2X1 U17602 ( .A(n37655), .B(n44791), .Y(n18905) );
  NOR2X1 U17606 ( .A(n37626), .B(n44794), .Y(n18906) );
  NOR2X1 U17609 ( .A(n37654), .B(n44791), .Y(n18911) );
  NOR2X1 U17613 ( .A(n37625), .B(n44794), .Y(n18912) );
  NOR2X1 U17616 ( .A(n37653), .B(n44791), .Y(n18917) );
  NOR2X1 U17620 ( .A(n37624), .B(n44794), .Y(n18918) );
  NOR2X1 U17623 ( .A(n37652), .B(n44791), .Y(n18923) );
  NOR2X1 U17627 ( .A(n37623), .B(n44794), .Y(n18924) );
  NOR2X1 U17630 ( .A(n37651), .B(n44791), .Y(n18929) );
  NOR2X1 U17634 ( .A(n37622), .B(n44794), .Y(n18930) );
  NOR2X1 U17637 ( .A(n37650), .B(n44791), .Y(n18935) );
  NOR2X1 U17641 ( .A(n37621), .B(n44794), .Y(n18936) );
  NOR2X1 U17644 ( .A(n37649), .B(n44791), .Y(n18941) );
  NOR2X1 U17648 ( .A(n37620), .B(n44794), .Y(n18942) );
  NOR2X1 U17651 ( .A(n37648), .B(n44791), .Y(n18947) );
  NOR2X1 U17655 ( .A(n37619), .B(n44794), .Y(n18948) );
  NOR2X1 U17658 ( .A(n37647), .B(n44791), .Y(n18953) );
  NOR2X1 U17662 ( .A(n37618), .B(n44794), .Y(n18954) );
  NOR2X1 U17665 ( .A(n37602), .B(n44791), .Y(n18959) );
  NOR2X1 U17669 ( .A(n37599), .B(n44794), .Y(n18960) );
  NOR2X1 U17672 ( .A(n37646), .B(n44792), .Y(n18965) );
  NOR2X1 U17676 ( .A(n37617), .B(n44795), .Y(n18966) );
  NOR2X1 U17679 ( .A(n37645), .B(n44792), .Y(n18971) );
  NOR2X1 U17683 ( .A(n37616), .B(n44795), .Y(n18972) );
  NOR2X1 U17686 ( .A(n37644), .B(n44792), .Y(n18977) );
  NOR2X1 U17690 ( .A(n37615), .B(n44795), .Y(n18978) );
  NOR2X1 U17693 ( .A(n37643), .B(n44792), .Y(n18983) );
  NOR2X1 U17697 ( .A(n37614), .B(n44795), .Y(n18984) );
  NOR2X1 U17700 ( .A(n37642), .B(n44792), .Y(n18989) );
  NOR2X1 U17704 ( .A(n37613), .B(n44795), .Y(n18990) );
  NOR2X1 U17707 ( .A(n37641), .B(n44792), .Y(n18995) );
  NOR2X1 U17711 ( .A(n37612), .B(n44795), .Y(n18996) );
  NOR2X1 U17714 ( .A(n37640), .B(n44792), .Y(n19001) );
  NOR2X1 U17718 ( .A(n37611), .B(n44795), .Y(n19002) );
  NOR2X1 U17721 ( .A(n37639), .B(n44792), .Y(n19007) );
  NOR2X1 U17725 ( .A(n37610), .B(n44795), .Y(n19008) );
  NOR2X1 U17728 ( .A(n37638), .B(n44792), .Y(n19013) );
  NOR2X1 U17732 ( .A(n37609), .B(n44795), .Y(n19014) );
  NOR2X1 U17735 ( .A(n37637), .B(n44792), .Y(n19019) );
  NOR2X1 U17739 ( .A(n37608), .B(n44795), .Y(n19020) );
  NOR2X1 U17742 ( .A(n37636), .B(n44792), .Y(n19025) );
  NOR2X1 U17746 ( .A(n37607), .B(n44795), .Y(n19026) );
  NOR2X1 U17749 ( .A(n37635), .B(n44792), .Y(n19031) );
  NOR2X1 U17753 ( .A(n37606), .B(n44795), .Y(n19032) );
  NOR2X1 U17756 ( .A(n37634), .B(n44793), .Y(n19037) );
  NOR2X1 U17760 ( .A(n37605), .B(n44796), .Y(n19038) );
  NOR2X1 U17763 ( .A(n37662), .B(n44793), .Y(n19043) );
  NOR2X1 U17767 ( .A(n37633), .B(n44796), .Y(n19044) );
  NOR2X1 U17770 ( .A(n37661), .B(n44793), .Y(n19049) );
  NOR2X1 U17774 ( .A(n37632), .B(n44796), .Y(n19050) );
  NOR2X1 U17777 ( .A(n37660), .B(n44793), .Y(n19055) );
  NOR2X1 U17781 ( .A(n37631), .B(n44796), .Y(n19056) );
  NOR2X1 U17784 ( .A(n37659), .B(n44793), .Y(n19061) );
  NOR2X1 U17788 ( .A(n37630), .B(n44796), .Y(n19062) );
  NOR2X1 U17791 ( .A(n37658), .B(n44793), .Y(n19067) );
  NOR2X1 U17795 ( .A(n37629), .B(n44796), .Y(n19068) );
  NOR2X1 U17798 ( .A(n37604), .B(n44793), .Y(n19073) );
  NOR2X1 U17802 ( .A(n37601), .B(n44796), .Y(n19074) );
  NOR2X1 U17805 ( .A(n37603), .B(n44793), .Y(n19079) );
  NOR2X1 U17810 ( .A(n37600), .B(n44796), .Y(n19081) );
  NOR2X1 U17813 ( .A(n37657), .B(n44769), .Y(n19087) );
  NOR2X1 U17817 ( .A(n37628), .B(n44772), .Y(n19089) );
  NOR2X1 U17820 ( .A(n37656), .B(n44769), .Y(n19095) );
  NOR2X1 U17824 ( .A(n37627), .B(n44772), .Y(n19096) );
  NOR2X1 U17827 ( .A(n37655), .B(n44769), .Y(n19101) );
  NOR2X1 U17831 ( .A(n37626), .B(n44772), .Y(n19102) );
  NOR2X1 U17834 ( .A(n37654), .B(n44769), .Y(n19107) );
  NOR2X1 U17838 ( .A(n37625), .B(n44772), .Y(n19108) );
  NOR2X1 U17841 ( .A(n37653), .B(n44769), .Y(n19113) );
  NOR2X1 U17845 ( .A(n37624), .B(n44772), .Y(n19114) );
  NOR2X1 U17848 ( .A(n37652), .B(n44769), .Y(n19119) );
  NOR2X1 U17852 ( .A(n37623), .B(n44772), .Y(n19120) );
  NOR2X1 U17855 ( .A(n37651), .B(n44769), .Y(n19125) );
  NOR2X1 U17859 ( .A(n37622), .B(n44772), .Y(n19126) );
  NOR2X1 U17862 ( .A(n37650), .B(n44769), .Y(n19131) );
  NOR2X1 U17866 ( .A(n37621), .B(n44772), .Y(n19132) );
  NOR2X1 U17869 ( .A(n37649), .B(n44769), .Y(n19137) );
  NOR2X1 U17873 ( .A(n37620), .B(n44772), .Y(n19138) );
  NOR2X1 U17876 ( .A(n37648), .B(n44769), .Y(n19143) );
  NOR2X1 U17880 ( .A(n37619), .B(n44772), .Y(n19144) );
  NOR2X1 U17883 ( .A(n37647), .B(n44769), .Y(n19149) );
  NOR2X1 U17887 ( .A(n37618), .B(n44772), .Y(n19150) );
  NOR2X1 U17890 ( .A(n37602), .B(n44769), .Y(n19155) );
  NOR2X1 U17894 ( .A(n37599), .B(n44772), .Y(n19156) );
  NOR2X1 U17897 ( .A(n37646), .B(n44770), .Y(n19161) );
  NOR2X1 U17901 ( .A(n37617), .B(n44773), .Y(n19162) );
  NOR2X1 U17904 ( .A(n37645), .B(n44770), .Y(n19167) );
  NOR2X1 U17908 ( .A(n37616), .B(n44773), .Y(n19168) );
  NOR2X1 U17911 ( .A(n37644), .B(n44770), .Y(n19173) );
  NOR2X1 U17915 ( .A(n37615), .B(n44773), .Y(n19174) );
  NOR2X1 U17918 ( .A(n37643), .B(n44770), .Y(n19179) );
  NOR2X1 U17922 ( .A(n37614), .B(n44773), .Y(n19180) );
  NOR2X1 U17925 ( .A(n37642), .B(n44770), .Y(n19185) );
  NOR2X1 U17929 ( .A(n37613), .B(n44773), .Y(n19186) );
  NOR2X1 U17932 ( .A(n37641), .B(n44770), .Y(n19191) );
  NOR2X1 U17936 ( .A(n37612), .B(n44773), .Y(n19192) );
  NOR2X1 U17939 ( .A(n37640), .B(n44770), .Y(n19197) );
  NOR2X1 U17943 ( .A(n37611), .B(n44773), .Y(n19198) );
  NOR2X1 U17946 ( .A(n37639), .B(n44770), .Y(n19203) );
  NOR2X1 U17950 ( .A(n37610), .B(n44773), .Y(n19204) );
  NOR2X1 U17953 ( .A(n37638), .B(n44770), .Y(n19209) );
  NOR2X1 U17957 ( .A(n37609), .B(n44773), .Y(n19210) );
  NOR2X1 U17960 ( .A(n37637), .B(n44770), .Y(n19215) );
  NOR2X1 U17964 ( .A(n37608), .B(n44773), .Y(n19216) );
  NOR2X1 U17967 ( .A(n37636), .B(n44770), .Y(n19221) );
  NOR2X1 U17971 ( .A(n37607), .B(n44773), .Y(n19222) );
  NOR2X1 U17974 ( .A(n37635), .B(n44770), .Y(n19227) );
  NOR2X1 U17978 ( .A(n37606), .B(n44773), .Y(n19228) );
  NOR2X1 U17981 ( .A(n37634), .B(n44771), .Y(n19233) );
  NOR2X1 U17985 ( .A(n37605), .B(n44774), .Y(n19234) );
  NOR2X1 U17988 ( .A(n37662), .B(n44771), .Y(n19239) );
  NOR2X1 U17992 ( .A(n37633), .B(n44774), .Y(n19240) );
  NOR2X1 U17995 ( .A(n37661), .B(n44771), .Y(n19245) );
  NOR2X1 U17999 ( .A(n37632), .B(n44774), .Y(n19246) );
  NOR2X1 U18002 ( .A(n37660), .B(n44771), .Y(n19251) );
  NOR2X1 U18006 ( .A(n37631), .B(n44774), .Y(n19252) );
  NOR2X1 U18009 ( .A(n37659), .B(n44771), .Y(n19257) );
  NOR2X1 U18013 ( .A(n37630), .B(n44774), .Y(n19258) );
  NOR2X1 U18016 ( .A(n37658), .B(n44771), .Y(n19263) );
  NOR2X1 U18020 ( .A(n37629), .B(n44774), .Y(n19264) );
  NOR2X1 U18023 ( .A(n37604), .B(n44771), .Y(n19269) );
  NOR2X1 U18027 ( .A(n37601), .B(n44774), .Y(n19270) );
  NOR2X1 U18030 ( .A(n37603), .B(n44771), .Y(n19275) );
  NAND2X1 U18032 ( .A(n559), .B(n44564), .Y(n19088) );
  NOR2X1 U18035 ( .A(n37600), .B(n44774), .Y(n19277) );
  NOR2X1 U18038 ( .A(n44680), .B(n44781), .Y(n19283) );
  NOR2X1 U18042 ( .A(n44708), .B(n44783), .Y(n19285) );
  NOR2X1 U18045 ( .A(n44642), .B(n44781), .Y(n19291) );
  NOR2X1 U18049 ( .A(n44706), .B(n44783), .Y(n19292) );
  NOR2X1 U18052 ( .A(n44648), .B(n44781), .Y(n19297) );
  NOR2X1 U18056 ( .A(n44714), .B(n44783), .Y(n19298) );
  NOR2X1 U18059 ( .A(n44650), .B(n44781), .Y(n19303) );
  NOR2X1 U18063 ( .A(n44716), .B(n44783), .Y(n19304) );
  NOR2X1 U18066 ( .A(n44672), .B(n44781), .Y(n19309) );
  NOR2X1 U18070 ( .A(n44738), .B(n44783), .Y(n19310) );
  NOR2X1 U18073 ( .A(n44664), .B(n44781), .Y(n19315) );
  NOR2X1 U18077 ( .A(n44730), .B(n44783), .Y(n19316) );
  NOR2X1 U18080 ( .A(n44674), .B(n44781), .Y(n19321) );
  NOR2X1 U18084 ( .A(n44740), .B(n44783), .Y(n19322) );
  NOR2X1 U18087 ( .A(n44676), .B(n44781), .Y(n19327) );
  NOR2X1 U18091 ( .A(n44742), .B(n44783), .Y(n19328) );
  NOR2X1 U18094 ( .A(n44656), .B(n44781), .Y(n19333) );
  NOR2X1 U18098 ( .A(n44722), .B(n44783), .Y(n19334) );
  NOR2X1 U18101 ( .A(n44658), .B(n44781), .Y(n19339) );
  NOR2X1 U18105 ( .A(n44724), .B(n44783), .Y(n19340) );
  NOR2X1 U18108 ( .A(n44662), .B(n44781), .Y(n19345) );
  NOR2X1 U18112 ( .A(n44728), .B(n44783), .Y(n19346) );
  NOR2X1 U18115 ( .A(n44654), .B(n44781), .Y(n19351) );
  NOR2X1 U18119 ( .A(n44720), .B(n44783), .Y(n19352) );
  NOR2X1 U18122 ( .A(n44652), .B(n44782), .Y(n19357) );
  NOR2X1 U18126 ( .A(n44718), .B(n44784), .Y(n19358) );
  NOR2X1 U18129 ( .A(n44666), .B(n44782), .Y(n19363) );
  NOR2X1 U18133 ( .A(n44732), .B(n44784), .Y(n19364) );
  NOR2X1 U18136 ( .A(n44678), .B(n44782), .Y(n19369) );
  NOR2X1 U18140 ( .A(n44744), .B(n44784), .Y(n19370) );
  NOR2X1 U18143 ( .A(n44660), .B(n44782), .Y(n19375) );
  NOR2X1 U18147 ( .A(n44726), .B(n44784), .Y(n19376) );
  NOR2X1 U18150 ( .A(n44644), .B(n44782), .Y(n19381) );
  NOR2X1 U18154 ( .A(n44710), .B(n44784), .Y(n19382) );
  NOR2X1 U18157 ( .A(n44646), .B(n44782), .Y(n19387) );
  NOR2X1 U18161 ( .A(n44712), .B(n44784), .Y(n19388) );
  NOR2X1 U18164 ( .A(n44670), .B(n44782), .Y(n19393) );
  NOR2X1 U18168 ( .A(n44736), .B(n44784), .Y(n19394) );
  NOR2X1 U18171 ( .A(n44668), .B(n44782), .Y(n19399) );
  NOR2X1 U18175 ( .A(n44734), .B(n44784), .Y(n19400) );
  NOR2X1 U18178 ( .A(n44694), .B(n44782), .Y(n19405) );
  NOR2X1 U18182 ( .A(n44758), .B(n44784), .Y(n19406) );
  NOR2X1 U18185 ( .A(n44698), .B(n44782), .Y(n19411) );
  NOR2X1 U18189 ( .A(n44762), .B(n44784), .Y(n19412) );
  NOR2X1 U18192 ( .A(n44700), .B(n44782), .Y(n19417) );
  NOR2X1 U18196 ( .A(n44764), .B(n44784), .Y(n19418) );
  NOR2X1 U18199 ( .A(n44704), .B(n44782), .Y(n19423) );
  NOR2X1 U18203 ( .A(n44768), .B(n44784), .Y(n19424) );
  NOR2X1 U18206 ( .A(n44702), .B(n541), .Y(n19429) );
  NOR2X1 U18210 ( .A(n44766), .B(n540), .Y(n19430) );
  NOR2X1 U18213 ( .A(n44696), .B(n541), .Y(n19435) );
  NOR2X1 U18217 ( .A(n44760), .B(n540), .Y(n19436) );
  NOR2X1 U18220 ( .A(n44692), .B(n541), .Y(n19441) );
  NOR2X1 U18224 ( .A(n44748), .B(n540), .Y(n19442) );
  NOR2X1 U18227 ( .A(n44690), .B(n541), .Y(n19447) );
  NOR2X1 U18231 ( .A(n44752), .B(n540), .Y(n19448) );
  NOR2X1 U18234 ( .A(n44688), .B(n541), .Y(n19453) );
  NOR2X1 U18238 ( .A(n44754), .B(n540), .Y(n19454) );
  NOR2X1 U18241 ( .A(n44686), .B(n541), .Y(n19459) );
  NOR2X1 U18245 ( .A(n44756), .B(n540), .Y(n19460) );
  NOR2X1 U18248 ( .A(n44684), .B(n541), .Y(n19465) );
  NOR2X1 U18252 ( .A(n44750), .B(n540), .Y(n19466) );
  NOR2X1 U18255 ( .A(n44682), .B(n541), .Y(n19471) );
  NOR2X1 U18260 ( .A(n44746), .B(n540), .Y(n19473) );
  NOR2X1 U18263 ( .A(n44680), .B(n44553), .Y(n19479) );
  NOR2X1 U18267 ( .A(n44708), .B(n44544), .Y(n19482) );
  NOR2X1 U18270 ( .A(n44642), .B(n44553), .Y(n19489) );
  NOR2X1 U18274 ( .A(n44706), .B(n44544), .Y(n19490) );
  NOR2X1 U18277 ( .A(n44648), .B(n44553), .Y(n19495) );
  NOR2X1 U18281 ( .A(n44714), .B(n44544), .Y(n19496) );
  NOR2X1 U18284 ( .A(n44650), .B(n44553), .Y(n19501) );
  NOR2X1 U18288 ( .A(n44716), .B(n44544), .Y(n19502) );
  NOR2X1 U18291 ( .A(n44672), .B(n44553), .Y(n19507) );
  NOR2X1 U18295 ( .A(n44738), .B(n44544), .Y(n19508) );
  NOR2X1 U18298 ( .A(n44664), .B(n44553), .Y(n19513) );
  NOR2X1 U18302 ( .A(n44730), .B(n44544), .Y(n19514) );
  NOR2X1 U18305 ( .A(n44674), .B(n44553), .Y(n19519) );
  NOR2X1 U18309 ( .A(n44740), .B(n44544), .Y(n19520) );
  NOR2X1 U18312 ( .A(n44676), .B(n44553), .Y(n19525) );
  NOR2X1 U18316 ( .A(n44742), .B(n44544), .Y(n19526) );
  NOR2X1 U18319 ( .A(n44656), .B(n44553), .Y(n19531) );
  NOR2X1 U18323 ( .A(n44722), .B(n44544), .Y(n19532) );
  NOR2X1 U18326 ( .A(n44658), .B(n44553), .Y(n19537) );
  NOR2X1 U18330 ( .A(n44724), .B(n44544), .Y(n19538) );
  NOR2X1 U18333 ( .A(n44662), .B(n44553), .Y(n19543) );
  NOR2X1 U18337 ( .A(n44728), .B(n44544), .Y(n19544) );
  NOR2X1 U18340 ( .A(n44654), .B(n44553), .Y(n19549) );
  NOR2X1 U18344 ( .A(n44720), .B(n44544), .Y(n19550) );
  NOR2X1 U18347 ( .A(n44652), .B(n44554), .Y(n19555) );
  NOR2X1 U18351 ( .A(n44718), .B(n44545), .Y(n19556) );
  NOR2X1 U18354 ( .A(n44666), .B(n44554), .Y(n19561) );
  NOR2X1 U18358 ( .A(n44732), .B(n44545), .Y(n19562) );
  NOR2X1 U18361 ( .A(n44678), .B(n44554), .Y(n19567) );
  NOR2X1 U18365 ( .A(n44744), .B(n44545), .Y(n19568) );
  NOR2X1 U18368 ( .A(n44660), .B(n44554), .Y(n19573) );
  NOR2X1 U18372 ( .A(n44726), .B(n44545), .Y(n19574) );
  NOR2X1 U18375 ( .A(n44644), .B(n44554), .Y(n19579) );
  NOR2X1 U18379 ( .A(n44710), .B(n44545), .Y(n19580) );
  NOR2X1 U18382 ( .A(n44646), .B(n44554), .Y(n19585) );
  NOR2X1 U18386 ( .A(n44712), .B(n44545), .Y(n19586) );
  NOR2X1 U18389 ( .A(n44670), .B(n44554), .Y(n19591) );
  NOR2X1 U18393 ( .A(n44736), .B(n44545), .Y(n19592) );
  NOR2X1 U18396 ( .A(n44668), .B(n44554), .Y(n19597) );
  NOR2X1 U18400 ( .A(n44734), .B(n44545), .Y(n19598) );
  NOR2X1 U18403 ( .A(n44694), .B(n44554), .Y(n19603) );
  NOR2X1 U18407 ( .A(n44758), .B(n44545), .Y(n19604) );
  NOR2X1 U18410 ( .A(n44698), .B(n44554), .Y(n19609) );
  NOR2X1 U18414 ( .A(n44762), .B(n44545), .Y(n19610) );
  NOR2X1 U18417 ( .A(n44700), .B(n44554), .Y(n19615) );
  NOR2X1 U18421 ( .A(n44764), .B(n44545), .Y(n19616) );
  NOR2X1 U18424 ( .A(n44704), .B(n44554), .Y(n19621) );
  NOR2X1 U18428 ( .A(n44768), .B(n44545), .Y(n19622) );
  NOR2X1 U18431 ( .A(n44702), .B(n44555), .Y(n19627) );
  NOR2X1 U18435 ( .A(n44766), .B(n44546), .Y(n19628) );
  NOR2X1 U18438 ( .A(n44696), .B(n44555), .Y(n19633) );
  NOR2X1 U18442 ( .A(n44760), .B(n44546), .Y(n19634) );
  NOR2X1 U18445 ( .A(n44692), .B(n44555), .Y(n19639) );
  NOR2X1 U18449 ( .A(n44748), .B(n44546), .Y(n19640) );
  NOR2X1 U18452 ( .A(n44690), .B(n44555), .Y(n19645) );
  NOR2X1 U18456 ( .A(n44752), .B(n44546), .Y(n19646) );
  NOR2X1 U18459 ( .A(n44688), .B(n44555), .Y(n19651) );
  NOR2X1 U18463 ( .A(n44754), .B(n44546), .Y(n19652) );
  NOR2X1 U18466 ( .A(n44686), .B(n44555), .Y(n19657) );
  NOR2X1 U18470 ( .A(n44756), .B(n44546), .Y(n19658) );
  NOR2X1 U18473 ( .A(n44684), .B(n44555), .Y(n19663) );
  NOR2X1 U18477 ( .A(n44750), .B(n44546), .Y(n19664) );
  NOR2X1 U18480 ( .A(n44682), .B(n44555), .Y(n19669) );
  NAND2X1 U18482 ( .A(n520), .B(n44549), .Y(n19481) );
  NOR2X1 U18485 ( .A(n44746), .B(n44546), .Y(n19671) );
  NOR2X1 U18488 ( .A(n44680), .B(n44541), .Y(n19676) );
  NOR2X1 U18492 ( .A(n44708), .B(n44532), .Y(n19679) );
  NOR2X1 U18495 ( .A(n44642), .B(n44541), .Y(n19686) );
  NOR2X1 U18499 ( .A(n44706), .B(n44532), .Y(n19687) );
  NOR2X1 U18502 ( .A(n44648), .B(n44541), .Y(n19692) );
  NOR2X1 U18506 ( .A(n44714), .B(n44532), .Y(n19693) );
  NOR2X1 U18509 ( .A(n44650), .B(n44541), .Y(n19698) );
  NOR2X1 U18513 ( .A(n44716), .B(n44532), .Y(n19699) );
  NOR2X1 U18516 ( .A(n44672), .B(n44541), .Y(n19704) );
  NOR2X1 U18520 ( .A(n44738), .B(n44532), .Y(n19705) );
  NOR2X1 U18523 ( .A(n44664), .B(n44541), .Y(n19710) );
  NOR2X1 U18527 ( .A(n44730), .B(n44532), .Y(n19711) );
  NOR2X1 U18530 ( .A(n44674), .B(n44541), .Y(n19716) );
  NOR2X1 U18534 ( .A(n44740), .B(n44532), .Y(n19717) );
  NOR2X1 U18537 ( .A(n44676), .B(n44541), .Y(n19722) );
  NOR2X1 U18541 ( .A(n44742), .B(n44532), .Y(n19723) );
  NOR2X1 U18544 ( .A(n44656), .B(n44541), .Y(n19728) );
  NOR2X1 U18548 ( .A(n44722), .B(n44532), .Y(n19729) );
  NOR2X1 U18551 ( .A(n44658), .B(n44541), .Y(n19734) );
  NOR2X1 U18555 ( .A(n44724), .B(n44532), .Y(n19735) );
  NOR2X1 U18558 ( .A(n44662), .B(n44541), .Y(n19740) );
  NOR2X1 U18562 ( .A(n44728), .B(n44532), .Y(n19741) );
  NOR2X1 U18565 ( .A(n44654), .B(n44541), .Y(n19746) );
  NOR2X1 U18569 ( .A(n44720), .B(n44532), .Y(n19747) );
  NOR2X1 U18572 ( .A(n44652), .B(n44542), .Y(n19752) );
  NOR2X1 U18576 ( .A(n44718), .B(n44533), .Y(n19753) );
  NOR2X1 U18579 ( .A(n44666), .B(n44542), .Y(n19758) );
  NOR2X1 U18583 ( .A(n44732), .B(n44533), .Y(n19759) );
  NOR2X1 U18586 ( .A(n44678), .B(n44542), .Y(n19764) );
  NOR2X1 U18590 ( .A(n44744), .B(n44533), .Y(n19765) );
  NOR2X1 U18593 ( .A(n44660), .B(n44542), .Y(n19770) );
  NOR2X1 U18597 ( .A(n44726), .B(n44533), .Y(n19771) );
  NOR2X1 U18600 ( .A(n44644), .B(n44542), .Y(n19776) );
  NOR2X1 U18604 ( .A(n44710), .B(n44533), .Y(n19777) );
  NOR2X1 U18607 ( .A(n44646), .B(n44542), .Y(n19782) );
  NOR2X1 U18611 ( .A(n44712), .B(n44533), .Y(n19783) );
  NOR2X1 U18614 ( .A(n44670), .B(n44542), .Y(n19788) );
  NOR2X1 U18618 ( .A(n44736), .B(n44533), .Y(n19789) );
  NOR2X1 U18621 ( .A(n44668), .B(n44542), .Y(n19794) );
  NOR2X1 U18625 ( .A(n44734), .B(n44533), .Y(n19795) );
  NOR2X1 U18628 ( .A(n44694), .B(n44542), .Y(n19800) );
  NOR2X1 U18632 ( .A(n44758), .B(n44533), .Y(n19801) );
  NOR2X1 U18635 ( .A(n44698), .B(n44542), .Y(n19806) );
  NOR2X1 U18639 ( .A(n44762), .B(n44533), .Y(n19807) );
  NOR2X1 U18642 ( .A(n44700), .B(n44542), .Y(n19812) );
  NOR2X1 U18646 ( .A(n44764), .B(n44533), .Y(n19813) );
  NOR2X1 U18649 ( .A(n44704), .B(n44542), .Y(n19818) );
  NOR2X1 U18653 ( .A(n44768), .B(n44533), .Y(n19819) );
  NOR2X1 U18656 ( .A(n44702), .B(n44543), .Y(n19824) );
  NOR2X1 U18660 ( .A(n44766), .B(n44534), .Y(n19825) );
  NOR2X1 U18663 ( .A(n44696), .B(n44543), .Y(n19830) );
  NOR2X1 U18667 ( .A(n44760), .B(n44534), .Y(n19831) );
  NOR2X1 U18670 ( .A(n44692), .B(n44543), .Y(n19836) );
  NOR2X1 U18674 ( .A(n44748), .B(n44534), .Y(n19837) );
  NOR2X1 U18677 ( .A(n44690), .B(n44543), .Y(n19842) );
  NOR2X1 U18681 ( .A(n44752), .B(n44534), .Y(n19843) );
  NOR2X1 U18684 ( .A(n44688), .B(n44543), .Y(n19848) );
  NOR2X1 U18688 ( .A(n44754), .B(n44534), .Y(n19849) );
  NOR2X1 U18691 ( .A(n44686), .B(n44543), .Y(n19854) );
  NOR2X1 U18695 ( .A(n44756), .B(n44534), .Y(n19855) );
  NOR2X1 U18698 ( .A(n44684), .B(n44543), .Y(n19860) );
  NOR2X1 U18702 ( .A(n44750), .B(n44534), .Y(n19861) );
  NOR2X1 U18705 ( .A(n44682), .B(n44543), .Y(n19866) );
  NAND2X1 U18707 ( .A(n513), .B(n44537), .Y(n19678) );
  NOR2X1 U18710 ( .A(n44746), .B(n44534), .Y(n19868) );
  NOR2X1 U18713 ( .A(n44680), .B(n44529), .Y(n19873) );
  NOR2X1 U18717 ( .A(n44708), .B(n44520), .Y(n19876) );
  NOR2X1 U18720 ( .A(n44642), .B(n44529), .Y(n19883) );
  NOR2X1 U18724 ( .A(n44706), .B(n44520), .Y(n19884) );
  NOR2X1 U18727 ( .A(n44648), .B(n44529), .Y(n19889) );
  NOR2X1 U18731 ( .A(n44714), .B(n44520), .Y(n19890) );
  NOR2X1 U18734 ( .A(n44650), .B(n44529), .Y(n19895) );
  NOR2X1 U18738 ( .A(n44716), .B(n44520), .Y(n19896) );
  NOR2X1 U18741 ( .A(n44672), .B(n44529), .Y(n19901) );
  NOR2X1 U18745 ( .A(n44738), .B(n44520), .Y(n19902) );
  NOR2X1 U18748 ( .A(n44664), .B(n44529), .Y(n19907) );
  NOR2X1 U18752 ( .A(n44730), .B(n44520), .Y(n19908) );
  NOR2X1 U18755 ( .A(n44674), .B(n44529), .Y(n19913) );
  NOR2X1 U18759 ( .A(n44740), .B(n44520), .Y(n19914) );
  NOR2X1 U18762 ( .A(n44676), .B(n44529), .Y(n19919) );
  NOR2X1 U18766 ( .A(n44742), .B(n44520), .Y(n19920) );
  NOR2X1 U18769 ( .A(n44656), .B(n44529), .Y(n19925) );
  NOR2X1 U18773 ( .A(n44722), .B(n44520), .Y(n19926) );
  NOR2X1 U18776 ( .A(n44658), .B(n44529), .Y(n19931) );
  NOR2X1 U18780 ( .A(n44724), .B(n44520), .Y(n19932) );
  NOR2X1 U18783 ( .A(n44662), .B(n44529), .Y(n19937) );
  NOR2X1 U18787 ( .A(n44728), .B(n44520), .Y(n19938) );
  NOR2X1 U18790 ( .A(n44654), .B(n44529), .Y(n19943) );
  NOR2X1 U18794 ( .A(n44720), .B(n44520), .Y(n19944) );
  NOR2X1 U18797 ( .A(n44652), .B(n44530), .Y(n19949) );
  NOR2X1 U18801 ( .A(n44718), .B(n44521), .Y(n19950) );
  NOR2X1 U18804 ( .A(n44666), .B(n44530), .Y(n19955) );
  NOR2X1 U18808 ( .A(n44732), .B(n44521), .Y(n19956) );
  NOR2X1 U18811 ( .A(n44678), .B(n44530), .Y(n19961) );
  NOR2X1 U18815 ( .A(n44744), .B(n44521), .Y(n19962) );
  NOR2X1 U18818 ( .A(n44660), .B(n44530), .Y(n19967) );
  NOR2X1 U18822 ( .A(n44726), .B(n44521), .Y(n19968) );
  NOR2X1 U18825 ( .A(n44644), .B(n44530), .Y(n19973) );
  NOR2X1 U18829 ( .A(n44710), .B(n44521), .Y(n19974) );
  NOR2X1 U18832 ( .A(n44646), .B(n44530), .Y(n19979) );
  NOR2X1 U18836 ( .A(n44712), .B(n44521), .Y(n19980) );
  NOR2X1 U18839 ( .A(n44670), .B(n44530), .Y(n19985) );
  NOR2X1 U18843 ( .A(n44736), .B(n44521), .Y(n19986) );
  NOR2X1 U18846 ( .A(n44668), .B(n44530), .Y(n19991) );
  NOR2X1 U18850 ( .A(n44734), .B(n44521), .Y(n19992) );
  NOR2X1 U18853 ( .A(n44694), .B(n44530), .Y(n19997) );
  NOR2X1 U18857 ( .A(n44758), .B(n44521), .Y(n19998) );
  NOR2X1 U18860 ( .A(n44698), .B(n44530), .Y(n20003) );
  NOR2X1 U18864 ( .A(n44762), .B(n44521), .Y(n20004) );
  NOR2X1 U18867 ( .A(n44700), .B(n44530), .Y(n20009) );
  NOR2X1 U18871 ( .A(n44764), .B(n44521), .Y(n20010) );
  NOR2X1 U18874 ( .A(n44704), .B(n44530), .Y(n20015) );
  NOR2X1 U18878 ( .A(n44768), .B(n44521), .Y(n20016) );
  NOR2X1 U18881 ( .A(n44702), .B(n44531), .Y(n20021) );
  NOR2X1 U18885 ( .A(n44766), .B(n44522), .Y(n20022) );
  NOR2X1 U18888 ( .A(n44696), .B(n44531), .Y(n20027) );
  NOR2X1 U18892 ( .A(n44760), .B(n44522), .Y(n20028) );
  NOR2X1 U18895 ( .A(n44692), .B(n44531), .Y(n20033) );
  NOR2X1 U18899 ( .A(n44748), .B(n44522), .Y(n20034) );
  NOR2X1 U18902 ( .A(n44690), .B(n44531), .Y(n20039) );
  NOR2X1 U18906 ( .A(n44752), .B(n44522), .Y(n20040) );
  NOR2X1 U18909 ( .A(n44688), .B(n44531), .Y(n20045) );
  NOR2X1 U18913 ( .A(n44754), .B(n44522), .Y(n20046) );
  NOR2X1 U18916 ( .A(n44686), .B(n44531), .Y(n20051) );
  NOR2X1 U18920 ( .A(n44756), .B(n44522), .Y(n20052) );
  NOR2X1 U18923 ( .A(n44684), .B(n44531), .Y(n20057) );
  NOR2X1 U18927 ( .A(n44750), .B(n44522), .Y(n20058) );
  NOR2X1 U18930 ( .A(n44682), .B(n44531), .Y(n20063) );
  NAND2X1 U18932 ( .A(n495), .B(n44525), .Y(n19875) );
  NOR2X1 U18935 ( .A(n44746), .B(n44522), .Y(n20064) );
  NOR2X1 U18938 ( .A(n44680), .B(n44517), .Y(n20069) );
  NOR2X1 U18942 ( .A(n44708), .B(n44508), .Y(n20072) );
  NOR2X1 U18945 ( .A(n44642), .B(n44517), .Y(n20079) );
  NOR2X1 U18949 ( .A(n44706), .B(n44508), .Y(n20080) );
  NOR2X1 U18952 ( .A(n44648), .B(n44517), .Y(n20085) );
  NOR2X1 U18956 ( .A(n44714), .B(n44508), .Y(n20086) );
  NOR2X1 U18959 ( .A(n44650), .B(n44517), .Y(n20091) );
  NOR2X1 U18963 ( .A(n44716), .B(n44508), .Y(n20092) );
  NOR2X1 U18966 ( .A(n44672), .B(n44517), .Y(n20097) );
  NOR2X1 U18970 ( .A(n44738), .B(n44508), .Y(n20098) );
  NOR2X1 U18973 ( .A(n44664), .B(n44517), .Y(n20103) );
  NOR2X1 U18977 ( .A(n44730), .B(n44508), .Y(n20104) );
  NOR2X1 U18980 ( .A(n44674), .B(n44517), .Y(n20109) );
  NOR2X1 U18984 ( .A(n44740), .B(n44508), .Y(n20110) );
  NOR2X1 U18987 ( .A(n44676), .B(n44517), .Y(n20115) );
  NOR2X1 U18991 ( .A(n44742), .B(n44508), .Y(n20116) );
  NOR2X1 U18994 ( .A(n44656), .B(n44517), .Y(n20121) );
  NOR2X1 U18998 ( .A(n44722), .B(n44508), .Y(n20122) );
  NOR2X1 U19001 ( .A(n44658), .B(n44517), .Y(n20127) );
  NOR2X1 U19005 ( .A(n44724), .B(n44508), .Y(n20128) );
  NOR2X1 U19008 ( .A(n44662), .B(n44517), .Y(n20133) );
  NOR2X1 U19012 ( .A(n44728), .B(n44508), .Y(n20134) );
  NOR2X1 U19015 ( .A(n44654), .B(n44517), .Y(n20139) );
  NOR2X1 U19019 ( .A(n44720), .B(n44508), .Y(n20140) );
  NOR2X1 U19022 ( .A(n44652), .B(n44518), .Y(n20145) );
  NOR2X1 U19026 ( .A(n44718), .B(n44509), .Y(n20146) );
  NOR2X1 U19029 ( .A(n44666), .B(n44518), .Y(n20151) );
  NOR2X1 U19033 ( .A(n44732), .B(n44509), .Y(n20152) );
  NOR2X1 U19036 ( .A(n44678), .B(n44518), .Y(n20157) );
  NOR2X1 U19040 ( .A(n44744), .B(n44509), .Y(n20158) );
  NOR2X1 U19043 ( .A(n44660), .B(n44518), .Y(n20163) );
  NOR2X1 U19047 ( .A(n44726), .B(n44509), .Y(n20164) );
  NOR2X1 U19050 ( .A(n44644), .B(n44518), .Y(n20169) );
  NOR2X1 U19054 ( .A(n44710), .B(n44509), .Y(n20170) );
  NOR2X1 U19057 ( .A(n44646), .B(n44518), .Y(n20175) );
  NOR2X1 U19061 ( .A(n44712), .B(n44509), .Y(n20176) );
  NOR2X1 U19064 ( .A(n44670), .B(n44518), .Y(n20181) );
  NOR2X1 U19068 ( .A(n44736), .B(n44509), .Y(n20182) );
  NOR2X1 U19071 ( .A(n44668), .B(n44518), .Y(n20187) );
  NOR2X1 U19075 ( .A(n44734), .B(n44509), .Y(n20188) );
  NOR2X1 U19078 ( .A(n44694), .B(n44518), .Y(n20193) );
  NOR2X1 U19082 ( .A(n44758), .B(n44509), .Y(n20194) );
  NOR2X1 U19085 ( .A(n44698), .B(n44518), .Y(n20199) );
  NOR2X1 U19089 ( .A(n44762), .B(n44509), .Y(n20200) );
  NOR2X1 U19092 ( .A(n44700), .B(n44518), .Y(n20205) );
  NOR2X1 U19096 ( .A(n44764), .B(n44509), .Y(n20206) );
  NOR2X1 U19099 ( .A(n44704), .B(n44518), .Y(n20211) );
  NOR2X1 U19103 ( .A(n44768), .B(n44509), .Y(n20212) );
  NOR2X1 U19106 ( .A(n44702), .B(n44519), .Y(n20217) );
  NOR2X1 U19110 ( .A(n44766), .B(n44510), .Y(n20218) );
  NOR2X1 U19113 ( .A(n44696), .B(n44519), .Y(n20223) );
  NOR2X1 U19117 ( .A(n44760), .B(n44510), .Y(n20224) );
  NOR2X1 U19120 ( .A(n44692), .B(n44519), .Y(n20229) );
  NOR2X1 U19124 ( .A(n44748), .B(n44510), .Y(n20230) );
  NOR2X1 U19127 ( .A(n44690), .B(n44519), .Y(n20235) );
  NOR2X1 U19131 ( .A(n44752), .B(n44510), .Y(n20236) );
  NOR2X1 U19134 ( .A(n44688), .B(n44519), .Y(n20241) );
  NOR2X1 U19138 ( .A(n44754), .B(n44510), .Y(n20242) );
  NOR2X1 U19141 ( .A(n44686), .B(n44519), .Y(n20247) );
  NOR2X1 U19145 ( .A(n44756), .B(n44510), .Y(n20248) );
  NOR2X1 U19148 ( .A(n44684), .B(n44519), .Y(n20253) );
  NOR2X1 U19152 ( .A(n44750), .B(n44510), .Y(n20254) );
  NOR2X1 U19155 ( .A(n44682), .B(n44519), .Y(n20259) );
  NAND2X1 U19157 ( .A(n503), .B(n44513), .Y(n20071) );
  NOR2X1 U19160 ( .A(n44746), .B(n44510), .Y(n20260) );
  NOR2X1 U19163 ( .A(n44680), .B(n44505), .Y(n20265) );
  NOR2X1 U19167 ( .A(n44708), .B(n44496), .Y(n20268) );
  NOR2X1 U19170 ( .A(n44642), .B(n44505), .Y(n20275) );
  NOR2X1 U19174 ( .A(n44706), .B(n44496), .Y(n20276) );
  NOR2X1 U19177 ( .A(n44648), .B(n44505), .Y(n20281) );
  NOR2X1 U19181 ( .A(n44714), .B(n44496), .Y(n20282) );
  NOR2X1 U19184 ( .A(n44650), .B(n44505), .Y(n20287) );
  NOR2X1 U19188 ( .A(n44716), .B(n44496), .Y(n20288) );
  NOR2X1 U19191 ( .A(n44672), .B(n44505), .Y(n20293) );
  NOR2X1 U19195 ( .A(n44738), .B(n44496), .Y(n20294) );
  NOR2X1 U19198 ( .A(n44664), .B(n44505), .Y(n20299) );
  NOR2X1 U19202 ( .A(n44730), .B(n44496), .Y(n20300) );
  NOR2X1 U19205 ( .A(n44674), .B(n44505), .Y(n20305) );
  NOR2X1 U19209 ( .A(n44740), .B(n44496), .Y(n20306) );
  NOR2X1 U19212 ( .A(n44676), .B(n44505), .Y(n20311) );
  NOR2X1 U19216 ( .A(n44742), .B(n44496), .Y(n20312) );
  NOR2X1 U19219 ( .A(n44656), .B(n44505), .Y(n20317) );
  NOR2X1 U19223 ( .A(n44722), .B(n44496), .Y(n20318) );
  NOR2X1 U19226 ( .A(n44658), .B(n44505), .Y(n20323) );
  NOR2X1 U19230 ( .A(n44724), .B(n44496), .Y(n20324) );
  NOR2X1 U19233 ( .A(n44662), .B(n44505), .Y(n20329) );
  NOR2X1 U19237 ( .A(n44728), .B(n44496), .Y(n20330) );
  NOR2X1 U19240 ( .A(n44654), .B(n44505), .Y(n20335) );
  NOR2X1 U19244 ( .A(n44720), .B(n44496), .Y(n20336) );
  NOR2X1 U19247 ( .A(n44652), .B(n44506), .Y(n20341) );
  NOR2X1 U19251 ( .A(n44718), .B(n44497), .Y(n20342) );
  NOR2X1 U19254 ( .A(n44666), .B(n44506), .Y(n20347) );
  NOR2X1 U19258 ( .A(n44732), .B(n44497), .Y(n20348) );
  NOR2X1 U19261 ( .A(n44678), .B(n44506), .Y(n20353) );
  NOR2X1 U19265 ( .A(n44744), .B(n44497), .Y(n20354) );
  NOR2X1 U19268 ( .A(n44660), .B(n44506), .Y(n20359) );
  NOR2X1 U19272 ( .A(n44726), .B(n44497), .Y(n20360) );
  NOR2X1 U19275 ( .A(n44644), .B(n44506), .Y(n20365) );
  NOR2X1 U19279 ( .A(n44710), .B(n44497), .Y(n20366) );
  NOR2X1 U19282 ( .A(n44646), .B(n44506), .Y(n20371) );
  NOR2X1 U19286 ( .A(n44712), .B(n44497), .Y(n20372) );
  NOR2X1 U19289 ( .A(n44670), .B(n44506), .Y(n20377) );
  NOR2X1 U19293 ( .A(n44736), .B(n44497), .Y(n20378) );
  NOR2X1 U19296 ( .A(n44668), .B(n44506), .Y(n20383) );
  NOR2X1 U19300 ( .A(n44734), .B(n44497), .Y(n20384) );
  NOR2X1 U19303 ( .A(n44694), .B(n44506), .Y(n20389) );
  NOR2X1 U19307 ( .A(n44758), .B(n44497), .Y(n20390) );
  NOR2X1 U19310 ( .A(n44698), .B(n44506), .Y(n20395) );
  NOR2X1 U19314 ( .A(n44762), .B(n44497), .Y(n20396) );
  NOR2X1 U19317 ( .A(n44700), .B(n44506), .Y(n20401) );
  NOR2X1 U19321 ( .A(n44764), .B(n44497), .Y(n20402) );
  NOR2X1 U19324 ( .A(n44704), .B(n44506), .Y(n20407) );
  NOR2X1 U19328 ( .A(n44768), .B(n44497), .Y(n20408) );
  NOR2X1 U19331 ( .A(n44702), .B(n44507), .Y(n20413) );
  NOR2X1 U19335 ( .A(n44766), .B(n44498), .Y(n20414) );
  NOR2X1 U19338 ( .A(n44696), .B(n44507), .Y(n20419) );
  NOR2X1 U19342 ( .A(n44760), .B(n44498), .Y(n20420) );
  NOR2X1 U19345 ( .A(n44692), .B(n44507), .Y(n20425) );
  NOR2X1 U19349 ( .A(n44748), .B(n44498), .Y(n20426) );
  NOR2X1 U19352 ( .A(n44690), .B(n44507), .Y(n20431) );
  NOR2X1 U19356 ( .A(n44752), .B(n44498), .Y(n20432) );
  NOR2X1 U19359 ( .A(n44688), .B(n44507), .Y(n20437) );
  NOR2X1 U19363 ( .A(n44754), .B(n44498), .Y(n20438) );
  NOR2X1 U19366 ( .A(n44686), .B(n44507), .Y(n20443) );
  NOR2X1 U19370 ( .A(n44756), .B(n44498), .Y(n20444) );
  NOR2X1 U19373 ( .A(n44684), .B(n44507), .Y(n20449) );
  NOR2X1 U19377 ( .A(n44750), .B(n44498), .Y(n20450) );
  NOR2X1 U19380 ( .A(n44682), .B(n44507), .Y(n20455) );
  NAND2X1 U19382 ( .A(n497), .B(n44501), .Y(n20267) );
  NOR2X1 U19385 ( .A(n44746), .B(n44498), .Y(n20456) );
  NOR2X1 U19388 ( .A(n44680), .B(n44493), .Y(n20461) );
  NOR2X1 U19392 ( .A(n44708), .B(n44490), .Y(n20464) );
  NOR2X1 U19395 ( .A(n44642), .B(n44493), .Y(n20471) );
  NOR2X1 U19399 ( .A(n44706), .B(n44490), .Y(n20472) );
  NOR2X1 U19402 ( .A(n44648), .B(n44493), .Y(n20477) );
  NOR2X1 U19406 ( .A(n44714), .B(n44490), .Y(n20478) );
  NOR2X1 U19409 ( .A(n44650), .B(n44493), .Y(n20483) );
  NOR2X1 U19413 ( .A(n44716), .B(n44490), .Y(n20484) );
  NOR2X1 U19416 ( .A(n44672), .B(n44493), .Y(n20489) );
  NOR2X1 U19420 ( .A(n44738), .B(n44490), .Y(n20490) );
  NOR2X1 U19423 ( .A(n44664), .B(n44493), .Y(n20495) );
  NOR2X1 U19427 ( .A(n44730), .B(n44490), .Y(n20496) );
  NOR2X1 U19430 ( .A(n44674), .B(n44493), .Y(n20501) );
  NOR2X1 U19434 ( .A(n44740), .B(n44490), .Y(n20502) );
  NOR2X1 U19437 ( .A(n44676), .B(n44493), .Y(n20507) );
  NOR2X1 U19441 ( .A(n44742), .B(n44490), .Y(n20508) );
  NOR2X1 U19444 ( .A(n44656), .B(n44493), .Y(n20513) );
  NOR2X1 U19448 ( .A(n44722), .B(n44490), .Y(n20514) );
  NOR2X1 U19451 ( .A(n44658), .B(n44493), .Y(n20519) );
  NOR2X1 U19455 ( .A(n44724), .B(n44490), .Y(n20520) );
  NOR2X1 U19458 ( .A(n44662), .B(n44493), .Y(n20525) );
  NOR2X1 U19462 ( .A(n44728), .B(n44490), .Y(n20526) );
  NOR2X1 U19465 ( .A(n44654), .B(n44493), .Y(n20531) );
  NOR2X1 U19469 ( .A(n44720), .B(n44490), .Y(n20532) );
  NOR2X1 U19472 ( .A(n44652), .B(n44494), .Y(n20537) );
  NOR2X1 U19476 ( .A(n44718), .B(n44491), .Y(n20538) );
  NOR2X1 U19479 ( .A(n44666), .B(n44494), .Y(n20543) );
  NOR2X1 U19483 ( .A(n44732), .B(n44491), .Y(n20544) );
  NOR2X1 U19486 ( .A(n44678), .B(n44494), .Y(n20549) );
  NOR2X1 U19490 ( .A(n44744), .B(n44491), .Y(n20550) );
  NOR2X1 U19493 ( .A(n44660), .B(n44494), .Y(n20555) );
  NOR2X1 U19497 ( .A(n44726), .B(n44491), .Y(n20556) );
  NOR2X1 U19500 ( .A(n44644), .B(n44494), .Y(n20561) );
  NOR2X1 U19504 ( .A(n44710), .B(n44491), .Y(n20562) );
  NOR2X1 U19507 ( .A(n44646), .B(n44494), .Y(n20567) );
  NOR2X1 U19511 ( .A(n44712), .B(n44491), .Y(n20568) );
  NOR2X1 U19514 ( .A(n44670), .B(n44494), .Y(n20573) );
  NOR2X1 U19518 ( .A(n44736), .B(n44491), .Y(n20574) );
  NOR2X1 U19521 ( .A(n44668), .B(n44494), .Y(n20579) );
  NOR2X1 U19525 ( .A(n44734), .B(n44491), .Y(n20580) );
  NOR2X1 U19528 ( .A(n44694), .B(n44494), .Y(n20585) );
  NOR2X1 U19532 ( .A(n44758), .B(n44491), .Y(n20586) );
  NOR2X1 U19535 ( .A(n44698), .B(n44494), .Y(n20591) );
  NOR2X1 U19539 ( .A(n44762), .B(n44491), .Y(n20592) );
  NOR2X1 U19542 ( .A(n44700), .B(n44494), .Y(n20597) );
  NOR2X1 U19546 ( .A(n44764), .B(n44491), .Y(n20598) );
  NOR2X1 U19549 ( .A(n44704), .B(n44494), .Y(n20603) );
  NOR2X1 U19553 ( .A(n44768), .B(n44491), .Y(n20604) );
  NOR2X1 U19556 ( .A(n44702), .B(n44495), .Y(n20609) );
  NOR2X1 U19560 ( .A(n44766), .B(n44492), .Y(n20610) );
  NOR2X1 U19563 ( .A(n44696), .B(n44495), .Y(n20615) );
  NOR2X1 U19567 ( .A(n44760), .B(n44492), .Y(n20616) );
  NOR2X1 U19570 ( .A(n44692), .B(n44495), .Y(n20621) );
  NOR2X1 U19574 ( .A(n44748), .B(n44492), .Y(n20622) );
  NOR2X1 U19577 ( .A(n44690), .B(n44495), .Y(n20627) );
  NOR2X1 U19581 ( .A(n44752), .B(n44492), .Y(n20628) );
  NOR2X1 U19584 ( .A(n44688), .B(n44495), .Y(n20633) );
  NOR2X1 U19588 ( .A(n44754), .B(n44492), .Y(n20634) );
  NOR2X1 U19591 ( .A(n44686), .B(n44495), .Y(n20639) );
  NOR2X1 U19595 ( .A(n44756), .B(n44492), .Y(n20640) );
  NOR2X1 U19598 ( .A(n44684), .B(n44495), .Y(n20645) );
  NOR2X1 U19602 ( .A(n44750), .B(n44492), .Y(n20646) );
  NOR2X1 U19605 ( .A(n44682), .B(n44495), .Y(n20651) );
  NOR2X1 U19610 ( .A(n44746), .B(n44492), .Y(n20652) );
  NOR2X1 U19613 ( .A(n44680), .B(n44487), .Y(n20657) );
  NOR2X1 U19617 ( .A(n44708), .B(n44478), .Y(n20660) );
  NOR2X1 U19620 ( .A(n44642), .B(n44487), .Y(n20667) );
  NOR2X1 U19624 ( .A(n44706), .B(n44478), .Y(n20668) );
  NOR2X1 U19627 ( .A(n44648), .B(n44487), .Y(n20673) );
  NOR2X1 U19631 ( .A(n44714), .B(n44478), .Y(n20674) );
  NOR2X1 U19634 ( .A(n44650), .B(n44487), .Y(n20679) );
  NOR2X1 U19638 ( .A(n44716), .B(n44478), .Y(n20680) );
  NOR2X1 U19641 ( .A(n44672), .B(n44487), .Y(n20685) );
  NOR2X1 U19645 ( .A(n44738), .B(n44478), .Y(n20686) );
  NOR2X1 U19648 ( .A(n44664), .B(n44487), .Y(n20691) );
  NOR2X1 U19652 ( .A(n44730), .B(n44478), .Y(n20692) );
  NOR2X1 U19655 ( .A(n44674), .B(n44487), .Y(n20697) );
  NOR2X1 U19659 ( .A(n44740), .B(n44478), .Y(n20698) );
  NOR2X1 U19662 ( .A(n44676), .B(n44487), .Y(n20703) );
  NOR2X1 U19666 ( .A(n44742), .B(n44478), .Y(n20704) );
  NOR2X1 U19669 ( .A(n44656), .B(n44487), .Y(n20709) );
  NOR2X1 U19673 ( .A(n44722), .B(n44478), .Y(n20710) );
  NOR2X1 U19676 ( .A(n44658), .B(n44487), .Y(n20715) );
  NOR2X1 U19680 ( .A(n44724), .B(n44478), .Y(n20716) );
  NOR2X1 U19683 ( .A(n44662), .B(n44487), .Y(n20721) );
  NOR2X1 U19687 ( .A(n44728), .B(n44478), .Y(n20722) );
  NOR2X1 U19690 ( .A(n44654), .B(n44487), .Y(n20727) );
  NOR2X1 U19694 ( .A(n44720), .B(n44478), .Y(n20728) );
  NOR2X1 U19697 ( .A(n44652), .B(n44488), .Y(n20733) );
  NOR2X1 U19701 ( .A(n44718), .B(n44479), .Y(n20734) );
  NOR2X1 U19704 ( .A(n44666), .B(n44488), .Y(n20739) );
  NOR2X1 U19708 ( .A(n44732), .B(n44479), .Y(n20740) );
  NOR2X1 U19711 ( .A(n44678), .B(n44488), .Y(n20745) );
  NOR2X1 U19715 ( .A(n44744), .B(n44479), .Y(n20746) );
  NOR2X1 U19718 ( .A(n44660), .B(n44488), .Y(n20751) );
  NOR2X1 U19722 ( .A(n44726), .B(n44479), .Y(n20752) );
  NOR2X1 U19725 ( .A(n44644), .B(n44488), .Y(n20757) );
  NOR2X1 U19729 ( .A(n44710), .B(n44479), .Y(n20758) );
  NOR2X1 U19732 ( .A(n44646), .B(n44488), .Y(n20763) );
  NOR2X1 U19736 ( .A(n44712), .B(n44479), .Y(n20764) );
  NOR2X1 U19739 ( .A(n44670), .B(n44488), .Y(n20769) );
  NOR2X1 U19743 ( .A(n44736), .B(n44479), .Y(n20770) );
  NOR2X1 U19746 ( .A(n44668), .B(n44488), .Y(n20775) );
  NOR2X1 U19750 ( .A(n44734), .B(n44479), .Y(n20776) );
  NOR2X1 U19753 ( .A(n44694), .B(n44488), .Y(n20781) );
  NOR2X1 U19757 ( .A(n44758), .B(n44479), .Y(n20782) );
  NOR2X1 U19760 ( .A(n44698), .B(n44488), .Y(n20787) );
  NOR2X1 U19764 ( .A(n44762), .B(n44479), .Y(n20788) );
  NOR2X1 U19767 ( .A(n44700), .B(n44488), .Y(n20793) );
  NOR2X1 U19771 ( .A(n44764), .B(n44479), .Y(n20794) );
  NOR2X1 U19774 ( .A(n44704), .B(n44488), .Y(n20799) );
  NOR2X1 U19778 ( .A(n44768), .B(n44479), .Y(n20800) );
  NOR2X1 U19781 ( .A(n44702), .B(n44489), .Y(n20805) );
  NOR2X1 U19785 ( .A(n44766), .B(n44480), .Y(n20806) );
  NOR2X1 U19788 ( .A(n44696), .B(n44489), .Y(n20811) );
  NOR2X1 U19792 ( .A(n44760), .B(n44480), .Y(n20812) );
  NOR2X1 U19795 ( .A(n44692), .B(n44489), .Y(n20817) );
  NOR2X1 U19799 ( .A(n44748), .B(n44480), .Y(n20818) );
  NOR2X1 U19802 ( .A(n44690), .B(n44489), .Y(n20823) );
  NOR2X1 U19806 ( .A(n44752), .B(n44480), .Y(n20824) );
  NOR2X1 U19809 ( .A(n44688), .B(n44489), .Y(n20829) );
  NOR2X1 U19813 ( .A(n44754), .B(n44480), .Y(n20830) );
  NOR2X1 U19816 ( .A(n44686), .B(n44489), .Y(n20835) );
  NOR2X1 U19820 ( .A(n44756), .B(n44480), .Y(n20836) );
  NOR2X1 U19823 ( .A(n44684), .B(n44489), .Y(n20841) );
  NOR2X1 U19827 ( .A(n44750), .B(n44480), .Y(n20842) );
  NOR2X1 U19830 ( .A(n44682), .B(n44489), .Y(n20847) );
  NAND2X1 U19832 ( .A(n493), .B(n44483), .Y(n20659) );
  NOR2X1 U19835 ( .A(n44746), .B(n44480), .Y(n20848) );
  NOR2X1 U19838 ( .A(n44680), .B(n44475), .Y(n20853) );
  NOR2X1 U19842 ( .A(n44708), .B(n44466), .Y(n20856) );
  NOR2X1 U19845 ( .A(n44642), .B(n44475), .Y(n20863) );
  NOR2X1 U19849 ( .A(n44706), .B(n44466), .Y(n20864) );
  NOR2X1 U19852 ( .A(n44648), .B(n44475), .Y(n20869) );
  NOR2X1 U19856 ( .A(n44714), .B(n44466), .Y(n20870) );
  NOR2X1 U19859 ( .A(n44650), .B(n44475), .Y(n20875) );
  NOR2X1 U19863 ( .A(n44716), .B(n44466), .Y(n20876) );
  NOR2X1 U19866 ( .A(n44672), .B(n44475), .Y(n20881) );
  NOR2X1 U19870 ( .A(n44738), .B(n44466), .Y(n20882) );
  NOR2X1 U19873 ( .A(n44664), .B(n44475), .Y(n20887) );
  NOR2X1 U19877 ( .A(n44730), .B(n44466), .Y(n20888) );
  NOR2X1 U19880 ( .A(n44674), .B(n44475), .Y(n20893) );
  NOR2X1 U19884 ( .A(n44740), .B(n44466), .Y(n20894) );
  NOR2X1 U19887 ( .A(n44676), .B(n44475), .Y(n20899) );
  NOR2X1 U19891 ( .A(n44742), .B(n44466), .Y(n20900) );
  NOR2X1 U19894 ( .A(n44656), .B(n44475), .Y(n20905) );
  NOR2X1 U19898 ( .A(n44722), .B(n44466), .Y(n20906) );
  NOR2X1 U19901 ( .A(n44658), .B(n44475), .Y(n20911) );
  NOR2X1 U19905 ( .A(n44724), .B(n44466), .Y(n20912) );
  NOR2X1 U19908 ( .A(n44662), .B(n44475), .Y(n20917) );
  NOR2X1 U19912 ( .A(n44728), .B(n44466), .Y(n20918) );
  NOR2X1 U19915 ( .A(n44654), .B(n44475), .Y(n20923) );
  NOR2X1 U19919 ( .A(n44720), .B(n44466), .Y(n20924) );
  NOR2X1 U19922 ( .A(n44652), .B(n44476), .Y(n20929) );
  NOR2X1 U19926 ( .A(n44718), .B(n44467), .Y(n20930) );
  NOR2X1 U19929 ( .A(n44666), .B(n44476), .Y(n20935) );
  NOR2X1 U19933 ( .A(n44732), .B(n44467), .Y(n20936) );
  NOR2X1 U19936 ( .A(n44678), .B(n44476), .Y(n20941) );
  NOR2X1 U19940 ( .A(n44744), .B(n44467), .Y(n20942) );
  NOR2X1 U19943 ( .A(n44660), .B(n44476), .Y(n20947) );
  NOR2X1 U19947 ( .A(n44726), .B(n44467), .Y(n20948) );
  NOR2X1 U19950 ( .A(n44644), .B(n44476), .Y(n20953) );
  NOR2X1 U19954 ( .A(n44710), .B(n44467), .Y(n20954) );
  NOR2X1 U19957 ( .A(n44646), .B(n44476), .Y(n20959) );
  NOR2X1 U19961 ( .A(n44712), .B(n44467), .Y(n20960) );
  NOR2X1 U19964 ( .A(n44670), .B(n44476), .Y(n20965) );
  NOR2X1 U19968 ( .A(n44736), .B(n44467), .Y(n20966) );
  NOR2X1 U19971 ( .A(n44668), .B(n44476), .Y(n20971) );
  NOR2X1 U19975 ( .A(n44734), .B(n44467), .Y(n20972) );
  NOR2X1 U19978 ( .A(n44694), .B(n44476), .Y(n20977) );
  NOR2X1 U19982 ( .A(n44758), .B(n44467), .Y(n20978) );
  NOR2X1 U19985 ( .A(n44698), .B(n44476), .Y(n20983) );
  NOR2X1 U19989 ( .A(n44762), .B(n44467), .Y(n20984) );
  NOR2X1 U19992 ( .A(n44700), .B(n44476), .Y(n20989) );
  NOR2X1 U19996 ( .A(n44764), .B(n44467), .Y(n20990) );
  NOR2X1 U19999 ( .A(n44704), .B(n44476), .Y(n20995) );
  NOR2X1 U20003 ( .A(n44768), .B(n44467), .Y(n20996) );
  NOR2X1 U20006 ( .A(n44702), .B(n44477), .Y(n21001) );
  NOR2X1 U20010 ( .A(n44766), .B(n44468), .Y(n21002) );
  NOR2X1 U20013 ( .A(n44696), .B(n44477), .Y(n21007) );
  NOR2X1 U20017 ( .A(n44760), .B(n44468), .Y(n21008) );
  NOR2X1 U20020 ( .A(n44692), .B(n44477), .Y(n21013) );
  NOR2X1 U20024 ( .A(n44748), .B(n44468), .Y(n21014) );
  NOR2X1 U20027 ( .A(n44690), .B(n44477), .Y(n21019) );
  NOR2X1 U20031 ( .A(n44752), .B(n44468), .Y(n21020) );
  NOR2X1 U20034 ( .A(n44688), .B(n44477), .Y(n21025) );
  NOR2X1 U20038 ( .A(n44754), .B(n44468), .Y(n21026) );
  NOR2X1 U20041 ( .A(n44686), .B(n44477), .Y(n21031) );
  NOR2X1 U20045 ( .A(n44756), .B(n44468), .Y(n21032) );
  NOR2X1 U20048 ( .A(n44684), .B(n44477), .Y(n21037) );
  NOR2X1 U20052 ( .A(n44750), .B(n44468), .Y(n21038) );
  NOR2X1 U20055 ( .A(n44682), .B(n44477), .Y(n21043) );
  NOR2X1 U20060 ( .A(n44746), .B(n44468), .Y(n21044) );
  NOR2X1 U20063 ( .A(n44680), .B(n44463), .Y(n21049) );
  NOR2X1 U20067 ( .A(n44708), .B(n44454), .Y(n21052) );
  NOR2X1 U20070 ( .A(n44642), .B(n44463), .Y(n21059) );
  NOR2X1 U20074 ( .A(n44706), .B(n44454), .Y(n21060) );
  NOR2X1 U20077 ( .A(n44648), .B(n44463), .Y(n21065) );
  NOR2X1 U20081 ( .A(n44714), .B(n44454), .Y(n21066) );
  NOR2X1 U20084 ( .A(n44650), .B(n44463), .Y(n21071) );
  NOR2X1 U20088 ( .A(n44716), .B(n44454), .Y(n21072) );
  NOR2X1 U20091 ( .A(n44672), .B(n44463), .Y(n21077) );
  NOR2X1 U20095 ( .A(n44738), .B(n44454), .Y(n21078) );
  NOR2X1 U20098 ( .A(n44664), .B(n44463), .Y(n21083) );
  NOR2X1 U20102 ( .A(n44730), .B(n44454), .Y(n21084) );
  NOR2X1 U20105 ( .A(n44674), .B(n44463), .Y(n21089) );
  NOR2X1 U20109 ( .A(n44740), .B(n44454), .Y(n21090) );
  NOR2X1 U20112 ( .A(n44676), .B(n44463), .Y(n21095) );
  NOR2X1 U20116 ( .A(n44742), .B(n44454), .Y(n21096) );
  NOR2X1 U20119 ( .A(n44656), .B(n44463), .Y(n21101) );
  NOR2X1 U20123 ( .A(n44722), .B(n44454), .Y(n21102) );
  NOR2X1 U20126 ( .A(n44658), .B(n44463), .Y(n21107) );
  NOR2X1 U20130 ( .A(n44724), .B(n44454), .Y(n21108) );
  NOR2X1 U20133 ( .A(n44662), .B(n44463), .Y(n21113) );
  NOR2X1 U20137 ( .A(n44728), .B(n44454), .Y(n21114) );
  NOR2X1 U20140 ( .A(n44654), .B(n44463), .Y(n21119) );
  NOR2X1 U20144 ( .A(n44720), .B(n44454), .Y(n21120) );
  NOR2X1 U20147 ( .A(n44652), .B(n44464), .Y(n21125) );
  NOR2X1 U20151 ( .A(n44718), .B(n44455), .Y(n21126) );
  NOR2X1 U20154 ( .A(n44666), .B(n44464), .Y(n21131) );
  NOR2X1 U20158 ( .A(n44732), .B(n44455), .Y(n21132) );
  NOR2X1 U20161 ( .A(n44678), .B(n44464), .Y(n21137) );
  NOR2X1 U20165 ( .A(n44744), .B(n44455), .Y(n21138) );
  NOR2X1 U20168 ( .A(n44660), .B(n44464), .Y(n21143) );
  NOR2X1 U20172 ( .A(n44726), .B(n44455), .Y(n21144) );
  NOR2X1 U20175 ( .A(n44644), .B(n44464), .Y(n21149) );
  NOR2X1 U20179 ( .A(n44710), .B(n44455), .Y(n21150) );
  NOR2X1 U20182 ( .A(n44646), .B(n44464), .Y(n21155) );
  NOR2X1 U20186 ( .A(n44712), .B(n44455), .Y(n21156) );
  NOR2X1 U20189 ( .A(n44670), .B(n44464), .Y(n21161) );
  NOR2X1 U20193 ( .A(n44736), .B(n44455), .Y(n21162) );
  NOR2X1 U20196 ( .A(n44668), .B(n44464), .Y(n21167) );
  NOR2X1 U20200 ( .A(n44734), .B(n44455), .Y(n21168) );
  NOR2X1 U20203 ( .A(n44694), .B(n44464), .Y(n21173) );
  NOR2X1 U20207 ( .A(n44758), .B(n44455), .Y(n21174) );
  NOR2X1 U20210 ( .A(n44698), .B(n44464), .Y(n21179) );
  NOR2X1 U20214 ( .A(n44762), .B(n44455), .Y(n21180) );
  NOR2X1 U20217 ( .A(n44700), .B(n44464), .Y(n21185) );
  NOR2X1 U20221 ( .A(n44764), .B(n44455), .Y(n21186) );
  NOR2X1 U20224 ( .A(n44704), .B(n44464), .Y(n21191) );
  NOR2X1 U20228 ( .A(n44768), .B(n44455), .Y(n21192) );
  NOR2X1 U20231 ( .A(n44702), .B(n44465), .Y(n21197) );
  NOR2X1 U20235 ( .A(n44766), .B(n44456), .Y(n21198) );
  NOR2X1 U20238 ( .A(n44696), .B(n44465), .Y(n21203) );
  NOR2X1 U20242 ( .A(n44760), .B(n44456), .Y(n21204) );
  NOR2X1 U20245 ( .A(n44692), .B(n44465), .Y(n21209) );
  NOR2X1 U20249 ( .A(n44748), .B(n44456), .Y(n21210) );
  NOR2X1 U20252 ( .A(n44690), .B(n44465), .Y(n21215) );
  NOR2X1 U20256 ( .A(n44752), .B(n44456), .Y(n21216) );
  NOR2X1 U20259 ( .A(n44688), .B(n44465), .Y(n21221) );
  NOR2X1 U20263 ( .A(n44754), .B(n44456), .Y(n21222) );
  NOR2X1 U20266 ( .A(n44686), .B(n44465), .Y(n21227) );
  NOR2X1 U20270 ( .A(n44756), .B(n44456), .Y(n21228) );
  NOR2X1 U20273 ( .A(n44684), .B(n44465), .Y(n21233) );
  NOR2X1 U20277 ( .A(n44750), .B(n44456), .Y(n21234) );
  NOR2X1 U20280 ( .A(n44682), .B(n44465), .Y(n21239) );
  NAND2X1 U20282 ( .A(n492), .B(n44459), .Y(n21051) );
  NOR2X1 U20285 ( .A(n44746), .B(n44456), .Y(n21241) );
  NOR2X1 U20288 ( .A(n44680), .B(n44451), .Y(n21246) );
  NOR2X1 U20292 ( .A(n44708), .B(n44448), .Y(n21249) );
  NOR2X1 U20295 ( .A(n44642), .B(n44451), .Y(n21256) );
  NOR2X1 U20299 ( .A(n44706), .B(n44448), .Y(n21257) );
  NOR2X1 U20302 ( .A(n44648), .B(n44451), .Y(n21262) );
  NOR2X1 U20306 ( .A(n44714), .B(n44448), .Y(n21263) );
  NOR2X1 U20309 ( .A(n44650), .B(n44451), .Y(n21268) );
  NOR2X1 U20313 ( .A(n44716), .B(n44448), .Y(n21269) );
  NOR2X1 U20316 ( .A(n44672), .B(n44451), .Y(n21274) );
  NOR2X1 U20320 ( .A(n44738), .B(n44448), .Y(n21275) );
  NOR2X1 U20323 ( .A(n44664), .B(n44451), .Y(n21280) );
  NOR2X1 U20327 ( .A(n44730), .B(n44448), .Y(n21281) );
  NOR2X1 U20330 ( .A(n44674), .B(n44451), .Y(n21286) );
  NOR2X1 U20334 ( .A(n44740), .B(n44448), .Y(n21287) );
  NOR2X1 U20337 ( .A(n44676), .B(n44451), .Y(n21292) );
  NOR2X1 U20341 ( .A(n44742), .B(n44448), .Y(n21293) );
  NOR2X1 U20344 ( .A(n44656), .B(n44451), .Y(n21298) );
  NOR2X1 U20348 ( .A(n44722), .B(n44448), .Y(n21299) );
  NOR2X1 U20351 ( .A(n44658), .B(n44451), .Y(n21304) );
  NOR2X1 U20355 ( .A(n44724), .B(n44448), .Y(n21305) );
  NOR2X1 U20358 ( .A(n44662), .B(n44451), .Y(n21310) );
  NOR2X1 U20362 ( .A(n44728), .B(n44448), .Y(n21311) );
  NOR2X1 U20365 ( .A(n44654), .B(n44451), .Y(n21316) );
  NOR2X1 U20369 ( .A(n44720), .B(n44448), .Y(n21317) );
  NOR2X1 U20372 ( .A(n44652), .B(n44452), .Y(n21322) );
  NOR2X1 U20376 ( .A(n44718), .B(n44449), .Y(n21323) );
  NOR2X1 U20379 ( .A(n44666), .B(n44452), .Y(n21328) );
  NOR2X1 U20383 ( .A(n44732), .B(n44449), .Y(n21329) );
  NOR2X1 U20386 ( .A(n44678), .B(n44452), .Y(n21334) );
  NOR2X1 U20390 ( .A(n44744), .B(n44449), .Y(n21335) );
  NOR2X1 U20393 ( .A(n44660), .B(n44452), .Y(n21340) );
  NOR2X1 U20397 ( .A(n44726), .B(n44449), .Y(n21341) );
  NOR2X1 U20400 ( .A(n44644), .B(n44452), .Y(n21346) );
  NOR2X1 U20404 ( .A(n44710), .B(n44449), .Y(n21347) );
  NOR2X1 U20407 ( .A(n44646), .B(n44452), .Y(n21352) );
  NOR2X1 U20411 ( .A(n44712), .B(n44449), .Y(n21353) );
  NOR2X1 U20414 ( .A(n44670), .B(n44452), .Y(n21358) );
  NOR2X1 U20418 ( .A(n44736), .B(n44449), .Y(n21359) );
  NOR2X1 U20421 ( .A(n44668), .B(n44452), .Y(n21364) );
  NOR2X1 U20425 ( .A(n44734), .B(n44449), .Y(n21365) );
  NOR2X1 U20428 ( .A(n44694), .B(n44452), .Y(n21370) );
  NOR2X1 U20432 ( .A(n44758), .B(n44449), .Y(n21371) );
  NOR2X1 U20435 ( .A(n44698), .B(n44452), .Y(n21376) );
  NOR2X1 U20439 ( .A(n44762), .B(n44449), .Y(n21377) );
  NOR2X1 U20442 ( .A(n44700), .B(n44452), .Y(n21382) );
  NOR2X1 U20446 ( .A(n44764), .B(n44449), .Y(n21383) );
  NOR2X1 U20449 ( .A(n44704), .B(n44452), .Y(n21388) );
  NOR2X1 U20453 ( .A(n44768), .B(n44449), .Y(n21389) );
  NOR2X1 U20456 ( .A(n44702), .B(n44453), .Y(n21394) );
  NOR2X1 U20460 ( .A(n44766), .B(n44450), .Y(n21395) );
  NOR2X1 U20463 ( .A(n44696), .B(n44453), .Y(n21400) );
  NOR2X1 U20467 ( .A(n44760), .B(n44450), .Y(n21401) );
  NOR2X1 U20470 ( .A(n44692), .B(n44453), .Y(n21406) );
  NOR2X1 U20474 ( .A(n44748), .B(n44450), .Y(n21407) );
  NOR2X1 U20477 ( .A(n44690), .B(n44453), .Y(n21412) );
  NOR2X1 U20481 ( .A(n44752), .B(n44450), .Y(n21413) );
  NOR2X1 U20484 ( .A(n44688), .B(n44453), .Y(n21418) );
  NOR2X1 U20488 ( .A(n44754), .B(n44450), .Y(n21419) );
  NOR2X1 U20491 ( .A(n44686), .B(n44453), .Y(n21424) );
  NOR2X1 U20495 ( .A(n44756), .B(n44450), .Y(n21425) );
  NOR2X1 U20498 ( .A(n44684), .B(n44453), .Y(n21430) );
  NOR2X1 U20502 ( .A(n44750), .B(n44450), .Y(n21431) );
  NOR2X1 U20505 ( .A(n44682), .B(n44453), .Y(n21436) );
  NOR2X1 U20510 ( .A(n44746), .B(n44450), .Y(n21438) );
  NOR2X1 U20513 ( .A(n44679), .B(n44445), .Y(n21443) );
  NOR2X1 U20517 ( .A(n44707), .B(n44436), .Y(n21446) );
  NOR2X1 U20520 ( .A(n44641), .B(n44445), .Y(n21453) );
  NOR2X1 U20524 ( .A(n44705), .B(n44436), .Y(n21454) );
  NOR2X1 U20527 ( .A(n44647), .B(n44445), .Y(n21459) );
  NOR2X1 U20531 ( .A(n44713), .B(n44436), .Y(n21460) );
  NOR2X1 U20534 ( .A(n44649), .B(n44445), .Y(n21465) );
  NOR2X1 U20538 ( .A(n44715), .B(n44436), .Y(n21466) );
  NOR2X1 U20541 ( .A(n44671), .B(n44445), .Y(n21471) );
  NOR2X1 U20545 ( .A(n44737), .B(n44436), .Y(n21472) );
  NOR2X1 U20548 ( .A(n44663), .B(n44445), .Y(n21477) );
  NOR2X1 U20552 ( .A(n44729), .B(n44436), .Y(n21478) );
  NOR2X1 U20555 ( .A(n44673), .B(n44445), .Y(n21483) );
  NOR2X1 U20559 ( .A(n44739), .B(n44436), .Y(n21484) );
  NOR2X1 U20562 ( .A(n44675), .B(n44445), .Y(n21489) );
  NOR2X1 U20566 ( .A(n44741), .B(n44436), .Y(n21490) );
  NOR2X1 U20569 ( .A(n44655), .B(n44445), .Y(n21495) );
  NOR2X1 U20573 ( .A(n44721), .B(n44436), .Y(n21496) );
  NOR2X1 U20576 ( .A(n44657), .B(n44445), .Y(n21501) );
  NOR2X1 U20580 ( .A(n44723), .B(n44436), .Y(n21502) );
  NOR2X1 U20583 ( .A(n44661), .B(n44445), .Y(n21507) );
  NOR2X1 U20587 ( .A(n44727), .B(n44436), .Y(n21508) );
  NOR2X1 U20590 ( .A(n44653), .B(n44445), .Y(n21513) );
  NOR2X1 U20594 ( .A(n44719), .B(n44436), .Y(n21514) );
  NOR2X1 U20597 ( .A(n44651), .B(n44446), .Y(n21519) );
  NOR2X1 U20601 ( .A(n44717), .B(n44437), .Y(n21520) );
  NOR2X1 U20604 ( .A(n44665), .B(n44446), .Y(n21525) );
  NOR2X1 U20608 ( .A(n44731), .B(n44437), .Y(n21526) );
  NOR2X1 U20611 ( .A(n44677), .B(n44446), .Y(n21531) );
  NOR2X1 U20615 ( .A(n44743), .B(n44437), .Y(n21532) );
  NOR2X1 U20618 ( .A(n44659), .B(n44446), .Y(n21537) );
  NOR2X1 U20622 ( .A(n44725), .B(n44437), .Y(n21538) );
  NOR2X1 U20625 ( .A(n44643), .B(n44446), .Y(n21543) );
  NOR2X1 U20629 ( .A(n44709), .B(n44437), .Y(n21544) );
  NOR2X1 U20632 ( .A(n44645), .B(n44446), .Y(n21549) );
  NOR2X1 U20636 ( .A(n44711), .B(n44437), .Y(n21550) );
  NOR2X1 U20639 ( .A(n44669), .B(n44446), .Y(n21555) );
  NOR2X1 U20643 ( .A(n44735), .B(n44437), .Y(n21556) );
  NOR2X1 U20646 ( .A(n44667), .B(n44446), .Y(n21561) );
  NOR2X1 U20650 ( .A(n44733), .B(n44437), .Y(n21562) );
  NOR2X1 U20653 ( .A(n44694), .B(n44446), .Y(n21567) );
  NOR2X1 U20657 ( .A(n44758), .B(n44437), .Y(n21568) );
  NOR2X1 U20660 ( .A(n44698), .B(n44446), .Y(n21573) );
  NOR2X1 U20664 ( .A(n44762), .B(n44437), .Y(n21574) );
  NOR2X1 U20667 ( .A(n44700), .B(n44446), .Y(n21579) );
  NOR2X1 U20671 ( .A(n44764), .B(n44437), .Y(n21580) );
  NOR2X1 U20674 ( .A(n44704), .B(n44446), .Y(n21585) );
  NOR2X1 U20678 ( .A(n44768), .B(n44437), .Y(n21586) );
  NOR2X1 U20681 ( .A(n44702), .B(n44447), .Y(n21591) );
  NOR2X1 U20685 ( .A(n44766), .B(n44438), .Y(n21592) );
  NOR2X1 U20688 ( .A(n44696), .B(n44447), .Y(n21597) );
  NOR2X1 U20692 ( .A(n44760), .B(n44438), .Y(n21598) );
  NOR2X1 U20695 ( .A(n44692), .B(n44447), .Y(n21603) );
  NOR2X1 U20699 ( .A(n44748), .B(n44438), .Y(n21604) );
  NOR2X1 U20702 ( .A(n44690), .B(n44447), .Y(n21609) );
  NOR2X1 U20706 ( .A(n44752), .B(n44438), .Y(n21610) );
  NOR2X1 U20709 ( .A(n44688), .B(n44447), .Y(n21615) );
  NOR2X1 U20713 ( .A(n44754), .B(n44438), .Y(n21616) );
  NOR2X1 U20716 ( .A(n44686), .B(n44447), .Y(n21621) );
  NOR2X1 U20720 ( .A(n44756), .B(n44438), .Y(n21622) );
  NOR2X1 U20723 ( .A(n44684), .B(n44447), .Y(n21627) );
  NOR2X1 U20727 ( .A(n44750), .B(n44438), .Y(n21628) );
  NOR2X1 U20730 ( .A(n44682), .B(n44447), .Y(n21633) );
  NAND2X1 U20732 ( .A(n569), .B(n44441), .Y(n21445) );
  NOR2X1 U20735 ( .A(n44746), .B(n44438), .Y(n21634) );
  NOR2X1 U20738 ( .A(n44679), .B(n44433), .Y(n21639) );
  NOR2X1 U20742 ( .A(n44707), .B(n44424), .Y(n21642) );
  NOR2X1 U20745 ( .A(n44641), .B(n44433), .Y(n21649) );
  NOR2X1 U20749 ( .A(n44705), .B(n44424), .Y(n21650) );
  NOR2X1 U20752 ( .A(n44647), .B(n44433), .Y(n21655) );
  NOR2X1 U20756 ( .A(n44713), .B(n44424), .Y(n21656) );
  NOR2X1 U20759 ( .A(n44649), .B(n44433), .Y(n21661) );
  NOR2X1 U20763 ( .A(n44715), .B(n44424), .Y(n21662) );
  NOR2X1 U20766 ( .A(n44671), .B(n44433), .Y(n21667) );
  NOR2X1 U20770 ( .A(n44737), .B(n44424), .Y(n21668) );
  NOR2X1 U20773 ( .A(n44663), .B(n44433), .Y(n21673) );
  NOR2X1 U20777 ( .A(n44729), .B(n44424), .Y(n21674) );
  NOR2X1 U20780 ( .A(n44673), .B(n44433), .Y(n21679) );
  NOR2X1 U20784 ( .A(n44739), .B(n44424), .Y(n21680) );
  NOR2X1 U20787 ( .A(n44675), .B(n44433), .Y(n21685) );
  NOR2X1 U20791 ( .A(n44741), .B(n44424), .Y(n21686) );
  NOR2X1 U20794 ( .A(n44655), .B(n44433), .Y(n21691) );
  NOR2X1 U20798 ( .A(n44721), .B(n44424), .Y(n21692) );
  NOR2X1 U20801 ( .A(n44657), .B(n44433), .Y(n21697) );
  NOR2X1 U20805 ( .A(n44723), .B(n44424), .Y(n21698) );
  NOR2X1 U20808 ( .A(n44661), .B(n44433), .Y(n21703) );
  NOR2X1 U20812 ( .A(n44727), .B(n44424), .Y(n21704) );
  NOR2X1 U20815 ( .A(n44653), .B(n44433), .Y(n21709) );
  NOR2X1 U20819 ( .A(n44719), .B(n44424), .Y(n21710) );
  NOR2X1 U20822 ( .A(n44651), .B(n44434), .Y(n21715) );
  NOR2X1 U20826 ( .A(n44717), .B(n44425), .Y(n21716) );
  NOR2X1 U20829 ( .A(n44665), .B(n44434), .Y(n21721) );
  NOR2X1 U20833 ( .A(n44731), .B(n44425), .Y(n21722) );
  NOR2X1 U20836 ( .A(n44677), .B(n44434), .Y(n21727) );
  NOR2X1 U20840 ( .A(n44743), .B(n44425), .Y(n21728) );
  NOR2X1 U20843 ( .A(n44659), .B(n44434), .Y(n21733) );
  NOR2X1 U20847 ( .A(n44725), .B(n44425), .Y(n21734) );
  NOR2X1 U20850 ( .A(n44643), .B(n44434), .Y(n21739) );
  NOR2X1 U20854 ( .A(n44709), .B(n44425), .Y(n21740) );
  NOR2X1 U20857 ( .A(n44645), .B(n44434), .Y(n21745) );
  NOR2X1 U20861 ( .A(n44711), .B(n44425), .Y(n21746) );
  NOR2X1 U20864 ( .A(n44669), .B(n44434), .Y(n21751) );
  NOR2X1 U20868 ( .A(n44735), .B(n44425), .Y(n21752) );
  NOR2X1 U20871 ( .A(n44667), .B(n44434), .Y(n21757) );
  NOR2X1 U20875 ( .A(n44733), .B(n44425), .Y(n21758) );
  NOR2X1 U20878 ( .A(n44693), .B(n44434), .Y(n21763) );
  NOR2X1 U20882 ( .A(n44757), .B(n44425), .Y(n21764) );
  NOR2X1 U20885 ( .A(n44697), .B(n44434), .Y(n21769) );
  NOR2X1 U20889 ( .A(n44761), .B(n44425), .Y(n21770) );
  NOR2X1 U20892 ( .A(n44699), .B(n44434), .Y(n21775) );
  NOR2X1 U20896 ( .A(n44763), .B(n44425), .Y(n21776) );
  NOR2X1 U20899 ( .A(n44703), .B(n44434), .Y(n21781) );
  NOR2X1 U20903 ( .A(n44767), .B(n44425), .Y(n21782) );
  NOR2X1 U20906 ( .A(n44701), .B(n44435), .Y(n21787) );
  NOR2X1 U20910 ( .A(n44765), .B(n44426), .Y(n21788) );
  NOR2X1 U20913 ( .A(n44695), .B(n44435), .Y(n21793) );
  NOR2X1 U20917 ( .A(n44759), .B(n44426), .Y(n21794) );
  NOR2X1 U20920 ( .A(n44691), .B(n44435), .Y(n21799) );
  NOR2X1 U20924 ( .A(n44747), .B(n44426), .Y(n21800) );
  NOR2X1 U20927 ( .A(n44689), .B(n44435), .Y(n21805) );
  NOR2X1 U20931 ( .A(n44751), .B(n44426), .Y(n21806) );
  NOR2X1 U20934 ( .A(n44687), .B(n44435), .Y(n21811) );
  NOR2X1 U20938 ( .A(n44753), .B(n44426), .Y(n21812) );
  NOR2X1 U20941 ( .A(n44685), .B(n44435), .Y(n21817) );
  NOR2X1 U20945 ( .A(n44755), .B(n44426), .Y(n21818) );
  NOR2X1 U20948 ( .A(n44683), .B(n44435), .Y(n21823) );
  NOR2X1 U20952 ( .A(n44749), .B(n44426), .Y(n21824) );
  NOR2X1 U20955 ( .A(n44681), .B(n44435), .Y(n21829) );
  NAND2X1 U20957 ( .A(n529), .B(n44429), .Y(n21641) );
  NOR2X1 U20960 ( .A(n44745), .B(n44426), .Y(n21830) );
  NOR2X1 U20963 ( .A(n44679), .B(n44421), .Y(n21835) );
  NOR2X1 U20967 ( .A(n44707), .B(n44412), .Y(n21838) );
  NOR2X1 U20970 ( .A(n44641), .B(n44421), .Y(n21845) );
  NOR2X1 U20974 ( .A(n44705), .B(n44412), .Y(n21846) );
  NOR2X1 U20977 ( .A(n44647), .B(n44421), .Y(n21851) );
  NOR2X1 U20981 ( .A(n44713), .B(n44412), .Y(n21852) );
  NOR2X1 U20984 ( .A(n44649), .B(n44421), .Y(n21857) );
  NOR2X1 U20988 ( .A(n44715), .B(n44412), .Y(n21858) );
  NOR2X1 U20991 ( .A(n44671), .B(n44421), .Y(n21863) );
  NOR2X1 U20995 ( .A(n44737), .B(n44412), .Y(n21864) );
  NOR2X1 U20998 ( .A(n44663), .B(n44421), .Y(n21869) );
  NOR2X1 U21002 ( .A(n44729), .B(n44412), .Y(n21870) );
  NOR2X1 U21005 ( .A(n44673), .B(n44421), .Y(n21875) );
  NOR2X1 U21009 ( .A(n44739), .B(n44412), .Y(n21876) );
  NOR2X1 U21012 ( .A(n44675), .B(n44421), .Y(n21881) );
  NOR2X1 U21016 ( .A(n44741), .B(n44412), .Y(n21882) );
  NOR2X1 U21019 ( .A(n44655), .B(n44421), .Y(n21887) );
  NOR2X1 U21023 ( .A(n44721), .B(n44412), .Y(n21888) );
  NOR2X1 U21026 ( .A(n44657), .B(n44421), .Y(n21893) );
  NOR2X1 U21030 ( .A(n44723), .B(n44412), .Y(n21894) );
  NOR2X1 U21033 ( .A(n44661), .B(n44421), .Y(n21899) );
  NOR2X1 U21037 ( .A(n44727), .B(n44412), .Y(n21900) );
  NOR2X1 U21040 ( .A(n44653), .B(n44421), .Y(n21905) );
  NOR2X1 U21044 ( .A(n44719), .B(n44412), .Y(n21906) );
  NOR2X1 U21047 ( .A(n44651), .B(n44422), .Y(n21911) );
  NOR2X1 U21051 ( .A(n44717), .B(n44413), .Y(n21912) );
  NOR2X1 U21054 ( .A(n44665), .B(n44422), .Y(n21917) );
  NOR2X1 U21058 ( .A(n44731), .B(n44413), .Y(n21918) );
  NOR2X1 U21061 ( .A(n44677), .B(n44422), .Y(n21923) );
  NOR2X1 U21065 ( .A(n44743), .B(n44413), .Y(n21924) );
  NOR2X1 U21068 ( .A(n44659), .B(n44422), .Y(n21929) );
  NOR2X1 U21072 ( .A(n44725), .B(n44413), .Y(n21930) );
  NOR2X1 U21075 ( .A(n44643), .B(n44422), .Y(n21935) );
  NOR2X1 U21079 ( .A(n44709), .B(n44413), .Y(n21936) );
  NOR2X1 U21082 ( .A(n44645), .B(n44422), .Y(n21941) );
  NOR2X1 U21086 ( .A(n44711), .B(n44413), .Y(n21942) );
  NOR2X1 U21089 ( .A(n44669), .B(n44422), .Y(n21947) );
  NOR2X1 U21093 ( .A(n44735), .B(n44413), .Y(n21948) );
  NOR2X1 U21096 ( .A(n44667), .B(n44422), .Y(n21953) );
  NOR2X1 U21100 ( .A(n44733), .B(n44413), .Y(n21954) );
  NOR2X1 U21103 ( .A(n44693), .B(n44422), .Y(n21959) );
  NOR2X1 U21107 ( .A(n44757), .B(n44413), .Y(n21960) );
  NOR2X1 U21110 ( .A(n44697), .B(n44422), .Y(n21965) );
  NOR2X1 U21114 ( .A(n44761), .B(n44413), .Y(n21966) );
  NOR2X1 U21117 ( .A(n44699), .B(n44422), .Y(n21971) );
  NOR2X1 U21121 ( .A(n44763), .B(n44413), .Y(n21972) );
  NOR2X1 U21124 ( .A(n44703), .B(n44422), .Y(n21977) );
  NOR2X1 U21128 ( .A(n44767), .B(n44413), .Y(n21978) );
  NOR2X1 U21131 ( .A(n44701), .B(n44423), .Y(n21983) );
  NOR2X1 U21135 ( .A(n44765), .B(n44414), .Y(n21984) );
  NOR2X1 U21138 ( .A(n44695), .B(n44423), .Y(n21989) );
  NOR2X1 U21142 ( .A(n44759), .B(n44414), .Y(n21990) );
  NOR2X1 U21145 ( .A(n44691), .B(n44423), .Y(n21995) );
  NOR2X1 U21149 ( .A(n44747), .B(n44414), .Y(n21996) );
  NOR2X1 U21152 ( .A(n44689), .B(n44423), .Y(n22001) );
  NOR2X1 U21156 ( .A(n44751), .B(n44414), .Y(n22002) );
  NOR2X1 U21159 ( .A(n44687), .B(n44423), .Y(n22007) );
  NOR2X1 U21163 ( .A(n44753), .B(n44414), .Y(n22008) );
  NOR2X1 U21166 ( .A(n44685), .B(n44423), .Y(n22013) );
  NOR2X1 U21170 ( .A(n44755), .B(n44414), .Y(n22014) );
  NOR2X1 U21173 ( .A(n44683), .B(n44423), .Y(n22019) );
  NOR2X1 U21177 ( .A(n44749), .B(n44414), .Y(n22020) );
  NOR2X1 U21180 ( .A(n44681), .B(n44423), .Y(n22025) );
  NAND2X1 U21182 ( .A(n571), .B(n44417), .Y(n21837) );
  NOR2X1 U21185 ( .A(n44745), .B(n44414), .Y(n22026) );
  NOR2X1 U21188 ( .A(n44679), .B(n44409), .Y(n22031) );
  NOR2X1 U21192 ( .A(n44707), .B(n44400), .Y(n22034) );
  NOR2X1 U21195 ( .A(n44641), .B(n44409), .Y(n22041) );
  NOR2X1 U21199 ( .A(n44705), .B(n44400), .Y(n22042) );
  NOR2X1 U21202 ( .A(n44647), .B(n44409), .Y(n22047) );
  NOR2X1 U21206 ( .A(n44713), .B(n44400), .Y(n22048) );
  NOR2X1 U21209 ( .A(n44649), .B(n44409), .Y(n22053) );
  NOR2X1 U21213 ( .A(n44715), .B(n44400), .Y(n22054) );
  NOR2X1 U21216 ( .A(n44671), .B(n44409), .Y(n22059) );
  NOR2X1 U21220 ( .A(n44737), .B(n44400), .Y(n22060) );
  NOR2X1 U21223 ( .A(n44663), .B(n44409), .Y(n22065) );
  NOR2X1 U21227 ( .A(n44729), .B(n44400), .Y(n22066) );
  NOR2X1 U21230 ( .A(n44673), .B(n44409), .Y(n22071) );
  NOR2X1 U21234 ( .A(n44739), .B(n44400), .Y(n22072) );
  NOR2X1 U21237 ( .A(n44675), .B(n44409), .Y(n22077) );
  NOR2X1 U21241 ( .A(n44741), .B(n44400), .Y(n22078) );
  NOR2X1 U21244 ( .A(n44655), .B(n44409), .Y(n22083) );
  NOR2X1 U21248 ( .A(n44721), .B(n44400), .Y(n22084) );
  NOR2X1 U21251 ( .A(n44657), .B(n44409), .Y(n22089) );
  NOR2X1 U21255 ( .A(n44723), .B(n44400), .Y(n22090) );
  NOR2X1 U21258 ( .A(n44661), .B(n44409), .Y(n22095) );
  NOR2X1 U21262 ( .A(n44727), .B(n44400), .Y(n22096) );
  NOR2X1 U21265 ( .A(n44653), .B(n44409), .Y(n22101) );
  NOR2X1 U21269 ( .A(n44719), .B(n44400), .Y(n22102) );
  NOR2X1 U21272 ( .A(n44651), .B(n44410), .Y(n22107) );
  NOR2X1 U21276 ( .A(n44717), .B(n44401), .Y(n22108) );
  NOR2X1 U21279 ( .A(n44665), .B(n44410), .Y(n22113) );
  NOR2X1 U21283 ( .A(n44731), .B(n44401), .Y(n22114) );
  NOR2X1 U21286 ( .A(n44677), .B(n44410), .Y(n22119) );
  NOR2X1 U21290 ( .A(n44743), .B(n44401), .Y(n22120) );
  NOR2X1 U21293 ( .A(n44659), .B(n44410), .Y(n22125) );
  NOR2X1 U21297 ( .A(n44725), .B(n44401), .Y(n22126) );
  NOR2X1 U21300 ( .A(n44643), .B(n44410), .Y(n22131) );
  NOR2X1 U21304 ( .A(n44709), .B(n44401), .Y(n22132) );
  NOR2X1 U21307 ( .A(n44645), .B(n44410), .Y(n22137) );
  NOR2X1 U21311 ( .A(n44711), .B(n44401), .Y(n22138) );
  NOR2X1 U21314 ( .A(n44669), .B(n44410), .Y(n22143) );
  NOR2X1 U21318 ( .A(n44735), .B(n44401), .Y(n22144) );
  NOR2X1 U21321 ( .A(n44667), .B(n44410), .Y(n22149) );
  NOR2X1 U21325 ( .A(n44733), .B(n44401), .Y(n22150) );
  NOR2X1 U21328 ( .A(n44693), .B(n44410), .Y(n22155) );
  NOR2X1 U21332 ( .A(n44757), .B(n44401), .Y(n22156) );
  NOR2X1 U21335 ( .A(n44697), .B(n44410), .Y(n22161) );
  NOR2X1 U21339 ( .A(n44761), .B(n44401), .Y(n22162) );
  NOR2X1 U21342 ( .A(n44699), .B(n44410), .Y(n22167) );
  NOR2X1 U21346 ( .A(n44763), .B(n44401), .Y(n22168) );
  NOR2X1 U21349 ( .A(n44703), .B(n44410), .Y(n22173) );
  NOR2X1 U21353 ( .A(n44767), .B(n44401), .Y(n22174) );
  NOR2X1 U21356 ( .A(n44701), .B(n44411), .Y(n22179) );
  NOR2X1 U21360 ( .A(n44765), .B(n44402), .Y(n22180) );
  NOR2X1 U21363 ( .A(n44695), .B(n44411), .Y(n22185) );
  NOR2X1 U21367 ( .A(n44759), .B(n44402), .Y(n22186) );
  NOR2X1 U21370 ( .A(n44691), .B(n44411), .Y(n22191) );
  NOR2X1 U21374 ( .A(n44747), .B(n44402), .Y(n22192) );
  NOR2X1 U21377 ( .A(n44689), .B(n44411), .Y(n22197) );
  NOR2X1 U21381 ( .A(n44751), .B(n44402), .Y(n22198) );
  NOR2X1 U21384 ( .A(n44687), .B(n44411), .Y(n22203) );
  NOR2X1 U21388 ( .A(n44753), .B(n44402), .Y(n22204) );
  NOR2X1 U21391 ( .A(n44685), .B(n44411), .Y(n22209) );
  NOR2X1 U21395 ( .A(n44755), .B(n44402), .Y(n22210) );
  NOR2X1 U21398 ( .A(n44683), .B(n44411), .Y(n22215) );
  NOR2X1 U21402 ( .A(n44749), .B(n44402), .Y(n22216) );
  NOR2X1 U21405 ( .A(n44681), .B(n44411), .Y(n22221) );
  NAND2X1 U21407 ( .A(n527), .B(n44405), .Y(n22033) );
  NOR2X1 U21410 ( .A(n44745), .B(n44402), .Y(n22222) );
  NOR2X1 U21413 ( .A(n44679), .B(n44397), .Y(n22227) );
  NOR2X1 U21417 ( .A(n44707), .B(n44388), .Y(n22230) );
  NOR2X1 U21420 ( .A(n44641), .B(n44397), .Y(n22237) );
  NOR2X1 U21424 ( .A(n44705), .B(n44388), .Y(n22238) );
  NOR2X1 U21427 ( .A(n44647), .B(n44397), .Y(n22243) );
  NOR2X1 U21431 ( .A(n44713), .B(n44388), .Y(n22244) );
  NOR2X1 U21434 ( .A(n44649), .B(n44397), .Y(n22249) );
  NOR2X1 U21438 ( .A(n44715), .B(n44388), .Y(n22250) );
  NOR2X1 U21441 ( .A(n44671), .B(n44397), .Y(n22255) );
  NOR2X1 U21445 ( .A(n44737), .B(n44388), .Y(n22256) );
  NOR2X1 U21448 ( .A(n44663), .B(n44397), .Y(n22261) );
  NOR2X1 U21452 ( .A(n44729), .B(n44388), .Y(n22262) );
  NOR2X1 U21455 ( .A(n44673), .B(n44397), .Y(n22267) );
  NOR2X1 U21459 ( .A(n44739), .B(n44388), .Y(n22268) );
  NOR2X1 U21462 ( .A(n44675), .B(n44397), .Y(n22273) );
  NOR2X1 U21466 ( .A(n44741), .B(n44388), .Y(n22274) );
  NOR2X1 U21469 ( .A(n44655), .B(n44397), .Y(n22279) );
  NOR2X1 U21473 ( .A(n44721), .B(n44388), .Y(n22280) );
  NOR2X1 U21476 ( .A(n44657), .B(n44397), .Y(n22285) );
  NOR2X1 U21480 ( .A(n44723), .B(n44388), .Y(n22286) );
  NOR2X1 U21483 ( .A(n44661), .B(n44397), .Y(n22291) );
  NOR2X1 U21487 ( .A(n44727), .B(n44388), .Y(n22292) );
  NOR2X1 U21490 ( .A(n44653), .B(n44397), .Y(n22297) );
  NOR2X1 U21494 ( .A(n44719), .B(n44388), .Y(n22298) );
  NOR2X1 U21497 ( .A(n44651), .B(n44398), .Y(n22303) );
  NOR2X1 U21501 ( .A(n44717), .B(n44389), .Y(n22304) );
  NOR2X1 U21504 ( .A(n44665), .B(n44398), .Y(n22309) );
  NOR2X1 U21508 ( .A(n44731), .B(n44389), .Y(n22310) );
  NOR2X1 U21511 ( .A(n44677), .B(n44398), .Y(n22315) );
  NOR2X1 U21515 ( .A(n44743), .B(n44389), .Y(n22316) );
  NOR2X1 U21518 ( .A(n44659), .B(n44398), .Y(n22321) );
  NOR2X1 U21522 ( .A(n44725), .B(n44389), .Y(n22322) );
  NOR2X1 U21525 ( .A(n44643), .B(n44398), .Y(n22327) );
  NOR2X1 U21529 ( .A(n44709), .B(n44389), .Y(n22328) );
  NOR2X1 U21532 ( .A(n44645), .B(n44398), .Y(n22333) );
  NOR2X1 U21536 ( .A(n44711), .B(n44389), .Y(n22334) );
  NOR2X1 U21539 ( .A(n44669), .B(n44398), .Y(n22339) );
  NOR2X1 U21543 ( .A(n44735), .B(n44389), .Y(n22340) );
  NOR2X1 U21546 ( .A(n44667), .B(n44398), .Y(n22345) );
  NOR2X1 U21550 ( .A(n44733), .B(n44389), .Y(n22346) );
  NOR2X1 U21553 ( .A(n44693), .B(n44398), .Y(n22351) );
  NOR2X1 U21557 ( .A(n44757), .B(n44389), .Y(n22352) );
  NOR2X1 U21560 ( .A(n44697), .B(n44398), .Y(n22357) );
  NOR2X1 U21564 ( .A(n44761), .B(n44389), .Y(n22358) );
  NOR2X1 U21567 ( .A(n44699), .B(n44398), .Y(n22363) );
  NOR2X1 U21571 ( .A(n44763), .B(n44389), .Y(n22364) );
  NOR2X1 U21574 ( .A(n44703), .B(n44398), .Y(n22369) );
  NOR2X1 U21578 ( .A(n44767), .B(n44389), .Y(n22370) );
  NOR2X1 U21581 ( .A(n44701), .B(n44399), .Y(n22375) );
  NOR2X1 U21585 ( .A(n44765), .B(n44390), .Y(n22376) );
  NOR2X1 U21588 ( .A(n44695), .B(n44399), .Y(n22381) );
  NOR2X1 U21592 ( .A(n44759), .B(n44390), .Y(n22382) );
  NOR2X1 U21595 ( .A(n44691), .B(n44399), .Y(n22387) );
  NOR2X1 U21599 ( .A(n44747), .B(n44390), .Y(n22388) );
  NOR2X1 U21602 ( .A(n44689), .B(n44399), .Y(n22393) );
  NOR2X1 U21606 ( .A(n44751), .B(n44390), .Y(n22394) );
  NOR2X1 U21609 ( .A(n44687), .B(n44399), .Y(n22399) );
  NOR2X1 U21613 ( .A(n44753), .B(n44390), .Y(n22400) );
  NOR2X1 U21616 ( .A(n44685), .B(n44399), .Y(n22405) );
  NOR2X1 U21620 ( .A(n44755), .B(n44390), .Y(n22406) );
  NOR2X1 U21623 ( .A(n44683), .B(n44399), .Y(n22411) );
  NOR2X1 U21627 ( .A(n44749), .B(n44390), .Y(n22412) );
  NOR2X1 U21630 ( .A(n44681), .B(n44399), .Y(n22417) );
  NAND2X1 U21632 ( .A(n567), .B(n44393), .Y(n22229) );
  NOR2X1 U21635 ( .A(n44745), .B(n44390), .Y(n22418) );
  NOR2X1 U21638 ( .A(n44679), .B(n44385), .Y(n22423) );
  NOR2X1 U21642 ( .A(n44707), .B(n44376), .Y(n22426) );
  NOR2X1 U21645 ( .A(n44641), .B(n44385), .Y(n22433) );
  NOR2X1 U21649 ( .A(n44705), .B(n44376), .Y(n22434) );
  NOR2X1 U21652 ( .A(n44647), .B(n44385), .Y(n22439) );
  NOR2X1 U21656 ( .A(n44713), .B(n44376), .Y(n22440) );
  NOR2X1 U21659 ( .A(n44649), .B(n44385), .Y(n22445) );
  NOR2X1 U21663 ( .A(n44715), .B(n44376), .Y(n22446) );
  NOR2X1 U21666 ( .A(n44671), .B(n44385), .Y(n22451) );
  NOR2X1 U21670 ( .A(n44737), .B(n44376), .Y(n22452) );
  NOR2X1 U21673 ( .A(n44663), .B(n44385), .Y(n22457) );
  NOR2X1 U21677 ( .A(n44729), .B(n44376), .Y(n22458) );
  NOR2X1 U21680 ( .A(n44673), .B(n44385), .Y(n22463) );
  NOR2X1 U21684 ( .A(n44739), .B(n44376), .Y(n22464) );
  NOR2X1 U21687 ( .A(n44675), .B(n44385), .Y(n22469) );
  NOR2X1 U21691 ( .A(n44741), .B(n44376), .Y(n22470) );
  NOR2X1 U21694 ( .A(n44655), .B(n44385), .Y(n22475) );
  NOR2X1 U21698 ( .A(n44721), .B(n44376), .Y(n22476) );
  NOR2X1 U21701 ( .A(n44657), .B(n44385), .Y(n22481) );
  NOR2X1 U21705 ( .A(n44723), .B(n44376), .Y(n22482) );
  NOR2X1 U21708 ( .A(n44661), .B(n44385), .Y(n22487) );
  NOR2X1 U21712 ( .A(n44727), .B(n44376), .Y(n22488) );
  NOR2X1 U21715 ( .A(n44653), .B(n44385), .Y(n22493) );
  NOR2X1 U21719 ( .A(n44719), .B(n44376), .Y(n22494) );
  NOR2X1 U21722 ( .A(n44651), .B(n44386), .Y(n22499) );
  NOR2X1 U21726 ( .A(n44717), .B(n44377), .Y(n22500) );
  NOR2X1 U21729 ( .A(n44665), .B(n44386), .Y(n22505) );
  NOR2X1 U21733 ( .A(n44731), .B(n44377), .Y(n22506) );
  NOR2X1 U21736 ( .A(n44677), .B(n44386), .Y(n22511) );
  NOR2X1 U21740 ( .A(n44743), .B(n44377), .Y(n22512) );
  NOR2X1 U21743 ( .A(n44659), .B(n44386), .Y(n22517) );
  NOR2X1 U21747 ( .A(n44725), .B(n44377), .Y(n22518) );
  NOR2X1 U21750 ( .A(n44643), .B(n44386), .Y(n22523) );
  NOR2X1 U21754 ( .A(n44709), .B(n44377), .Y(n22524) );
  NOR2X1 U21757 ( .A(n44645), .B(n44386), .Y(n22529) );
  NOR2X1 U21761 ( .A(n44711), .B(n44377), .Y(n22530) );
  NOR2X1 U21764 ( .A(n44669), .B(n44386), .Y(n22535) );
  NOR2X1 U21768 ( .A(n44735), .B(n44377), .Y(n22536) );
  NOR2X1 U21771 ( .A(n44667), .B(n44386), .Y(n22541) );
  NOR2X1 U21775 ( .A(n44733), .B(n44377), .Y(n22542) );
  NOR2X1 U21778 ( .A(n44693), .B(n44386), .Y(n22547) );
  NOR2X1 U21782 ( .A(n44757), .B(n44377), .Y(n22548) );
  NOR2X1 U21785 ( .A(n44697), .B(n44386), .Y(n22553) );
  NOR2X1 U21789 ( .A(n44761), .B(n44377), .Y(n22554) );
  NOR2X1 U21792 ( .A(n44699), .B(n44386), .Y(n22559) );
  NOR2X1 U21796 ( .A(n44763), .B(n44377), .Y(n22560) );
  NOR2X1 U21799 ( .A(n44703), .B(n44386), .Y(n22565) );
  NOR2X1 U21803 ( .A(n44767), .B(n44377), .Y(n22566) );
  NOR2X1 U21806 ( .A(n44701), .B(n44387), .Y(n22571) );
  NOR2X1 U21810 ( .A(n44765), .B(n44378), .Y(n22572) );
  NOR2X1 U21813 ( .A(n44695), .B(n44387), .Y(n22577) );
  NOR2X1 U21817 ( .A(n44759), .B(n44378), .Y(n22578) );
  NOR2X1 U21820 ( .A(n44691), .B(n44387), .Y(n22583) );
  NOR2X1 U21824 ( .A(n44747), .B(n44378), .Y(n22584) );
  NOR2X1 U21827 ( .A(n44689), .B(n44387), .Y(n22589) );
  NOR2X1 U21831 ( .A(n44751), .B(n44378), .Y(n22590) );
  NOR2X1 U21834 ( .A(n44687), .B(n44387), .Y(n22595) );
  NOR2X1 U21838 ( .A(n44753), .B(n44378), .Y(n22596) );
  NOR2X1 U21841 ( .A(n44685), .B(n44387), .Y(n22601) );
  NOR2X1 U21845 ( .A(n44755), .B(n44378), .Y(n22602) );
  NOR2X1 U21848 ( .A(n44683), .B(n44387), .Y(n22607) );
  NOR2X1 U21852 ( .A(n44749), .B(n44378), .Y(n22608) );
  NOR2X1 U21855 ( .A(n44681), .B(n44387), .Y(n22613) );
  NAND2X1 U21857 ( .A(n525), .B(n44381), .Y(n22425) );
  NOR2X1 U21860 ( .A(n44745), .B(n44378), .Y(n22614) );
  NOR2X1 U21863 ( .A(n44707), .B(n44373), .Y(n22619) );
  NOR2X1 U21867 ( .A(n44679), .B(n44370), .Y(n22622) );
  NOR2X1 U21870 ( .A(n44705), .B(n44373), .Y(n22629) );
  NOR2X1 U21874 ( .A(n44641), .B(n44370), .Y(n22630) );
  NOR2X1 U21877 ( .A(n44713), .B(n44373), .Y(n22635) );
  NOR2X1 U21881 ( .A(n44647), .B(n44370), .Y(n22636) );
  NOR2X1 U21884 ( .A(n44715), .B(n44373), .Y(n22641) );
  NOR2X1 U21888 ( .A(n44649), .B(n44370), .Y(n22642) );
  NOR2X1 U21891 ( .A(n44737), .B(n44373), .Y(n22647) );
  NOR2X1 U21895 ( .A(n44671), .B(n44370), .Y(n22648) );
  NOR2X1 U21898 ( .A(n44729), .B(n44373), .Y(n22653) );
  NOR2X1 U21902 ( .A(n44663), .B(n44370), .Y(n22654) );
  NOR2X1 U21905 ( .A(n44739), .B(n44373), .Y(n22659) );
  NOR2X1 U21909 ( .A(n44673), .B(n44370), .Y(n22660) );
  NOR2X1 U21912 ( .A(n44680), .B(n44367), .Y(n22665) );
  NOR2X1 U21916 ( .A(n44708), .B(n44358), .Y(n22668) );
  NOR2X1 U21919 ( .A(n44642), .B(n44367), .Y(n22675) );
  NOR2X1 U21923 ( .A(n44706), .B(n44358), .Y(n22676) );
  NOR2X1 U21926 ( .A(n44741), .B(n44373), .Y(n22681) );
  NOR2X1 U21930 ( .A(n44675), .B(n44370), .Y(n22682) );
  NOR2X1 U21933 ( .A(n44648), .B(n44367), .Y(n22687) );
  NOR2X1 U21937 ( .A(n44714), .B(n44358), .Y(n22688) );
  NOR2X1 U21940 ( .A(n44650), .B(n44367), .Y(n22693) );
  NOR2X1 U21944 ( .A(n44716), .B(n44358), .Y(n22694) );
  NOR2X1 U21947 ( .A(n44672), .B(n44367), .Y(n22699) );
  NOR2X1 U21951 ( .A(n44738), .B(n44358), .Y(n22700) );
  NOR2X1 U21954 ( .A(n44664), .B(n44367), .Y(n22705) );
  NOR2X1 U21958 ( .A(n44730), .B(n44358), .Y(n22706) );
  NOR2X1 U21961 ( .A(n44674), .B(n44367), .Y(n22711) );
  NOR2X1 U21965 ( .A(n44740), .B(n44358), .Y(n22712) );
  NOR2X1 U21968 ( .A(n44676), .B(n44367), .Y(n22717) );
  NOR2X1 U21972 ( .A(n44742), .B(n44358), .Y(n22718) );
  NOR2X1 U21975 ( .A(n44655), .B(n44367), .Y(n22723) );
  NOR2X1 U21979 ( .A(n44721), .B(n44358), .Y(n22724) );
  NOR2X1 U21982 ( .A(n44657), .B(n44367), .Y(n22729) );
  NOR2X1 U21986 ( .A(n44723), .B(n44358), .Y(n22730) );
  NOR2X1 U21989 ( .A(n44661), .B(n44367), .Y(n22735) );
  NOR2X1 U21993 ( .A(n44727), .B(n44358), .Y(n22736) );
  NOR2X1 U21996 ( .A(n44653), .B(n44367), .Y(n22741) );
  NOR2X1 U22000 ( .A(n44719), .B(n44358), .Y(n22742) );
  NOR2X1 U22003 ( .A(n44722), .B(n44373), .Y(n22747) );
  NOR2X1 U22007 ( .A(n44656), .B(n44370), .Y(n22748) );
  NOR2X1 U22010 ( .A(n44651), .B(n44368), .Y(n22753) );
  NOR2X1 U22014 ( .A(n44717), .B(n44359), .Y(n22754) );
  NOR2X1 U22017 ( .A(n44665), .B(n44368), .Y(n22759) );
  NOR2X1 U22021 ( .A(n44731), .B(n44359), .Y(n22760) );
  NOR2X1 U22024 ( .A(n44677), .B(n44368), .Y(n22765) );
  NOR2X1 U22028 ( .A(n44743), .B(n44359), .Y(n22766) );
  NOR2X1 U22031 ( .A(n44659), .B(n44368), .Y(n22771) );
  NOR2X1 U22035 ( .A(n44725), .B(n44359), .Y(n22772) );
  NOR2X1 U22038 ( .A(n44643), .B(n44368), .Y(n22777) );
  NOR2X1 U22042 ( .A(n44709), .B(n44359), .Y(n22778) );
  NOR2X1 U22045 ( .A(n44645), .B(n44368), .Y(n22783) );
  NOR2X1 U22049 ( .A(n44711), .B(n44359), .Y(n22784) );
  NOR2X1 U22052 ( .A(n44669), .B(n44368), .Y(n22789) );
  NOR2X1 U22056 ( .A(n44735), .B(n44359), .Y(n22790) );
  NOR2X1 U22059 ( .A(n44667), .B(n44368), .Y(n22795) );
  NOR2X1 U22063 ( .A(n44733), .B(n44359), .Y(n22796) );
  NOR2X1 U22066 ( .A(n44693), .B(n44368), .Y(n22801) );
  NOR2X1 U22070 ( .A(n44757), .B(n44359), .Y(n22802) );
  NOR2X1 U22073 ( .A(n44697), .B(n44368), .Y(n22807) );
  NOR2X1 U22077 ( .A(n44761), .B(n44359), .Y(n22808) );
  NOR2X1 U22080 ( .A(n44724), .B(n44373), .Y(n22813) );
  NOR2X1 U22084 ( .A(n44658), .B(n44370), .Y(n22814) );
  NOR2X1 U22087 ( .A(n44699), .B(n44368), .Y(n22819) );
  NOR2X1 U22091 ( .A(n44763), .B(n44359), .Y(n22820) );
  NOR2X1 U22094 ( .A(n44703), .B(n44368), .Y(n22825) );
  NOR2X1 U22098 ( .A(n44767), .B(n44359), .Y(n22826) );
  NOR2X1 U22101 ( .A(n44701), .B(n44369), .Y(n22831) );
  NOR2X1 U22105 ( .A(n44765), .B(n44360), .Y(n22832) );
  NOR2X1 U22108 ( .A(n44695), .B(n44369), .Y(n22837) );
  NOR2X1 U22112 ( .A(n44759), .B(n44360), .Y(n22838) );
  NOR2X1 U22115 ( .A(n44691), .B(n44369), .Y(n22843) );
  NOR2X1 U22119 ( .A(n44747), .B(n44360), .Y(n22844) );
  NOR2X1 U22122 ( .A(n44689), .B(n44369), .Y(n22849) );
  NOR2X1 U22126 ( .A(n44751), .B(n44360), .Y(n22850) );
  NOR2X1 U22129 ( .A(n44687), .B(n44369), .Y(n22855) );
  NOR2X1 U22133 ( .A(n44753), .B(n44360), .Y(n22856) );
  NOR2X1 U22136 ( .A(n44685), .B(n44369), .Y(n22861) );
  NOR2X1 U22140 ( .A(n44755), .B(n44360), .Y(n22862) );
  NOR2X1 U22143 ( .A(n44683), .B(n44369), .Y(n22867) );
  NOR2X1 U22147 ( .A(n44749), .B(n44360), .Y(n22868) );
  NOR2X1 U22150 ( .A(n44681), .B(n44369), .Y(n22873) );
  NAND2X1 U22152 ( .A(n553), .B(n44363), .Y(n22667) );
  NOR2X1 U22155 ( .A(n44745), .B(n44360), .Y(n22874) );
  NOR2X1 U22158 ( .A(n44728), .B(n44373), .Y(n22879) );
  NOR2X1 U22162 ( .A(n44662), .B(n44370), .Y(n22880) );
  NOR2X1 U22165 ( .A(n44679), .B(n44355), .Y(n22885) );
  NOR2X1 U22169 ( .A(n44707), .B(n44346), .Y(n22888) );
  NOR2X1 U22172 ( .A(n44641), .B(n44355), .Y(n22895) );
  NOR2X1 U22176 ( .A(n44705), .B(n44346), .Y(n22896) );
  NOR2X1 U22179 ( .A(n44647), .B(n44355), .Y(n22901) );
  NOR2X1 U22183 ( .A(n44713), .B(n44346), .Y(n22902) );
  NOR2X1 U22186 ( .A(n44649), .B(n44355), .Y(n22907) );
  NOR2X1 U22190 ( .A(n44715), .B(n44346), .Y(n22908) );
  NOR2X1 U22193 ( .A(n44671), .B(n44355), .Y(n22913) );
  NOR2X1 U22197 ( .A(n44737), .B(n44346), .Y(n22914) );
  NOR2X1 U22200 ( .A(n44720), .B(n44373), .Y(n22919) );
  NOR2X1 U22204 ( .A(n44654), .B(n44370), .Y(n22920) );
  NOR2X1 U22207 ( .A(n44663), .B(n44355), .Y(n22925) );
  NOR2X1 U22211 ( .A(n44729), .B(n44346), .Y(n22926) );
  NOR2X1 U22214 ( .A(n44673), .B(n44355), .Y(n22931) );
  NOR2X1 U22218 ( .A(n44739), .B(n44346), .Y(n22932) );
  NOR2X1 U22221 ( .A(n44675), .B(n44355), .Y(n22937) );
  NOR2X1 U22225 ( .A(n44741), .B(n44346), .Y(n22938) );
  NOR2X1 U22228 ( .A(n44655), .B(n44355), .Y(n22943) );
  NOR2X1 U22232 ( .A(n44721), .B(n44346), .Y(n22944) );
  NOR2X1 U22235 ( .A(n44657), .B(n44355), .Y(n22949) );
  NOR2X1 U22239 ( .A(n44723), .B(n44346), .Y(n22950) );
  NOR2X1 U22242 ( .A(n44661), .B(n44355), .Y(n22955) );
  NOR2X1 U22246 ( .A(n44727), .B(n44346), .Y(n22956) );
  NOR2X1 U22249 ( .A(n44653), .B(n44355), .Y(n22961) );
  NOR2X1 U22253 ( .A(n44719), .B(n44346), .Y(n22962) );
  NOR2X1 U22256 ( .A(n44652), .B(n44356), .Y(n22967) );
  NOR2X1 U22260 ( .A(n44718), .B(n44347), .Y(n22968) );
  NOR2X1 U22263 ( .A(n44666), .B(n44356), .Y(n22973) );
  NOR2X1 U22267 ( .A(n44732), .B(n44347), .Y(n22974) );
  NOR2X1 U22270 ( .A(n44678), .B(n44356), .Y(n22979) );
  NOR2X1 U22274 ( .A(n44744), .B(n44347), .Y(n22980) );
  NOR2X1 U22277 ( .A(n44717), .B(n44374), .Y(n22985) );
  NOR2X1 U22281 ( .A(n44651), .B(n44371), .Y(n22986) );
  NOR2X1 U22284 ( .A(n44660), .B(n44356), .Y(n22991) );
  NOR2X1 U22288 ( .A(n44726), .B(n44347), .Y(n22992) );
  NOR2X1 U22291 ( .A(n44644), .B(n44356), .Y(n22997) );
  NOR2X1 U22295 ( .A(n44710), .B(n44347), .Y(n22998) );
  NOR2X1 U22298 ( .A(n44646), .B(n44356), .Y(n23003) );
  NOR2X1 U22302 ( .A(n44712), .B(n44347), .Y(n23004) );
  NOR2X1 U22305 ( .A(n44670), .B(n44356), .Y(n23009) );
  NOR2X1 U22309 ( .A(n44736), .B(n44347), .Y(n23010) );
  NOR2X1 U22312 ( .A(n44668), .B(n44356), .Y(n23015) );
  NOR2X1 U22316 ( .A(n44734), .B(n44347), .Y(n23016) );
  NOR2X1 U22319 ( .A(n44693), .B(n44356), .Y(n23021) );
  NOR2X1 U22323 ( .A(n44757), .B(n44347), .Y(n23022) );
  NOR2X1 U22326 ( .A(n44697), .B(n44356), .Y(n23027) );
  NOR2X1 U22330 ( .A(n44761), .B(n44347), .Y(n23028) );
  NOR2X1 U22333 ( .A(n44699), .B(n44356), .Y(n23033) );
  NOR2X1 U22337 ( .A(n44763), .B(n44347), .Y(n23034) );
  NOR2X1 U22340 ( .A(n44703), .B(n44356), .Y(n23039) );
  NOR2X1 U22344 ( .A(n44767), .B(n44347), .Y(n23040) );
  NOR2X1 U22347 ( .A(n44701), .B(n44357), .Y(n23045) );
  NOR2X1 U22351 ( .A(n44765), .B(n44348), .Y(n23046) );
  NOR2X1 U22354 ( .A(n44731), .B(n44374), .Y(n23051) );
  NOR2X1 U22358 ( .A(n44665), .B(n44371), .Y(n23052) );
  NOR2X1 U22361 ( .A(n44695), .B(n44357), .Y(n23057) );
  NOR2X1 U22365 ( .A(n44759), .B(n44348), .Y(n23058) );
  NOR2X1 U22368 ( .A(n44691), .B(n44357), .Y(n23063) );
  NOR2X1 U22372 ( .A(n44747), .B(n44348), .Y(n23064) );
  NOR2X1 U22375 ( .A(n44689), .B(n44357), .Y(n23069) );
  NOR2X1 U22379 ( .A(n44751), .B(n44348), .Y(n23070) );
  NOR2X1 U22382 ( .A(n44687), .B(n44357), .Y(n23075) );
  NOR2X1 U22386 ( .A(n44753), .B(n44348), .Y(n23076) );
  NOR2X1 U22389 ( .A(n44685), .B(n44357), .Y(n23081) );
  NOR2X1 U22393 ( .A(n44755), .B(n44348), .Y(n23082) );
  NOR2X1 U22396 ( .A(n44683), .B(n44357), .Y(n23087) );
  NOR2X1 U22400 ( .A(n44749), .B(n44348), .Y(n23088) );
  NOR2X1 U22403 ( .A(n44681), .B(n44357), .Y(n23093) );
  NAND2X1 U22405 ( .A(n73425), .B(n44351), .Y(n22887) );
  NOR2X1 U22408 ( .A(n44745), .B(n44348), .Y(n23094) );
  NOR2X1 U22411 ( .A(n44743), .B(n44374), .Y(n23099) );
  NOR2X1 U22415 ( .A(n44677), .B(n44371), .Y(n23100) );
  NOR2X1 U22418 ( .A(n44679), .B(n44343), .Y(n23105) );
  NOR2X1 U22422 ( .A(n44707), .B(n44334), .Y(n23108) );
  NOR2X1 U22425 ( .A(n44641), .B(n44343), .Y(n23115) );
  NOR2X1 U22429 ( .A(n44705), .B(n44334), .Y(n23116) );
  NOR2X1 U22432 ( .A(n44647), .B(n44343), .Y(n23121) );
  NOR2X1 U22436 ( .A(n44713), .B(n44334), .Y(n23122) );
  NOR2X1 U22439 ( .A(n44649), .B(n44343), .Y(n23127) );
  NOR2X1 U22443 ( .A(n44715), .B(n44334), .Y(n23128) );
  NOR2X1 U22446 ( .A(n44671), .B(n44343), .Y(n23133) );
  NOR2X1 U22450 ( .A(n44737), .B(n44334), .Y(n23134) );
  NOR2X1 U22453 ( .A(n44663), .B(n44343), .Y(n23139) );
  NOR2X1 U22457 ( .A(n44729), .B(n44334), .Y(n23140) );
  NOR2X1 U22460 ( .A(n44673), .B(n44343), .Y(n23145) );
  NOR2X1 U22464 ( .A(n44739), .B(n44334), .Y(n23146) );
  NOR2X1 U22467 ( .A(n44675), .B(n44343), .Y(n23151) );
  NOR2X1 U22471 ( .A(n44741), .B(n44334), .Y(n23152) );
  NOR2X1 U22474 ( .A(n44725), .B(n44374), .Y(n23157) );
  NOR2X1 U22478 ( .A(n44659), .B(n44371), .Y(n23158) );
  NOR2X1 U22481 ( .A(n44655), .B(n44343), .Y(n23163) );
  NOR2X1 U22485 ( .A(n44721), .B(n44334), .Y(n23164) );
  NOR2X1 U22488 ( .A(n44657), .B(n44343), .Y(n23169) );
  NOR2X1 U22492 ( .A(n44723), .B(n44334), .Y(n23170) );
  NOR2X1 U22495 ( .A(n44661), .B(n44343), .Y(n23175) );
  NOR2X1 U22499 ( .A(n44727), .B(n44334), .Y(n23176) );
  NOR2X1 U22502 ( .A(n44653), .B(n44343), .Y(n23181) );
  NOR2X1 U22506 ( .A(n44719), .B(n44334), .Y(n23182) );
  NOR2X1 U22509 ( .A(n44651), .B(n44344), .Y(n23187) );
  NOR2X1 U22513 ( .A(n44717), .B(n44335), .Y(n23188) );
  NOR2X1 U22516 ( .A(n44665), .B(n44344), .Y(n23193) );
  NOR2X1 U22520 ( .A(n44731), .B(n44335), .Y(n23194) );
  NOR2X1 U22523 ( .A(n44677), .B(n44344), .Y(n23199) );
  NOR2X1 U22527 ( .A(n44743), .B(n44335), .Y(n23200) );
  NOR2X1 U22530 ( .A(n44659), .B(n44344), .Y(n23205) );
  NOR2X1 U22534 ( .A(n44725), .B(n44335), .Y(n23206) );
  NOR2X1 U22537 ( .A(n44643), .B(n44344), .Y(n23211) );
  NOR2X1 U22541 ( .A(n44709), .B(n44335), .Y(n23212) );
  NOR2X1 U22544 ( .A(n44645), .B(n44344), .Y(n23217) );
  NOR2X1 U22548 ( .A(n44711), .B(n44335), .Y(n23218) );
  NOR2X1 U22551 ( .A(n44709), .B(n44374), .Y(n23223) );
  NOR2X1 U22555 ( .A(n44643), .B(n44371), .Y(n23224) );
  NOR2X1 U22558 ( .A(n44669), .B(n44344), .Y(n23229) );
  NOR2X1 U22562 ( .A(n44735), .B(n44335), .Y(n23230) );
  NOR2X1 U22565 ( .A(n44667), .B(n44344), .Y(n23235) );
  NOR2X1 U22569 ( .A(n44733), .B(n44335), .Y(n23236) );
  NOR2X1 U22572 ( .A(n44693), .B(n44344), .Y(n23241) );
  NOR2X1 U22576 ( .A(n44757), .B(n44335), .Y(n23242) );
  NOR2X1 U22579 ( .A(n44697), .B(n44344), .Y(n23247) );
  NOR2X1 U22583 ( .A(n44761), .B(n44335), .Y(n23248) );
  NOR2X1 U22586 ( .A(n44699), .B(n44344), .Y(n23253) );
  NOR2X1 U22590 ( .A(n44763), .B(n44335), .Y(n23254) );
  NOR2X1 U22593 ( .A(n44703), .B(n44344), .Y(n23259) );
  NOR2X1 U22597 ( .A(n44767), .B(n44335), .Y(n23260) );
  NOR2X1 U22600 ( .A(n44701), .B(n44345), .Y(n23265) );
  NOR2X1 U22604 ( .A(n44765), .B(n44336), .Y(n23266) );
  NOR2X1 U22607 ( .A(n44695), .B(n44345), .Y(n23271) );
  NOR2X1 U22611 ( .A(n44759), .B(n44336), .Y(n23272) );
  NOR2X1 U22614 ( .A(n44691), .B(n44345), .Y(n23277) );
  NOR2X1 U22618 ( .A(n44747), .B(n44336), .Y(n23278) );
  NOR2X1 U22621 ( .A(n44689), .B(n44345), .Y(n23283) );
  NOR2X1 U22625 ( .A(n44751), .B(n44336), .Y(n23284) );
  NOR2X1 U22628 ( .A(n44711), .B(n44374), .Y(n23289) );
  NOR2X1 U22632 ( .A(n44645), .B(n44371), .Y(n23290) );
  NOR2X1 U22635 ( .A(n44687), .B(n44345), .Y(n23295) );
  NOR2X1 U22639 ( .A(n44753), .B(n44336), .Y(n23296) );
  NOR2X1 U22642 ( .A(n44685), .B(n44345), .Y(n23301) );
  NOR2X1 U22646 ( .A(n44755), .B(n44336), .Y(n23302) );
  NOR2X1 U22649 ( .A(n44683), .B(n44345), .Y(n23307) );
  NOR2X1 U22653 ( .A(n44749), .B(n44336), .Y(n23308) );
  NOR2X1 U22656 ( .A(n44681), .B(n44345), .Y(n23313) );
  NAND2X1 U22658 ( .A(n549), .B(n44339), .Y(n23107) );
  NOR2X1 U22661 ( .A(n44745), .B(n44336), .Y(n23314) );
  NOR2X1 U22664 ( .A(n44679), .B(n44331), .Y(n23319) );
  NOR2X1 U22668 ( .A(n44707), .B(n44322), .Y(n23322) );
  NOR2X1 U22671 ( .A(n44735), .B(n44374), .Y(n23329) );
  NOR2X1 U22675 ( .A(n44669), .B(n44371), .Y(n23330) );
  NOR2X1 U22678 ( .A(n44641), .B(n44331), .Y(n23335) );
  NOR2X1 U22682 ( .A(n44705), .B(n44322), .Y(n23336) );
  NOR2X1 U22685 ( .A(n44647), .B(n44331), .Y(n23341) );
  NOR2X1 U22689 ( .A(n44713), .B(n44322), .Y(n23342) );
  NOR2X1 U22692 ( .A(n44649), .B(n44331), .Y(n23347) );
  NOR2X1 U22696 ( .A(n44715), .B(n44322), .Y(n23348) );
  NOR2X1 U22699 ( .A(n44671), .B(n44331), .Y(n23353) );
  NOR2X1 U22703 ( .A(n44737), .B(n44322), .Y(n23354) );
  NOR2X1 U22706 ( .A(n44663), .B(n44331), .Y(n23359) );
  NOR2X1 U22710 ( .A(n44729), .B(n44322), .Y(n23360) );
  NOR2X1 U22713 ( .A(n44673), .B(n44331), .Y(n23365) );
  NOR2X1 U22717 ( .A(n44739), .B(n44322), .Y(n23366) );
  NOR2X1 U22720 ( .A(n44675), .B(n44331), .Y(n23371) );
  NOR2X1 U22724 ( .A(n44741), .B(n44322), .Y(n23372) );
  NOR2X1 U22727 ( .A(n44655), .B(n44331), .Y(n23377) );
  NOR2X1 U22731 ( .A(n44721), .B(n44322), .Y(n23378) );
  NOR2X1 U22734 ( .A(n44657), .B(n44331), .Y(n23383) );
  NOR2X1 U22738 ( .A(n44723), .B(n44322), .Y(n23384) );
  NOR2X1 U22741 ( .A(n44661), .B(n44331), .Y(n23389) );
  NOR2X1 U22745 ( .A(n44727), .B(n44322), .Y(n23390) );
  NOR2X1 U22748 ( .A(n44733), .B(n44374), .Y(n23395) );
  NOR2X1 U22752 ( .A(n44667), .B(n44371), .Y(n23396) );
  NOR2X1 U22755 ( .A(n44653), .B(n44331), .Y(n23401) );
  NOR2X1 U22759 ( .A(n44719), .B(n44322), .Y(n23402) );
  NOR2X1 U22762 ( .A(n44651), .B(n44332), .Y(n23407) );
  NOR2X1 U22766 ( .A(n44717), .B(n44323), .Y(n23408) );
  NOR2X1 U22769 ( .A(n44665), .B(n44332), .Y(n23413) );
  NOR2X1 U22773 ( .A(n44731), .B(n44323), .Y(n23414) );
  NOR2X1 U22776 ( .A(n44677), .B(n44332), .Y(n23419) );
  NOR2X1 U22780 ( .A(n44743), .B(n44323), .Y(n23420) );
  NOR2X1 U22783 ( .A(n44659), .B(n44332), .Y(n23425) );
  NOR2X1 U22787 ( .A(n44725), .B(n44323), .Y(n23426) );
  NOR2X1 U22790 ( .A(n44643), .B(n44332), .Y(n23431) );
  NOR2X1 U22794 ( .A(n44709), .B(n44323), .Y(n23432) );
  NOR2X1 U22797 ( .A(n44645), .B(n44332), .Y(n23437) );
  NOR2X1 U22801 ( .A(n44711), .B(n44323), .Y(n23438) );
  NOR2X1 U22804 ( .A(n44669), .B(n44332), .Y(n23443) );
  NOR2X1 U22808 ( .A(n44735), .B(n44323), .Y(n23444) );
  NOR2X1 U22811 ( .A(n44667), .B(n44332), .Y(n23449) );
  NOR2X1 U22815 ( .A(n44733), .B(n44323), .Y(n23450) );
  NOR2X1 U22818 ( .A(n44693), .B(n44332), .Y(n23455) );
  NOR2X1 U22822 ( .A(n44757), .B(n44323), .Y(n23456) );
  NOR2X1 U22825 ( .A(n44757), .B(n44374), .Y(n23461) );
  NOR2X1 U22829 ( .A(n44693), .B(n44371), .Y(n23462) );
  NOR2X1 U22832 ( .A(n44697), .B(n44332), .Y(n23467) );
  NOR2X1 U22836 ( .A(n44761), .B(n44323), .Y(n23468) );
  NOR2X1 U22839 ( .A(n44699), .B(n44332), .Y(n23473) );
  NOR2X1 U22843 ( .A(n44763), .B(n44323), .Y(n23474) );
  NOR2X1 U22846 ( .A(n44703), .B(n44332), .Y(n23479) );
  NOR2X1 U22850 ( .A(n44767), .B(n44323), .Y(n23480) );
  NOR2X1 U22853 ( .A(n44701), .B(n44333), .Y(n23485) );
  NOR2X1 U22857 ( .A(n44765), .B(n44324), .Y(n23486) );
  NOR2X1 U22860 ( .A(n44695), .B(n44333), .Y(n23491) );
  NOR2X1 U22864 ( .A(n44759), .B(n44324), .Y(n23492) );
  NOR2X1 U22867 ( .A(n44691), .B(n44333), .Y(n23497) );
  NOR2X1 U22871 ( .A(n44747), .B(n44324), .Y(n23498) );
  NOR2X1 U22874 ( .A(n44689), .B(n44333), .Y(n23503) );
  NOR2X1 U22878 ( .A(n44751), .B(n44324), .Y(n23504) );
  NOR2X1 U22881 ( .A(n44687), .B(n44333), .Y(n23509) );
  NOR2X1 U22885 ( .A(n44753), .B(n44324), .Y(n23510) );
  NOR2X1 U22888 ( .A(n44685), .B(n44333), .Y(n23515) );
  NOR2X1 U22892 ( .A(n44755), .B(n44324), .Y(n23516) );
  NOR2X1 U22895 ( .A(n44683), .B(n44333), .Y(n23521) );
  NOR2X1 U22899 ( .A(n44749), .B(n44324), .Y(n23522) );
  NOR2X1 U22902 ( .A(n44761), .B(n44374), .Y(n23527) );
  NOR2X1 U22906 ( .A(n44697), .B(n44371), .Y(n23528) );
  NOR2X1 U22909 ( .A(n44681), .B(n44333), .Y(n23533) );
  NAND2X1 U22911 ( .A(n547), .B(n44327), .Y(n23321) );
  NOR2X1 U22914 ( .A(n44745), .B(n44324), .Y(n23534) );
  NOR2X1 U22917 ( .A(n44679), .B(n44319), .Y(n23539) );
  NOR2X1 U22921 ( .A(n44707), .B(n44310), .Y(n23542) );
  NOR2X1 U22924 ( .A(n44641), .B(n44319), .Y(n23549) );
  NOR2X1 U22928 ( .A(n44705), .B(n44310), .Y(n23550) );
  NOR2X1 U22931 ( .A(n44647), .B(n44319), .Y(n23555) );
  NOR2X1 U22935 ( .A(n44713), .B(n44310), .Y(n23556) );
  NOR2X1 U22938 ( .A(n44649), .B(n44319), .Y(n23561) );
  NOR2X1 U22942 ( .A(n44715), .B(n44310), .Y(n23562) );
  NOR2X1 U22945 ( .A(n44763), .B(n44374), .Y(n23567) );
  NOR2X1 U22949 ( .A(n44699), .B(n44371), .Y(n23568) );
  NOR2X1 U22952 ( .A(n44671), .B(n44319), .Y(n23573) );
  NOR2X1 U22956 ( .A(n44737), .B(n44310), .Y(n23574) );
  NOR2X1 U22959 ( .A(n44663), .B(n44319), .Y(n23579) );
  NOR2X1 U22963 ( .A(n44729), .B(n44310), .Y(n23580) );
  NOR2X1 U22966 ( .A(n44673), .B(n44319), .Y(n23585) );
  NOR2X1 U22970 ( .A(n44739), .B(n44310), .Y(n23586) );
  NOR2X1 U22973 ( .A(n44675), .B(n44319), .Y(n23591) );
  NOR2X1 U22977 ( .A(n44741), .B(n44310), .Y(n23592) );
  NOR2X1 U22980 ( .A(n44655), .B(n44319), .Y(n23597) );
  NOR2X1 U22984 ( .A(n44721), .B(n44310), .Y(n23598) );
  NOR2X1 U22987 ( .A(n44657), .B(n44319), .Y(n23603) );
  NOR2X1 U22991 ( .A(n44723), .B(n44310), .Y(n23604) );
  NOR2X1 U22994 ( .A(n44661), .B(n44319), .Y(n23609) );
  NOR2X1 U22998 ( .A(n44727), .B(n44310), .Y(n23610) );
  NOR2X1 U23001 ( .A(n44653), .B(n44319), .Y(n23615) );
  NOR2X1 U23005 ( .A(n44719), .B(n44310), .Y(n23616) );
  NOR2X1 U23008 ( .A(n44651), .B(n44320), .Y(n23621) );
  NOR2X1 U23012 ( .A(n44717), .B(n44311), .Y(n23622) );
  NOR2X1 U23015 ( .A(n44665), .B(n44320), .Y(n23627) );
  NOR2X1 U23019 ( .A(n44731), .B(n44311), .Y(n23628) );
  NOR2X1 U23022 ( .A(n44767), .B(n44374), .Y(n23633) );
  NOR2X1 U23026 ( .A(n44703), .B(n44371), .Y(n23634) );
  NOR2X1 U23029 ( .A(n44677), .B(n44320), .Y(n23639) );
  NOR2X1 U23033 ( .A(n44743), .B(n44311), .Y(n23640) );
  NOR2X1 U23036 ( .A(n44659), .B(n44320), .Y(n23645) );
  NOR2X1 U23040 ( .A(n44725), .B(n44311), .Y(n23646) );
  NOR2X1 U23043 ( .A(n44643), .B(n44320), .Y(n23651) );
  NOR2X1 U23047 ( .A(n44709), .B(n44311), .Y(n23652) );
  NOR2X1 U23050 ( .A(n44645), .B(n44320), .Y(n23657) );
  NOR2X1 U23054 ( .A(n44711), .B(n44311), .Y(n23658) );
  NOR2X1 U23057 ( .A(n44669), .B(n44320), .Y(n23663) );
  NOR2X1 U23061 ( .A(n44735), .B(n44311), .Y(n23664) );
  NOR2X1 U23064 ( .A(n44667), .B(n44320), .Y(n23669) );
  NOR2X1 U23068 ( .A(n44733), .B(n44311), .Y(n23670) );
  NOR2X1 U23071 ( .A(n44693), .B(n44320), .Y(n23675) );
  NOR2X1 U23075 ( .A(n44757), .B(n44311), .Y(n23676) );
  NOR2X1 U23078 ( .A(n44697), .B(n44320), .Y(n23681) );
  NOR2X1 U23082 ( .A(n44761), .B(n44311), .Y(n23682) );
  NOR2X1 U23085 ( .A(n44699), .B(n44320), .Y(n23687) );
  NOR2X1 U23089 ( .A(n44763), .B(n44311), .Y(n23688) );
  NOR2X1 U23092 ( .A(n44703), .B(n44320), .Y(n23693) );
  NOR2X1 U23096 ( .A(n44767), .B(n44311), .Y(n23694) );
  NOR2X1 U23099 ( .A(n44765), .B(n44375), .Y(n23699) );
  NOR2X1 U23103 ( .A(n44701), .B(n44372), .Y(n23700) );
  NOR2X1 U23106 ( .A(n44701), .B(n44321), .Y(n23705) );
  NOR2X1 U23110 ( .A(n44765), .B(n44312), .Y(n23706) );
  NOR2X1 U23113 ( .A(n44695), .B(n44321), .Y(n23711) );
  NOR2X1 U23117 ( .A(n44759), .B(n44312), .Y(n23712) );
  NOR2X1 U23120 ( .A(n44691), .B(n44321), .Y(n23717) );
  NOR2X1 U23124 ( .A(n44747), .B(n44312), .Y(n23718) );
  NOR2X1 U23127 ( .A(n44689), .B(n44321), .Y(n23723) );
  NOR2X1 U23131 ( .A(n44751), .B(n44312), .Y(n23724) );
  NOR2X1 U23134 ( .A(n44687), .B(n44321), .Y(n23729) );
  NOR2X1 U23138 ( .A(n44753), .B(n44312), .Y(n23730) );
  NOR2X1 U23141 ( .A(n44685), .B(n44321), .Y(n23735) );
  NOR2X1 U23145 ( .A(n44755), .B(n44312), .Y(n23736) );
  NOR2X1 U23148 ( .A(n44683), .B(n44321), .Y(n23741) );
  NOR2X1 U23152 ( .A(n44749), .B(n44312), .Y(n23742) );
  NOR2X1 U23155 ( .A(n44681), .B(n44321), .Y(n23747) );
  NAND2X1 U23157 ( .A(n552), .B(n44315), .Y(n23541) );
  NOR2X1 U23160 ( .A(n44745), .B(n44312), .Y(n23748) );
  NOR2X1 U23163 ( .A(n44759), .B(n44375), .Y(n23753) );
  NOR2X1 U23167 ( .A(n44695), .B(n44372), .Y(n23754) );
  NOR2X1 U23170 ( .A(n44679), .B(n44307), .Y(n23759) );
  NOR2X1 U23174 ( .A(n44707), .B(n44298), .Y(n23762) );
  NOR2X1 U23177 ( .A(n44641), .B(n44307), .Y(n23769) );
  NOR2X1 U23181 ( .A(n44705), .B(n44298), .Y(n23770) );
  NOR2X1 U23184 ( .A(n44647), .B(n44307), .Y(n23775) );
  NOR2X1 U23188 ( .A(n44713), .B(n44298), .Y(n23776) );
  NOR2X1 U23191 ( .A(n44649), .B(n44307), .Y(n23781) );
  NOR2X1 U23195 ( .A(n44715), .B(n44298), .Y(n23782) );
  NOR2X1 U23198 ( .A(n44671), .B(n44307), .Y(n23787) );
  NOR2X1 U23202 ( .A(n44737), .B(n44298), .Y(n23788) );
  NOR2X1 U23205 ( .A(n44663), .B(n44307), .Y(n23793) );
  NOR2X1 U23209 ( .A(n44729), .B(n44298), .Y(n23794) );
  NOR2X1 U23212 ( .A(n44673), .B(n44307), .Y(n23799) );
  NOR2X1 U23216 ( .A(n44739), .B(n44298), .Y(n23800) );
  NOR2X1 U23219 ( .A(n44747), .B(n44375), .Y(n23805) );
  NOR2X1 U23223 ( .A(n44691), .B(n44372), .Y(n23806) );
  NOR2X1 U23226 ( .A(n44675), .B(n44307), .Y(n23811) );
  NOR2X1 U23230 ( .A(n44741), .B(n44298), .Y(n23812) );
  NOR2X1 U23233 ( .A(n44655), .B(n44307), .Y(n23817) );
  NOR2X1 U23237 ( .A(n44721), .B(n44298), .Y(n23818) );
  NOR2X1 U23240 ( .A(n44657), .B(n44307), .Y(n23823) );
  NOR2X1 U23244 ( .A(n44723), .B(n44298), .Y(n23824) );
  NOR2X1 U23247 ( .A(n44661), .B(n44307), .Y(n23829) );
  NOR2X1 U23251 ( .A(n44727), .B(n44298), .Y(n23830) );
  NOR2X1 U23254 ( .A(n44653), .B(n44307), .Y(n23835) );
  NOR2X1 U23258 ( .A(n44719), .B(n44298), .Y(n23836) );
  NOR2X1 U23261 ( .A(n44651), .B(n44308), .Y(n23841) );
  NOR2X1 U23265 ( .A(n44717), .B(n44299), .Y(n23842) );
  NOR2X1 U23268 ( .A(n44665), .B(n44308), .Y(n23847) );
  NOR2X1 U23272 ( .A(n44731), .B(n44299), .Y(n23848) );
  NOR2X1 U23275 ( .A(n44677), .B(n44308), .Y(n23853) );
  NOR2X1 U23279 ( .A(n44743), .B(n44299), .Y(n23854) );
  NOR2X1 U23282 ( .A(n44659), .B(n44308), .Y(n23859) );
  NOR2X1 U23286 ( .A(n44725), .B(n44299), .Y(n23860) );
  NOR2X1 U23289 ( .A(n44643), .B(n44308), .Y(n23865) );
  NOR2X1 U23293 ( .A(n44709), .B(n44299), .Y(n23866) );
  NOR2X1 U23296 ( .A(n44751), .B(n44375), .Y(n23871) );
  NOR2X1 U23300 ( .A(n44689), .B(n44372), .Y(n23872) );
  NOR2X1 U23303 ( .A(n44645), .B(n44308), .Y(n23877) );
  NOR2X1 U23307 ( .A(n44711), .B(n44299), .Y(n23878) );
  NOR2X1 U23310 ( .A(n44669), .B(n44308), .Y(n23883) );
  NOR2X1 U23314 ( .A(n44735), .B(n44299), .Y(n23884) );
  NOR2X1 U23317 ( .A(n44667), .B(n44308), .Y(n23889) );
  NOR2X1 U23321 ( .A(n44733), .B(n44299), .Y(n23890) );
  NOR2X1 U23324 ( .A(n44693), .B(n44308), .Y(n23895) );
  NOR2X1 U23328 ( .A(n44757), .B(n44299), .Y(n23896) );
  NOR2X1 U23331 ( .A(n44697), .B(n44308), .Y(n23901) );
  NOR2X1 U23335 ( .A(n44761), .B(n44299), .Y(n23902) );
  NOR2X1 U23338 ( .A(n44699), .B(n44308), .Y(n23907) );
  NOR2X1 U23342 ( .A(n44763), .B(n44299), .Y(n23908) );
  NOR2X1 U23345 ( .A(n44703), .B(n44308), .Y(n23913) );
  NOR2X1 U23349 ( .A(n44767), .B(n44299), .Y(n23914) );
  NOR2X1 U23352 ( .A(n44701), .B(n44309), .Y(n23919) );
  NOR2X1 U23356 ( .A(n44765), .B(n44300), .Y(n23920) );
  NOR2X1 U23359 ( .A(n44695), .B(n44309), .Y(n23925) );
  NOR2X1 U23363 ( .A(n44759), .B(n44300), .Y(n23926) );
  NOR2X1 U23366 ( .A(n44691), .B(n44309), .Y(n23931) );
  NOR2X1 U23370 ( .A(n44747), .B(n44300), .Y(n23932) );
  NOR2X1 U23373 ( .A(n44753), .B(n44375), .Y(n23937) );
  NOR2X1 U23377 ( .A(n44687), .B(n44372), .Y(n23938) );
  NOR2X1 U23380 ( .A(n44689), .B(n44309), .Y(n23943) );
  NOR2X1 U23384 ( .A(n44751), .B(n44300), .Y(n23944) );
  NOR2X1 U23387 ( .A(n44687), .B(n44309), .Y(n23949) );
  NOR2X1 U23391 ( .A(n44753), .B(n44300), .Y(n23950) );
  NOR2X1 U23394 ( .A(n44685), .B(n44309), .Y(n23955) );
  NOR2X1 U23398 ( .A(n44755), .B(n44300), .Y(n23956) );
  NOR2X1 U23401 ( .A(n44683), .B(n44309), .Y(n23961) );
  NOR2X1 U23405 ( .A(n44749), .B(n44300), .Y(n23962) );
  NOR2X1 U23408 ( .A(n44681), .B(n44309), .Y(n23967) );
  NAND2X1 U23410 ( .A(n543), .B(n44303), .Y(n23761) );
  NOR2X1 U23413 ( .A(n44745), .B(n44300), .Y(n23968) );
  NOR2X1 U23416 ( .A(n44755), .B(n44375), .Y(n23973) );
  NOR2X1 U23420 ( .A(n44685), .B(n44372), .Y(n23974) );
  NOR2X1 U23423 ( .A(n44804), .B(n37657), .Y(n23979) );
  NOR2X1 U23427 ( .A(n44807), .B(n37628), .Y(n23980) );
  NOR2X1 U23430 ( .A(n44804), .B(n37656), .Y(n23985) );
  NOR2X1 U23434 ( .A(n44807), .B(n37627), .Y(n23986) );
  NOR2X1 U23437 ( .A(n44804), .B(n37655), .Y(n23991) );
  NOR2X1 U23441 ( .A(n44807), .B(n37626), .Y(n23992) );
  NOR2X1 U23444 ( .A(n44804), .B(n37654), .Y(n23997) );
  NOR2X1 U23448 ( .A(n44807), .B(n37625), .Y(n23998) );
  NOR2X1 U23451 ( .A(n44804), .B(n37653), .Y(n24003) );
  NOR2X1 U23455 ( .A(n44807), .B(n37624), .Y(n24004) );
  NOR2X1 U23458 ( .A(n44804), .B(n37652), .Y(n24009) );
  NOR2X1 U23462 ( .A(n44807), .B(n37623), .Y(n24010) );
  NOR2X1 U23465 ( .A(n44804), .B(n37651), .Y(n24015) );
  NOR2X1 U23469 ( .A(n44807), .B(n37622), .Y(n24016) );
  NOR2X1 U23472 ( .A(n44804), .B(n37650), .Y(n24021) );
  NOR2X1 U23476 ( .A(n44807), .B(n37621), .Y(n24022) );
  NOR2X1 U23479 ( .A(n44804), .B(n37649), .Y(n24027) );
  NOR2X1 U23483 ( .A(n44807), .B(n37620), .Y(n24028) );
  NOR2X1 U23486 ( .A(n44804), .B(n37648), .Y(n24033) );
  NOR2X1 U23490 ( .A(n44807), .B(n37619), .Y(n24034) );
  NOR2X1 U23493 ( .A(n44749), .B(n44375), .Y(n24039) );
  NOR2X1 U23497 ( .A(n44683), .B(n44372), .Y(n24040) );
  NOR2X1 U23500 ( .A(n44804), .B(n37647), .Y(n24045) );
  NOR2X1 U23504 ( .A(n44807), .B(n37618), .Y(n24046) );
  NOR2X1 U23507 ( .A(n44804), .B(n37602), .Y(n24051) );
  NOR2X1 U23511 ( .A(n44807), .B(n37599), .Y(n24052) );
  NOR2X1 U23514 ( .A(n44805), .B(n37646), .Y(n24057) );
  NOR2X1 U23518 ( .A(n44808), .B(n37617), .Y(n24058) );
  NOR2X1 U23521 ( .A(n44805), .B(n37645), .Y(n24063) );
  NOR2X1 U23525 ( .A(n44808), .B(n37616), .Y(n24064) );
  NOR2X1 U23528 ( .A(n44805), .B(n37644), .Y(n24069) );
  NOR2X1 U23532 ( .A(n44808), .B(n37615), .Y(n24070) );
  NOR2X1 U23535 ( .A(n44805), .B(n37643), .Y(n24075) );
  NOR2X1 U23539 ( .A(n44808), .B(n37614), .Y(n24076) );
  NOR2X1 U23542 ( .A(n44805), .B(n37642), .Y(n24081) );
  NOR2X1 U23546 ( .A(n44808), .B(n37613), .Y(n24082) );
  NOR2X1 U23549 ( .A(n44805), .B(n37641), .Y(n24087) );
  NOR2X1 U23553 ( .A(n44808), .B(n37612), .Y(n24088) );
  NOR2X1 U23556 ( .A(n44805), .B(n37640), .Y(n24093) );
  NOR2X1 U23560 ( .A(n44808), .B(n37611), .Y(n24094) );
  NOR2X1 U23563 ( .A(n44805), .B(n37639), .Y(n24099) );
  NAND2X1 U23565 ( .A(n518), .B(n44606), .Y(n18002) );
  NOR2X1 U23568 ( .A(n44808), .B(n37610), .Y(n24102) );
  NOR2X1 U23571 ( .A(n44745), .B(n44375), .Y(n24108) );
  NOR2X1 U23576 ( .A(n44681), .B(n44372), .Y(n24110) );
  NOR2X1 U23577 ( .A(n24112), .B(n24113), .Y(u_decode_scoreboard_r[9]) );
  NAND2X1 U23578 ( .A(n24114), .B(n24115), .Y(n24113) );
  NAND2X1 U23579 ( .A(n73423), .B(n1054), .Y(n24114) );
  NOR2X1 U23582 ( .A(n24119), .B(n24120), .Y(u_decode_scoreboard_r[8]) );
  NAND2X1 U23583 ( .A(n24121), .B(n24122), .Y(n24120) );
  NAND2X1 U23584 ( .A(n24123), .B(n73423), .Y(n24121) );
  NAND2X1 U23612 ( .A(n24165), .B(n24166), .Y(n24164) );
  NAND2X1 U23613 ( .A(n24167), .B(n73422), .Y(n24165) );
  NAND2X1 U23630 ( .A(n24191), .B(n24192), .Y(n24190) );
  NAND2X1 U23631 ( .A(n24193), .B(n73422), .Y(n24191) );
  NAND2X1 U23648 ( .A(n24213), .B(n24214), .Y(n24212) );
  NAND2X1 U23649 ( .A(n73424), .B(n24167), .Y(n24213) );
  NAND2X1 U23654 ( .A(n24220), .B(n24221), .Y(n24219) );
  NAND2X1 U23655 ( .A(n24193), .B(n73424), .Y(n24220) );
  NOR2X1 U23659 ( .A(n24225), .B(n24226), .Y(u_decode_scoreboard_r[25]) );
  NAND2X1 U23660 ( .A(n24227), .B(n24228), .Y(n24226) );
  NOR2X1 U23663 ( .A(n24231), .B(n24180), .Y(n24225) );
  NOR2X1 U23664 ( .A(n24232), .B(n24233), .Y(u_decode_scoreboard_r[24]) );
  NAND2X1 U23665 ( .A(n24234), .B(n24235), .Y(n24233) );
  NAND2X1 U23666 ( .A(n73424), .B(n24123), .Y(n24234) );
  NOR2X1 U23695 ( .A(n24271), .B(n24272), .Y(u_decode_scoreboard_r[1]) );
  NAND2X1 U23696 ( .A(n24273), .B(n24274), .Y(n24272) );
  NOR2X1 U23699 ( .A(n24231), .B(n24135), .Y(n24271) );
  NAND2X1 U23702 ( .A(n24279), .B(n24280), .Y(n24278) );
  NAND2X1 U23703 ( .A(n73426), .B(n24167), .Y(n24279) );
  NAND2X1 U23708 ( .A(n24286), .B(n24287), .Y(n24285) );
  NAND2X1 U23709 ( .A(n73426), .B(n24193), .Y(n24286) );
  NOR2X1 U23713 ( .A(n24291), .B(n24292), .Y(u_decode_scoreboard_r[17]) );
  NAND2X1 U23714 ( .A(n24293), .B(n24294), .Y(n24292) );
  NAND2X1 U23715 ( .A(n73426), .B(n1054), .Y(n24293) );
  NAND2X1 U23716 ( .A(n24295), .B(n24296), .Y(n24231) );
  NOR2X1 U23717 ( .A(u_csr_writeback_idx_q[2]), .B(u_csr_writeback_idx_q[1]), 
        .Y(n24296) );
  NOR2X1 U23721 ( .A(n24299), .B(n24300), .Y(u_decode_scoreboard_r[16]) );
  NAND2X1 U23722 ( .A(n24301), .B(n24302), .Y(n24300) );
  NAND2X1 U23723 ( .A(n73426), .B(n24123), .Y(n24301) );
  AND2X1 U23724 ( .A(n36767), .B(n37483), .Y(n24123) );
  NAND2X1 U23737 ( .A(n37597), .B(n24319), .Y(n24136) );
  NAND2X1 U23746 ( .A(n24319), .B(n37337), .Y(n24145) );
  NAND2X1 U23753 ( .A(n24337), .B(n24319), .Y(n24154) );
  NAND2X1 U23763 ( .A(n24319), .B(n36767), .Y(n24162) );
  NOR2X1 U23764 ( .A(n37483), .B(n24237), .Y(n24319) );
  NAND2X1 U23766 ( .A(n24348), .B(n24349), .Y(n24347) );
  NAND2X1 U23767 ( .A(n24167), .B(n73423), .Y(n24348) );
  AND2X1 U23768 ( .A(n37597), .B(n24350), .Y(n24167) );
  NAND2X1 U23774 ( .A(n24356), .B(n24357), .Y(n24355) );
  NAND2X1 U23775 ( .A(n24193), .B(n73423), .Y(n24356) );
  AND2X1 U23778 ( .A(n24350), .B(n37337), .Y(n24193) );
  NOR2X1 U23779 ( .A(u_csr_writeback_idx_q[2]), .B(n24237), .Y(n24350) );
  NAND2X1 U23788 ( .A(n24366), .B(n44082), .Y(n24365) );
  NOR2X1 U23789 ( .A(n15219), .B(n24367), .Y(n24366) );
  NOR2X1 U23795 ( .A(n73535), .B(n24378), .Y(n24376) );
  NOR2X1 U23798 ( .A(n24382), .B(n24383), .Y(n24379) );
  NOR2X1 U23799 ( .A(n24384), .B(n24385), .Y(n24383) );
  NOR2X1 U23800 ( .A(n73537), .B(n24386), .Y(n24382) );
  NOR2X1 U23801 ( .A(n24387), .B(n73528), .Y(n24386) );
  NOR2X1 U23802 ( .A(n24388), .B(n24389), .Y(n24387) );
  AND2X1 U23813 ( .A(n24405), .B(n24406), .Y(n24403) );
  AND2X1 U23815 ( .A(n24409), .B(n24410), .Y(n24407) );
  NAND2X1 U23817 ( .A(n24413), .B(n24414), .Y(n24412) );
  NAND2X1 U23818 ( .A(n73531), .B(n24415), .Y(n24414) );
  NAND2X1 U23819 ( .A(n24397), .B(n24416), .Y(n24415) );
  NOR2X1 U23820 ( .A(n73534), .B(n73533), .Y(n24397) );
  NOR2X1 U23821 ( .A(n24419), .B(n24420), .Y(n24413) );
  NOR2X1 U23822 ( .A(n24421), .B(n24422), .Y(n24420) );
  NOR2X1 U23823 ( .A(n37572), .B(n24381), .Y(n24421) );
  OR2X1 U23824 ( .A(n73535), .B(n37570), .Y(n24381) );
  NOR2X1 U23825 ( .A(n24425), .B(n24426), .Y(n24419) );
  NAND2X1 U23826 ( .A(n73398), .B(n73537), .Y(n24426) );
  NAND2X1 U23827 ( .A(n73536), .B(n24429), .Y(n24425) );
  NAND2X1 U23828 ( .A(n24430), .B(n24431), .Y(n24411) );
  NAND2X1 U23829 ( .A(n24432), .B(n24433), .Y(n24431) );
  NOR2X1 U23830 ( .A(n73541), .B(n24434), .Y(n24433) );
  NAND2X1 U23831 ( .A(n24435), .B(n24436), .Y(n24434) );
  NOR2X1 U23832 ( .A(n24437), .B(n24438), .Y(n24432) );
  NAND2X1 U23833 ( .A(n596), .B(n73529), .Y(n24438) );
  NOR2X1 U23834 ( .A(n73515), .B(n24441), .Y(n24430) );
  NOR2X1 U23835 ( .A(n24442), .B(n24443), .Y(n24441) );
  NAND2X1 U23836 ( .A(n24444), .B(n73530), .Y(n24443) );
  NOR2X1 U23837 ( .A(n24445), .B(n24446), .Y(n24444) );
  NAND2X1 U23838 ( .A(n24447), .B(n24448), .Y(n24442) );
  NOR2X1 U23839 ( .A(n602), .B(n24449), .Y(n24447) );
  NOR2X1 U23840 ( .A(n24450), .B(n24451), .Y(n24449) );
  NOR2X1 U23841 ( .A(n24452), .B(n24453), .Y(n24451) );
  NAND2X1 U23842 ( .A(n621), .B(n24454), .Y(n24453) );
  NAND2X1 U23843 ( .A(n73533), .B(n24455), .Y(n24452) );
  NOR2X1 U23844 ( .A(n24456), .B(n24457), .Y(n24450) );
  NAND2X1 U23845 ( .A(n73541), .B(n24458), .Y(n24457) );
  NAND2X1 U23846 ( .A(n24459), .B(n24460), .Y(n24456) );
  NOR2X1 U23847 ( .A(n24461), .B(n24455), .Y(n24459) );
  NOR2X1 U23848 ( .A(n24462), .B(n24463), .Y(n24461) );
  NOR2X1 U23849 ( .A(n73558), .B(n24435), .Y(n24463) );
  NOR2X1 U23888 ( .A(n73558), .B(n24504), .Y(n24502) );
  NAND2X1 U23898 ( .A(n24464), .B(n24473), .Y(n24511) );
  NOR2X1 U23899 ( .A(n24446), .B(n24512), .Y(n24508) );
  NAND2X1 U23900 ( .A(n24458), .B(n24460), .Y(n24512) );
  AND2X1 U23901 ( .A(n24513), .B(n24514), .Y(n24460) );
  NOR2X1 U23902 ( .A(n24515), .B(n24516), .Y(n24514) );
  NAND2X1 U23903 ( .A(n24517), .B(n24518), .Y(n24516) );
  NOR2X1 U23904 ( .A(n24519), .B(n24520), .Y(n24513) );
  NAND2X1 U23905 ( .A(n37561), .B(n24522), .Y(n24520) );
  AND2X1 U23906 ( .A(n24523), .B(n24454), .Y(n24458) );
  NOR2X1 U23907 ( .A(n24524), .B(n24525), .Y(n24523) );
  NAND2X1 U23908 ( .A(n24526), .B(n24527), .Y(n24446) );
  NOR2X1 U23909 ( .A(n24384), .B(n24528), .Y(n24527) );
  NOR2X1 U23910 ( .A(n24529), .B(n24530), .Y(n24526) );
  NOR2X1 U23940 ( .A(n24539), .B(n24535), .Y(n24538) );
  NOR2X1 U23970 ( .A(n24555), .B(n24556), .Y(n24448) );
  OR2X1 U23971 ( .A(n24557), .B(n24469), .Y(n24555) );
  NOR2X1 U23985 ( .A(n24564), .B(n24474), .Y(n24488) );
  NAND2X1 U23986 ( .A(n24552), .B(n24565), .Y(n24474) );
  NOR2X1 U23987 ( .A(n606), .B(n24566), .Y(n24565) );
  OR2X1 U23988 ( .A(n24556), .B(n24557), .Y(n24566) );
  NOR2X1 U23989 ( .A(n24445), .B(n24436), .Y(n24552) );
  OR2X1 U23990 ( .A(n24469), .B(n24473), .Y(n24564) );
  NAND2X1 U24012 ( .A(n24570), .B(n24571), .Y(n24533) );
  NOR2X1 U24013 ( .A(n24572), .B(n612), .Y(n24571) );
  NOR2X1 U24014 ( .A(n24574), .B(n24429), .Y(n24570) );
  NOR2X1 U24282 ( .A(n37562), .B(n24842), .Y(n24839) );
  AND2X1 U24283 ( .A(n44085), .B(mem_i_inst_i[4]), .Y(n24842) );
  NOR2X1 U24291 ( .A(n37562), .B(n24847), .Y(n24845) );
  AND2X1 U24292 ( .A(n44086), .B(mem_i_inst_i[6]), .Y(n24847) );
  NAND2X1 U24293 ( .A(n24848), .B(n24573), .Y(n24539) );
  NAND2X1 U24294 ( .A(n24849), .B(n24850), .Y(n24573) );
  NOR2X1 U24296 ( .A(n37562), .B(n24851), .Y(n24849) );
  AND2X1 U24297 ( .A(n44086), .B(mem_i_inst_i[1]), .Y(n24851) );
  NOR2X1 U24298 ( .A(n24572), .B(n611), .Y(n24848) );
  NAND2X1 U24299 ( .A(n24852), .B(n24853), .Y(n24574) );
  NAND2X1 U24300 ( .A(mem_i_inst_i[2]), .B(n44085), .Y(n24853) );
  AND2X1 U24302 ( .A(n24854), .B(n24855), .Y(n24572) );
  NOR2X1 U24304 ( .A(n37562), .B(n24856), .Y(n24854) );
  AND2X1 U24305 ( .A(n44086), .B(mem_i_inst_i[0]), .Y(n24856) );
  NAND2X1 U24311 ( .A(n24861), .B(n24862), .Y(u_csr_result_r[9]) );
  NOR2X1 U24312 ( .A(n24863), .B(n24864), .Y(n24862) );
  NAND2X1 U24313 ( .A(n24865), .B(n24866), .Y(n24864) );
  NAND2X1 U24314 ( .A(n457), .B(n73413), .Y(n24866) );
  NOR2X1 U24315 ( .A(n24867), .B(n24868), .Y(n24865) );
  NOR2X1 U24316 ( .A(n44297), .B(n1165), .Y(n24868) );
  NOR2X1 U24317 ( .A(n44293), .B(n37726), .Y(n24867) );
  NAND2X1 U24318 ( .A(n24871), .B(n24872), .Y(n24863) );
  NOR2X1 U24319 ( .A(n24873), .B(n24874), .Y(n24872) );
  NOR2X1 U24320 ( .A(n44292), .B(n37694), .Y(n24874) );
  NOR2X1 U24321 ( .A(n24876), .B(n24877), .Y(n24873) );
  NOR2X1 U24322 ( .A(n24878), .B(n24879), .Y(n24876) );
  NOR2X1 U24323 ( .A(n889), .B(n37549), .Y(n24879) );
  NOR2X1 U24324 ( .A(n896), .B(n37334), .Y(n24878) );
  AND2X1 U24325 ( .A(n24880), .B(n24881), .Y(n24871) );
  NAND2X1 U24326 ( .A(cpu_id_i[9]), .B(n44288), .Y(n24881) );
  NAND2X1 U24327 ( .A(u_csr_csr_sr_q[9]), .B(n42144), .Y(n24880) );
  NOR2X1 U24328 ( .A(n24884), .B(n24885), .Y(n24861) );
  NAND2X1 U24329 ( .A(n24886), .B(n24887), .Y(n24885) );
  NAND2X1 U24330 ( .A(n42205), .B(u_csr_csr_mideleg_q[9]), .Y(n24887) );
  NOR2X1 U24331 ( .A(n24889), .B(n24890), .Y(n24886) );
  NOR2X1 U24332 ( .A(n42982), .B(n37716), .Y(n24890) );
  NAND2X1 U24334 ( .A(n24892), .B(n24893), .Y(n24884) );
  NOR2X1 U24335 ( .A(n24894), .B(n24895), .Y(n24893) );
  AND2X1 U24337 ( .A(n44079), .B(u_csr_csr_stval_q[9]), .Y(n24894) );
  NOR2X1 U24338 ( .A(n24898), .B(n24899), .Y(n24892) );
  AND2X1 U24339 ( .A(n73399), .B(u_csr_csr_medeleg_q[9]), .Y(n24899) );
  AND2X1 U24340 ( .A(n42848), .B(u_csr_csr_mscratch_q[9]), .Y(n24898) );
  NAND2X1 U24341 ( .A(n24900), .B(n24901), .Y(u_csr_result_r[8]) );
  NOR2X1 U24342 ( .A(n24902), .B(n24903), .Y(n24901) );
  NAND2X1 U24343 ( .A(n24904), .B(n24905), .Y(n24903) );
  NAND2X1 U24344 ( .A(n457), .B(n73414), .Y(n24905) );
  NOR2X1 U24345 ( .A(n24906), .B(n24907), .Y(n24904) );
  NOR2X1 U24346 ( .A(n44297), .B(n1166), .Y(n24907) );
  NOR2X1 U24347 ( .A(n44293), .B(n37725), .Y(n24906) );
  NAND2X1 U24348 ( .A(n24908), .B(n24909), .Y(n24902) );
  NOR2X1 U24349 ( .A(n24910), .B(n24911), .Y(n24909) );
  NOR2X1 U24350 ( .A(n44292), .B(n37571), .Y(n24911) );
  AND2X1 U24351 ( .A(n24912), .B(n24913), .Y(n24908) );
  NAND2X1 U24352 ( .A(cpu_id_i[8]), .B(n44288), .Y(n24913) );
  NAND2X1 U24353 ( .A(u_csr_csr_sr_q[8]), .B(n458), .Y(n24912) );
  NOR2X1 U24354 ( .A(n24914), .B(n24915), .Y(n24900) );
  NAND2X1 U24355 ( .A(n24916), .B(n24917), .Y(n24915) );
  NAND2X1 U24356 ( .A(u_csr_csr_mideleg_q[8]), .B(n42205), .Y(n24917) );
  NOR2X1 U24357 ( .A(n24918), .B(n24919), .Y(n24916) );
  NOR2X1 U24358 ( .A(n42982), .B(n37710), .Y(n24919) );
  NAND2X1 U24360 ( .A(n24920), .B(n24921), .Y(n24914) );
  NOR2X1 U24361 ( .A(n24922), .B(n24923), .Y(n24921) );
  AND2X1 U24363 ( .A(n44079), .B(u_csr_csr_stval_q[8]), .Y(n24922) );
  NOR2X1 U24364 ( .A(n24924), .B(n24925), .Y(n24920) );
  AND2X1 U24365 ( .A(n73399), .B(u_csr_csr_medeleg_q[8]), .Y(n24925) );
  AND2X1 U24366 ( .A(n42849), .B(u_csr_csr_mscratch_q[8]), .Y(n24924) );
  NAND2X1 U24367 ( .A(n24926), .B(n24927), .Y(u_csr_result_r[7]) );
  NOR2X1 U24368 ( .A(n24928), .B(n24929), .Y(n24927) );
  NAND2X1 U24369 ( .A(n24930), .B(n24931), .Y(n24929) );
  NAND2X1 U24370 ( .A(n457), .B(n73415), .Y(n24931) );
  NOR2X1 U24371 ( .A(n24932), .B(n24933), .Y(n24930) );
  NOR2X1 U24372 ( .A(n44297), .B(n1167), .Y(n24933) );
  NOR2X1 U24373 ( .A(n44293), .B(n37724), .Y(n24932) );
  NAND2X1 U24374 ( .A(n24934), .B(n24935), .Y(n24928) );
  NOR2X1 U24375 ( .A(n24936), .B(n24937), .Y(n24935) );
  NOR2X1 U24376 ( .A(n44292), .B(n37346), .Y(n24937) );
  NOR2X1 U24378 ( .A(n24940), .B(n24941), .Y(n24938) );
  NOR2X1 U24379 ( .A(n37330), .B(n24942), .Y(n24941) );
  NOR2X1 U24380 ( .A(n37545), .B(n24943), .Y(n24940) );
  AND2X1 U24381 ( .A(n24944), .B(n24945), .Y(n24934) );
  NAND2X1 U24382 ( .A(cpu_id_i[7]), .B(n44288), .Y(n24945) );
  NAND2X1 U24383 ( .A(u_csr_csr_sr_q[7]), .B(n42144), .Y(n24944) );
  NOR2X1 U24384 ( .A(n24946), .B(n24947), .Y(n24926) );
  NAND2X1 U24385 ( .A(n24948), .B(n24949), .Y(n24947) );
  NAND2X1 U24386 ( .A(n42205), .B(u_csr_csr_mideleg_q[7]), .Y(n24949) );
  NOR2X1 U24387 ( .A(n24950), .B(n24951), .Y(n24948) );
  NOR2X1 U24388 ( .A(n42983), .B(n37715), .Y(n24951) );
  NAND2X1 U24390 ( .A(n24952), .B(n24953), .Y(n24946) );
  NOR2X1 U24391 ( .A(n24954), .B(n24955), .Y(n24953) );
  AND2X1 U24393 ( .A(n44079), .B(u_csr_csr_stval_q[7]), .Y(n24954) );
  NOR2X1 U24394 ( .A(n24956), .B(n24957), .Y(n24952) );
  NOR2X1 U24395 ( .A(n24958), .B(n37566), .Y(n24957) );
  AND2X1 U24396 ( .A(n42849), .B(u_csr_csr_mscratch_q[7]), .Y(n24956) );
  NAND2X1 U24397 ( .A(n24959), .B(n24960), .Y(u_csr_result_r[6]) );
  NOR2X1 U24398 ( .A(n24961), .B(n24962), .Y(n24960) );
  NAND2X1 U24399 ( .A(n24963), .B(n24964), .Y(n24962) );
  NAND2X1 U24400 ( .A(u_csr_csr_stval_q[6]), .B(n44078), .Y(n24964) );
  NOR2X1 U24401 ( .A(n24965), .B(n24966), .Y(n24963) );
  NOR2X1 U24402 ( .A(n1898), .B(n40682), .Y(n24966) );
  NOR2X1 U24403 ( .A(n44297), .B(n1168), .Y(n24965) );
  NAND2X1 U24404 ( .A(n24968), .B(n24969), .Y(n24961) );
  NOR2X1 U24405 ( .A(n24970), .B(n24971), .Y(n24969) );
  AND2X1 U24406 ( .A(cpu_id_i[6]), .B(n44289), .Y(n24971) );
  NOR2X1 U24407 ( .A(n44292), .B(n37569), .Y(n24970) );
  NOR2X1 U24408 ( .A(n24972), .B(n24973), .Y(n24968) );
  NOR2X1 U24409 ( .A(n44293), .B(n1137), .Y(n24973) );
  AND2X1 U24410 ( .A(n44286), .B(u_csr_csr_sr_q[6]), .Y(n24972) );
  NOR2X1 U24411 ( .A(n24974), .B(n24975), .Y(n24959) );
  NAND2X1 U24412 ( .A(n24976), .B(n24977), .Y(n24975) );
  NAND2X1 U24413 ( .A(u_csr_csr_mideleg_q[6]), .B(n42205), .Y(n24977) );
  NOR2X1 U24414 ( .A(n24978), .B(n24979), .Y(n24976) );
  NOR2X1 U24415 ( .A(n42982), .B(n37706), .Y(n24979) );
  NAND2X1 U24417 ( .A(n24980), .B(n24981), .Y(n24974) );
  NAND2X1 U24418 ( .A(u_csr_csr_medeleg_q[6]), .B(n73399), .Y(n24981) );
  NOR2X1 U24419 ( .A(n24982), .B(n24983), .Y(n24980) );
  AND2X1 U24420 ( .A(n42848), .B(u_csr_csr_mscratch_q[6]), .Y(n24983) );
  NAND2X1 U24422 ( .A(n24984), .B(n24985), .Y(u_csr_result_r[5]) );
  NOR2X1 U24423 ( .A(n24986), .B(n24987), .Y(n24985) );
  NAND2X1 U24424 ( .A(n24988), .B(n24989), .Y(n24987) );
  NAND2X1 U24425 ( .A(n457), .B(n73416), .Y(n24989) );
  NOR2X1 U24426 ( .A(n24990), .B(n24991), .Y(n24988) );
  NOR2X1 U24427 ( .A(n44296), .B(n1169), .Y(n24991) );
  NOR2X1 U24428 ( .A(n44293), .B(n1138), .Y(n24990) );
  NAND2X1 U24429 ( .A(n24992), .B(n24993), .Y(n24986) );
  NOR2X1 U24430 ( .A(n24994), .B(n24995), .Y(n24993) );
  NOR2X1 U24431 ( .A(n44292), .B(n37345), .Y(n24995) );
  NOR2X1 U24432 ( .A(n24996), .B(n24877), .Y(n24994) );
  NOR2X1 U24433 ( .A(n24997), .B(n24998), .Y(n24996) );
  NOR2X1 U24434 ( .A(n889), .B(n37331), .Y(n24998) );
  NOR2X1 U24435 ( .A(n896), .B(n37546), .Y(n24997) );
  AND2X1 U24436 ( .A(n24999), .B(n25000), .Y(n24992) );
  NAND2X1 U24437 ( .A(cpu_id_i[5]), .B(n44288), .Y(n25000) );
  NAND2X1 U24438 ( .A(u_csr_csr_sr_q[5]), .B(n458), .Y(n24999) );
  NOR2X1 U24439 ( .A(n25001), .B(n25002), .Y(n24984) );
  NAND2X1 U24440 ( .A(n25003), .B(n25004), .Y(n25002) );
  NAND2X1 U24441 ( .A(n42205), .B(u_csr_csr_mideleg_q[5]), .Y(n25004) );
  NOR2X1 U24442 ( .A(n25005), .B(n25006), .Y(n25003) );
  NOR2X1 U24443 ( .A(n42982), .B(n37714), .Y(n25006) );
  NAND2X1 U24445 ( .A(n25007), .B(n25008), .Y(n25001) );
  NOR2X1 U24446 ( .A(n25009), .B(n25010), .Y(n25008) );
  AND2X1 U24448 ( .A(n44079), .B(u_csr_csr_stval_q[5]), .Y(n25009) );
  NOR2X1 U24449 ( .A(n25011), .B(n25012), .Y(n25007) );
  AND2X1 U24450 ( .A(n73399), .B(u_csr_csr_medeleg_q[5]), .Y(n25012) );
  AND2X1 U24451 ( .A(n42849), .B(u_csr_csr_mscratch_q[5]), .Y(n25011) );
  NAND2X1 U24452 ( .A(n25013), .B(n25014), .Y(u_csr_result_r[4]) );
  NOR2X1 U24453 ( .A(n25015), .B(n25016), .Y(n25014) );
  NAND2X1 U24454 ( .A(n25017), .B(n25018), .Y(n25016) );
  NAND2X1 U24455 ( .A(u_csr_csr_stval_q[4]), .B(n44078), .Y(n25018) );
  NOR2X1 U24456 ( .A(n25019), .B(n25020), .Y(n25017) );
  NOR2X1 U24457 ( .A(n1899), .B(n40681), .Y(n25020) );
  NOR2X1 U24458 ( .A(n44296), .B(n37701), .Y(n25019) );
  NAND2X1 U24459 ( .A(n25021), .B(n25022), .Y(n25015) );
  NOR2X1 U24460 ( .A(n25023), .B(n25024), .Y(n25022) );
  AND2X1 U24461 ( .A(cpu_id_i[4]), .B(n44289), .Y(n25024) );
  NOR2X1 U24462 ( .A(n44292), .B(n37721), .Y(n25023) );
  NOR2X1 U24463 ( .A(n25025), .B(n25026), .Y(n25021) );
  NOR2X1 U24464 ( .A(n44293), .B(n1139), .Y(n25026) );
  AND2X1 U24465 ( .A(n458), .B(u_csr_csr_sr_q[4]), .Y(n25025) );
  NOR2X1 U24466 ( .A(n25027), .B(n25028), .Y(n25013) );
  NAND2X1 U24467 ( .A(n25029), .B(n25030), .Y(n25028) );
  NAND2X1 U24468 ( .A(u_csr_csr_mideleg_q[4]), .B(n42205), .Y(n25030) );
  NOR2X1 U24469 ( .A(n25031), .B(n25032), .Y(n25029) );
  NOR2X1 U24470 ( .A(n42983), .B(n37705), .Y(n25032) );
  NAND2X1 U24472 ( .A(n25033), .B(n25034), .Y(n25027) );
  NAND2X1 U24473 ( .A(u_csr_csr_medeleg_q[4]), .B(n73399), .Y(n25034) );
  NOR2X1 U24474 ( .A(n25035), .B(n25036), .Y(n25033) );
  AND2X1 U24475 ( .A(n42849), .B(u_csr_csr_mscratch_q[4]), .Y(n25036) );
  NAND2X1 U24477 ( .A(n25037), .B(n25038), .Y(u_csr_result_r[3]) );
  NOR2X1 U24478 ( .A(n25039), .B(n25040), .Y(n25038) );
  NAND2X1 U24479 ( .A(n25041), .B(n25042), .Y(n25040) );
  AND2X1 U24480 ( .A(n25043), .B(n25044), .Y(n25042) );
  NAND2X1 U24481 ( .A(cpu_id_i[3]), .B(n44288), .Y(n25044) );
  NAND2X1 U24482 ( .A(u_csr_csr_sr_q[3]), .B(n44286), .Y(n25043) );
  NOR2X1 U24483 ( .A(n25045), .B(n25046), .Y(n25041) );
  NOR2X1 U24484 ( .A(n44296), .B(n37723), .Y(n25046) );
  NOR2X1 U24485 ( .A(n44293), .B(n1140), .Y(n25045) );
  NAND2X1 U24486 ( .A(n25047), .B(n25048), .Y(n25039) );
  NOR2X1 U24487 ( .A(n25049), .B(n25050), .Y(n25048) );
  AND2X1 U24488 ( .A(n73400), .B(u_csr_csr_scause_q[3]), .Y(n25050) );
  NOR2X1 U24490 ( .A(n25052), .B(n25053), .Y(n25051) );
  NOR2X1 U24491 ( .A(n37544), .B(n24942), .Y(n25053) );
  NOR2X1 U24492 ( .A(n37335), .B(n24943), .Y(n25052) );
  NOR2X1 U24493 ( .A(n25054), .B(n25055), .Y(n25047) );
  NOR2X1 U24494 ( .A(n44292), .B(n37693), .Y(n25055) );
  AND2X1 U24495 ( .A(n42145), .B(u_csr_csr_mcause_q[3]), .Y(n25054) );
  NOR2X1 U24496 ( .A(n25057), .B(n25058), .Y(n25037) );
  NAND2X1 U24497 ( .A(n25059), .B(n25060), .Y(n25058) );
  NOR2X1 U24498 ( .A(n25061), .B(n25062), .Y(n25060) );
  AND2X1 U24500 ( .A(n73399), .B(u_csr_csr_medeleg_q[3]), .Y(n25061) );
  NOR2X1 U24501 ( .A(n25063), .B(n25064), .Y(n25059) );
  AND2X1 U24502 ( .A(u_csr_csr_mideleg_q[3]), .B(n42205), .Y(n25064) );
  NOR2X1 U24503 ( .A(n42982), .B(n37700), .Y(n25063) );
  NAND2X1 U24504 ( .A(n25065), .B(n25066), .Y(n25057) );
  NOR2X1 U24505 ( .A(n25067), .B(n25068), .Y(n25066) );
  AND2X1 U24506 ( .A(n44079), .B(u_csr_csr_stval_q[3]), .Y(n25068) );
  NOR2X1 U24507 ( .A(n1895), .B(n40682), .Y(n25067) );
  NOR2X1 U24508 ( .A(n25069), .B(n25070), .Y(n25065) );
  AND2X1 U24509 ( .A(n42848), .B(u_csr_csr_mscratch_q[3]), .Y(n25070) );
  NAND2X1 U24511 ( .A(n25071), .B(n25072), .Y(u_csr_result_r[31]) );
  NOR2X1 U24512 ( .A(n25073), .B(n25074), .Y(n25072) );
  NAND2X1 U24513 ( .A(n25075), .B(n25076), .Y(n25074) );
  NAND2X1 U24514 ( .A(u_csr_csr_stvec_q[31]), .B(n36765), .Y(n25076) );
  NOR2X1 U24515 ( .A(n25077), .B(n25078), .Y(n25075) );
  NOR2X1 U24516 ( .A(n44293), .B(n1141), .Y(n25078) );
  AND2X1 U24517 ( .A(n44286), .B(u_csr_csr_sr_q_31), .Y(n25077) );
  NAND2X1 U24518 ( .A(n25079), .B(n25080), .Y(n25073) );
  NOR2X1 U24519 ( .A(n25081), .B(n25082), .Y(n25080) );
  AND2X1 U24520 ( .A(n42145), .B(u_csr_csr_mcause_q_31), .Y(n25082) );
  AND2X1 U24521 ( .A(n73400), .B(u_csr_csr_scause_q_31), .Y(n25081) );
  NOR2X1 U24522 ( .A(n25084), .B(n25085), .Y(n25079) );
  AND2X1 U24523 ( .A(cpu_id_i[31]), .B(n44289), .Y(n25085) );
  NOR2X1 U24524 ( .A(n44292), .B(n37729), .Y(n25084) );
  NOR2X1 U24525 ( .A(n25086), .B(n25087), .Y(n25071) );
  NAND2X1 U24526 ( .A(n25088), .B(n25089), .Y(n25087) );
  NAND2X1 U24527 ( .A(u_csr_csr_mtvec_q[31]), .B(n41738), .Y(n25089) );
  NOR2X1 U24528 ( .A(n25090), .B(n25091), .Y(n25088) );
  AND2X1 U24530 ( .A(n42848), .B(u_csr_csr_mscratch_q[31]), .Y(n25090) );
  NAND2X1 U24531 ( .A(n25092), .B(n25093), .Y(n25086) );
  NOR2X1 U24533 ( .A(n25094), .B(n25095), .Y(n25092) );
  AND2X1 U24534 ( .A(n44079), .B(u_csr_csr_stval_q[31]), .Y(n25095) );
  AND2X1 U24535 ( .A(u_csr_csr_satp_q_31_), .B(n457), .Y(n25094) );
  NAND2X1 U24536 ( .A(n25096), .B(n25097), .Y(u_csr_result_r[30]) );
  NOR2X1 U24537 ( .A(n25098), .B(n25099), .Y(n25097) );
  NAND2X1 U24538 ( .A(n25100), .B(n25101), .Y(n25099) );
  NAND2X1 U24539 ( .A(u_csr_csr_stvec_q[30]), .B(n36765), .Y(n25101) );
  NOR2X1 U24540 ( .A(n25102), .B(n25103), .Y(n25100) );
  NOR2X1 U24541 ( .A(n44293), .B(n1142), .Y(n25103) );
  AND2X1 U24542 ( .A(n44286), .B(u_csr_csr_sr_q_30), .Y(n25102) );
  NAND2X1 U24543 ( .A(n25104), .B(n25105), .Y(n25098) );
  NAND2X1 U24544 ( .A(cpu_id_i[30]), .B(n44288), .Y(n25105) );
  NOR2X1 U24545 ( .A(n24910), .B(n25106), .Y(n25104) );
  NOR2X1 U24546 ( .A(n44291), .B(n37699), .Y(n25106) );
  NOR2X1 U24547 ( .A(n25107), .B(n25108), .Y(n25096) );
  NAND2X1 U24548 ( .A(n25109), .B(n25110), .Y(n25108) );
  NAND2X1 U24549 ( .A(u_csr_csr_mtvec_q[30]), .B(n41738), .Y(n25110) );
  NOR2X1 U24550 ( .A(n25111), .B(n25112), .Y(n25109) );
  AND2X1 U24552 ( .A(n42849), .B(u_csr_csr_mscratch_q[30]), .Y(n25111) );
  NAND2X1 U24553 ( .A(n25113), .B(n25114), .Y(n25107) );
  NOR2X1 U24555 ( .A(n25115), .B(n25116), .Y(n25113) );
  AND2X1 U24556 ( .A(n44079), .B(u_csr_csr_stval_q[30]), .Y(n25116) );
  NOR2X1 U24557 ( .A(n1902), .B(n40681), .Y(n25115) );
  NAND2X1 U24558 ( .A(n25117), .B(n25118), .Y(u_csr_result_r[2]) );
  NOR2X1 U24559 ( .A(n25119), .B(n25120), .Y(n25118) );
  NAND2X1 U24560 ( .A(n25121), .B(n25122), .Y(n25120) );
  NOR2X1 U24561 ( .A(n25123), .B(n25124), .Y(n25122) );
  NOR2X1 U24562 ( .A(n44293), .B(n1143), .Y(n25124) );
  AND2X1 U24563 ( .A(n44286), .B(u_csr_csr_sr_q[2]), .Y(n25123) );
  NOR2X1 U24564 ( .A(n25125), .B(n25126), .Y(n25121) );
  NOR2X1 U24565 ( .A(n1903), .B(n40681), .Y(n25126) );
  NOR2X1 U24566 ( .A(n44296), .B(n37703), .Y(n25125) );
  NAND2X1 U24567 ( .A(n25127), .B(n25128), .Y(n25119) );
  NOR2X1 U24568 ( .A(n25129), .B(n25130), .Y(n25128) );
  AND2X1 U24569 ( .A(n42145), .B(u_csr_csr_mcause_q[2]), .Y(n25130) );
  NOR2X1 U24570 ( .A(n25083), .B(n37728), .Y(n25129) );
  NOR2X1 U24571 ( .A(n25131), .B(n25132), .Y(n25127) );
  AND2X1 U24572 ( .A(cpu_id_i[2]), .B(n44289), .Y(n25132) );
  NOR2X1 U24573 ( .A(n44291), .B(n37563), .Y(n25131) );
  NOR2X1 U24574 ( .A(n25133), .B(n25134), .Y(n25117) );
  NAND2X1 U24575 ( .A(n25135), .B(n25136), .Y(n25134) );
  NAND2X1 U24576 ( .A(u_csr_csr_mideleg_q[2]), .B(n42205), .Y(n25136) );
  NOR2X1 U24577 ( .A(n25137), .B(n25138), .Y(n25135) );
  NOR2X1 U24578 ( .A(n42982), .B(n37709), .Y(n25138) );
  NAND2X1 U24580 ( .A(n25139), .B(n25140), .Y(n25133) );
  NOR2X1 U24581 ( .A(n25141), .B(n25142), .Y(n25140) );
  AND2X1 U24583 ( .A(n44079), .B(u_csr_csr_stval_q[2]), .Y(n25141) );
  NOR2X1 U24584 ( .A(n25143), .B(n25144), .Y(n25139) );
  AND2X1 U24585 ( .A(n73399), .B(u_csr_csr_medeleg_q[2]), .Y(n25144) );
  AND2X1 U24586 ( .A(n42848), .B(u_csr_csr_mscratch_q[2]), .Y(n25143) );
  NAND2X1 U24587 ( .A(n25145), .B(n25146), .Y(u_csr_result_r[29]) );
  NOR2X1 U24588 ( .A(n25147), .B(n25148), .Y(n25146) );
  NAND2X1 U24589 ( .A(n25149), .B(n25150), .Y(n25148) );
  NAND2X1 U24590 ( .A(n457), .B(n73559), .Y(n25150) );
  NOR2X1 U24591 ( .A(n25151), .B(n25152), .Y(n25149) );
  NOR2X1 U24592 ( .A(n44296), .B(n1175), .Y(n25152) );
  NOR2X1 U24593 ( .A(n44293), .B(n1144), .Y(n25151) );
  NAND2X1 U24594 ( .A(n25153), .B(n25154), .Y(n25147) );
  NAND2X1 U24595 ( .A(u_csr_csr_sr_q_29), .B(n42144), .Y(n25154) );
  NOR2X1 U24596 ( .A(n25155), .B(n25156), .Y(n25153) );
  AND2X1 U24597 ( .A(cpu_id_i[29]), .B(n44289), .Y(n25156) );
  NOR2X1 U24598 ( .A(n44291), .B(n37695), .Y(n25155) );
  NOR2X1 U24599 ( .A(n25157), .B(n25158), .Y(n25145) );
  NAND2X1 U24600 ( .A(n25159), .B(n25160), .Y(n25158) );
  NAND2X1 U24602 ( .A(u_csr_csr_mtvec_q[29]), .B(n41738), .Y(n25159) );
  NAND2X1 U24603 ( .A(n25161), .B(n25162), .Y(n25157) );
  NAND2X1 U24604 ( .A(u_csr_csr_mscratch_q[29]), .B(n44080), .Y(n25162) );
  NOR2X1 U24605 ( .A(n25163), .B(n25164), .Y(n25161) );
  AND2X1 U24607 ( .A(n44079), .B(u_csr_csr_stval_q[29]), .Y(n25163) );
  NAND2X1 U24608 ( .A(n25165), .B(n25166), .Y(u_csr_result_r[28]) );
  NOR2X1 U24609 ( .A(n25167), .B(n25168), .Y(n25166) );
  NAND2X1 U24610 ( .A(n25169), .B(n25170), .Y(n25168) );
  NAND2X1 U24611 ( .A(n457), .B(n73560), .Y(n25170) );
  NOR2X1 U24612 ( .A(n25171), .B(n25172), .Y(n25169) );
  NOR2X1 U24613 ( .A(n44296), .B(n1176), .Y(n25172) );
  NOR2X1 U24614 ( .A(n44293), .B(n1145), .Y(n25171) );
  NAND2X1 U24615 ( .A(n25173), .B(n25174), .Y(n25167) );
  NAND2X1 U24616 ( .A(u_csr_csr_sr_q_28), .B(n42144), .Y(n25174) );
  NOR2X1 U24617 ( .A(n25175), .B(n25176), .Y(n25173) );
  AND2X1 U24618 ( .A(cpu_id_i[28]), .B(n44289), .Y(n25176) );
  NOR2X1 U24619 ( .A(n44291), .B(n37598), .Y(n25175) );
  NOR2X1 U24620 ( .A(n25177), .B(n25178), .Y(n25165) );
  NAND2X1 U24621 ( .A(n25179), .B(n25180), .Y(n25178) );
  NAND2X1 U24623 ( .A(u_csr_csr_mtvec_q[28]), .B(n41738), .Y(n25179) );
  NAND2X1 U24624 ( .A(n25181), .B(n25182), .Y(n25177) );
  NAND2X1 U24625 ( .A(u_csr_csr_mscratch_q[28]), .B(n42848), .Y(n25182) );
  NOR2X1 U24626 ( .A(n25183), .B(n25184), .Y(n25181) );
  AND2X1 U24628 ( .A(n44079), .B(u_csr_csr_stval_q[28]), .Y(n25183) );
  NAND2X1 U24629 ( .A(n25185), .B(n25186), .Y(u_csr_result_r[27]) );
  NOR2X1 U24630 ( .A(n25187), .B(n25188), .Y(n25186) );
  NAND2X1 U24631 ( .A(n25189), .B(n25190), .Y(n25188) );
  NAND2X1 U24632 ( .A(n457), .B(n73561), .Y(n25190) );
  NOR2X1 U24633 ( .A(n25191), .B(n25192), .Y(n25189) );
  NOR2X1 U24634 ( .A(n44296), .B(n1177), .Y(n25192) );
  NOR2X1 U24635 ( .A(n44293), .B(n1146), .Y(n25191) );
  NAND2X1 U24636 ( .A(n25193), .B(n25194), .Y(n25187) );
  NAND2X1 U24637 ( .A(u_csr_csr_sr_q_27), .B(n42144), .Y(n25194) );
  NOR2X1 U24638 ( .A(n25195), .B(n25196), .Y(n25193) );
  AND2X1 U24639 ( .A(cpu_id_i[27]), .B(n44289), .Y(n25196) );
  NOR2X1 U24640 ( .A(n44291), .B(n37352), .Y(n25195) );
  NOR2X1 U24641 ( .A(n25197), .B(n25198), .Y(n25185) );
  NAND2X1 U24642 ( .A(n25199), .B(n25200), .Y(n25198) );
  NAND2X1 U24644 ( .A(u_csr_csr_mtvec_q[27]), .B(n41738), .Y(n25199) );
  NAND2X1 U24645 ( .A(n25201), .B(n25202), .Y(n25197) );
  NAND2X1 U24646 ( .A(u_csr_csr_mscratch_q[27]), .B(n44080), .Y(n25202) );
  NOR2X1 U24647 ( .A(n25203), .B(n25204), .Y(n25201) );
  AND2X1 U24649 ( .A(n44079), .B(u_csr_csr_stval_q[27]), .Y(n25203) );
  NAND2X1 U24650 ( .A(n25205), .B(n25206), .Y(u_csr_result_r[26]) );
  NOR2X1 U24651 ( .A(n25207), .B(n25208), .Y(n25206) );
  NAND2X1 U24652 ( .A(n25209), .B(n25210), .Y(n25208) );
  NAND2X1 U24653 ( .A(n457), .B(n73562), .Y(n25210) );
  NOR2X1 U24654 ( .A(n25211), .B(n25212), .Y(n25209) );
  NOR2X1 U24655 ( .A(n44296), .B(n1178), .Y(n25212) );
  NOR2X1 U24656 ( .A(n44293), .B(n1147), .Y(n25211) );
  NAND2X1 U24657 ( .A(n25213), .B(n25214), .Y(n25207) );
  NAND2X1 U24658 ( .A(u_csr_csr_sr_q_26), .B(n42144), .Y(n25214) );
  NOR2X1 U24659 ( .A(n25215), .B(n25216), .Y(n25213) );
  AND2X1 U24660 ( .A(cpu_id_i[26]), .B(n44289), .Y(n25216) );
  NOR2X1 U24661 ( .A(n44291), .B(n37698), .Y(n25215) );
  NOR2X1 U24662 ( .A(n25217), .B(n25218), .Y(n25205) );
  NAND2X1 U24663 ( .A(n25219), .B(n25220), .Y(n25218) );
  NAND2X1 U24665 ( .A(u_csr_csr_mtvec_q[26]), .B(n41738), .Y(n25219) );
  NAND2X1 U24666 ( .A(n25221), .B(n25222), .Y(n25217) );
  NAND2X1 U24667 ( .A(u_csr_csr_mscratch_q[26]), .B(n44080), .Y(n25222) );
  NOR2X1 U24668 ( .A(n25223), .B(n25224), .Y(n25221) );
  AND2X1 U24670 ( .A(n44079), .B(u_csr_csr_stval_q[26]), .Y(n25223) );
  NAND2X1 U24671 ( .A(n25225), .B(n25226), .Y(u_csr_result_r[25]) );
  NOR2X1 U24672 ( .A(n25227), .B(n25228), .Y(n25226) );
  NAND2X1 U24673 ( .A(n25229), .B(n25230), .Y(n25228) );
  NAND2X1 U24674 ( .A(n457), .B(n73563), .Y(n25230) );
  NOR2X1 U24675 ( .A(n25231), .B(n25232), .Y(n25229) );
  NOR2X1 U24676 ( .A(n44296), .B(n1179), .Y(n25232) );
  NOR2X1 U24677 ( .A(n44293), .B(n1148), .Y(n25231) );
  NAND2X1 U24678 ( .A(n25233), .B(n25234), .Y(n25227) );
  NAND2X1 U24679 ( .A(u_csr_csr_sr_q_25), .B(n42144), .Y(n25234) );
  NOR2X1 U24680 ( .A(n25235), .B(n25236), .Y(n25233) );
  AND2X1 U24681 ( .A(cpu_id_i[25]), .B(n44289), .Y(n25236) );
  NOR2X1 U24682 ( .A(n44291), .B(n37691), .Y(n25235) );
  NOR2X1 U24683 ( .A(n25237), .B(n25238), .Y(n25225) );
  NAND2X1 U24684 ( .A(n25239), .B(n25240), .Y(n25238) );
  NAND2X1 U24686 ( .A(u_csr_csr_mtvec_q[25]), .B(n41738), .Y(n25239) );
  NAND2X1 U24687 ( .A(n25241), .B(n25242), .Y(n25237) );
  NAND2X1 U24688 ( .A(u_csr_csr_mscratch_q[25]), .B(n44080), .Y(n25242) );
  NOR2X1 U24689 ( .A(n25243), .B(n25244), .Y(n25241) );
  AND2X1 U24691 ( .A(n44079), .B(u_csr_csr_stval_q[25]), .Y(n25243) );
  NAND2X1 U24692 ( .A(n25245), .B(n25246), .Y(u_csr_result_r[24]) );
  NOR2X1 U24693 ( .A(n25247), .B(n25248), .Y(n25246) );
  NAND2X1 U24694 ( .A(n25249), .B(n25250), .Y(n25248) );
  NAND2X1 U24695 ( .A(n457), .B(n73564), .Y(n25250) );
  NOR2X1 U24696 ( .A(n25251), .B(n25252), .Y(n25249) );
  NOR2X1 U24697 ( .A(n44296), .B(n1180), .Y(n25252) );
  NOR2X1 U24698 ( .A(n44293), .B(n1149), .Y(n25251) );
  NAND2X1 U24699 ( .A(n25253), .B(n25254), .Y(n25247) );
  NAND2X1 U24700 ( .A(u_csr_csr_sr_q_24), .B(n42144), .Y(n25254) );
  NOR2X1 U24701 ( .A(n25255), .B(n25256), .Y(n25253) );
  AND2X1 U24702 ( .A(cpu_id_i[24]), .B(n44289), .Y(n25256) );
  NOR2X1 U24703 ( .A(n44291), .B(n37588), .Y(n25255) );
  NOR2X1 U24704 ( .A(n25257), .B(n25258), .Y(n25245) );
  NAND2X1 U24705 ( .A(n25259), .B(n25260), .Y(n25258) );
  NAND2X1 U24707 ( .A(u_csr_csr_mtvec_q[24]), .B(n41738), .Y(n25259) );
  NAND2X1 U24708 ( .A(n25261), .B(n25262), .Y(n25257) );
  NAND2X1 U24709 ( .A(u_csr_csr_mscratch_q[24]), .B(n44080), .Y(n25262) );
  NOR2X1 U24710 ( .A(n25263), .B(n25264), .Y(n25261) );
  AND2X1 U24712 ( .A(n44079), .B(u_csr_csr_stval_q[24]), .Y(n25263) );
  NAND2X1 U24713 ( .A(n25265), .B(n25266), .Y(u_csr_result_r[23]) );
  NOR2X1 U24714 ( .A(n25267), .B(n25268), .Y(n25266) );
  NAND2X1 U24715 ( .A(n25269), .B(n25270), .Y(n25268) );
  NAND2X1 U24716 ( .A(n457), .B(n73565), .Y(n25270) );
  NOR2X1 U24717 ( .A(n25271), .B(n25272), .Y(n25269) );
  NOR2X1 U24718 ( .A(n44296), .B(n1181), .Y(n25272) );
  NOR2X1 U24719 ( .A(n44293), .B(n1150), .Y(n25271) );
  NAND2X1 U24720 ( .A(n25273), .B(n25274), .Y(n25267) );
  NAND2X1 U24721 ( .A(u_csr_csr_sr_q_23), .B(n42144), .Y(n25274) );
  NOR2X1 U24722 ( .A(n25275), .B(n25276), .Y(n25273) );
  AND2X1 U24723 ( .A(cpu_id_i[23]), .B(n44289), .Y(n25276) );
  NOR2X1 U24724 ( .A(n44291), .B(n37350), .Y(n25275) );
  NOR2X1 U24725 ( .A(n25277), .B(n25278), .Y(n25265) );
  NAND2X1 U24726 ( .A(n25279), .B(n25280), .Y(n25278) );
  NAND2X1 U24728 ( .A(u_csr_csr_mtvec_q[23]), .B(n41738), .Y(n25279) );
  NAND2X1 U24729 ( .A(n25281), .B(n25282), .Y(n25277) );
  NAND2X1 U24730 ( .A(u_csr_csr_mscratch_q[23]), .B(n44080), .Y(n25282) );
  NOR2X1 U24731 ( .A(n25283), .B(n25284), .Y(n25281) );
  AND2X1 U24733 ( .A(n44079), .B(u_csr_csr_stval_q[23]), .Y(n25283) );
  NAND2X1 U24734 ( .A(n25285), .B(n25286), .Y(u_csr_result_r[22]) );
  NOR2X1 U24735 ( .A(n25287), .B(n25288), .Y(n25286) );
  NAND2X1 U24736 ( .A(n25289), .B(n25290), .Y(n25288) );
  NAND2X1 U24737 ( .A(n457), .B(n73566), .Y(n25290) );
  NOR2X1 U24738 ( .A(n25291), .B(n25292), .Y(n25289) );
  NOR2X1 U24739 ( .A(n44296), .B(n1182), .Y(n25292) );
  NOR2X1 U24740 ( .A(n44293), .B(n1151), .Y(n25291) );
  NAND2X1 U24741 ( .A(n25293), .B(n25294), .Y(n25287) );
  NAND2X1 U24742 ( .A(u_csr_csr_sr_q_22), .B(n42144), .Y(n25294) );
  NOR2X1 U24743 ( .A(n25295), .B(n25296), .Y(n25293) );
  AND2X1 U24744 ( .A(cpu_id_i[22]), .B(n44289), .Y(n25296) );
  NOR2X1 U24745 ( .A(n44291), .B(n37697), .Y(n25295) );
  NOR2X1 U24746 ( .A(n25297), .B(n25298), .Y(n25285) );
  NAND2X1 U24747 ( .A(n25299), .B(n25300), .Y(n25298) );
  NAND2X1 U24749 ( .A(u_csr_csr_mtvec_q[22]), .B(n41738), .Y(n25299) );
  NAND2X1 U24750 ( .A(n25301), .B(n25302), .Y(n25297) );
  NAND2X1 U24751 ( .A(u_csr_csr_mscratch_q[22]), .B(n44080), .Y(n25302) );
  NOR2X1 U24752 ( .A(n25303), .B(n25304), .Y(n25301) );
  AND2X1 U24754 ( .A(n44079), .B(u_csr_csr_stval_q[22]), .Y(n25303) );
  NAND2X1 U24755 ( .A(n25305), .B(n25306), .Y(u_csr_result_r[21]) );
  NOR2X1 U24756 ( .A(n25307), .B(n25308), .Y(n25306) );
  NAND2X1 U24757 ( .A(n25309), .B(n25310), .Y(n25308) );
  NAND2X1 U24758 ( .A(n457), .B(n73567), .Y(n25310) );
  NOR2X1 U24759 ( .A(n25311), .B(n25312), .Y(n25309) );
  NOR2X1 U24760 ( .A(n44295), .B(n1183), .Y(n25312) );
  NOR2X1 U24761 ( .A(n44293), .B(n1152), .Y(n25311) );
  NAND2X1 U24762 ( .A(n25313), .B(n25314), .Y(n25307) );
  NAND2X1 U24763 ( .A(u_csr_csr_sr_q_21), .B(n44286), .Y(n25314) );
  NOR2X1 U24764 ( .A(n25315), .B(n25316), .Y(n25313) );
  AND2X1 U24765 ( .A(cpu_id_i[21]), .B(n44289), .Y(n25316) );
  NOR2X1 U24766 ( .A(n44291), .B(n37690), .Y(n25315) );
  NOR2X1 U24767 ( .A(n25317), .B(n25318), .Y(n25305) );
  NAND2X1 U24768 ( .A(n25319), .B(n25320), .Y(n25318) );
  NAND2X1 U24770 ( .A(u_csr_csr_mtvec_q[21]), .B(n41738), .Y(n25319) );
  NAND2X1 U24771 ( .A(n25321), .B(n25322), .Y(n25317) );
  NAND2X1 U24772 ( .A(u_csr_csr_mscratch_q[21]), .B(n44080), .Y(n25322) );
  NOR2X1 U24773 ( .A(n25323), .B(n42570), .Y(n25321) );
  AND2X1 U24775 ( .A(n44079), .B(u_csr_csr_stval_q[21]), .Y(n25323) );
  NAND2X1 U24776 ( .A(n25325), .B(n25326), .Y(u_csr_result_r[20]) );
  NOR2X1 U24777 ( .A(n25327), .B(n25328), .Y(n25326) );
  NAND2X1 U24778 ( .A(n25329), .B(n25330), .Y(n25328) );
  NAND2X1 U24779 ( .A(u_csr_csr_stvec_q[20]), .B(n36765), .Y(n25330) );
  NOR2X1 U24780 ( .A(n25331), .B(n25332), .Y(n25329) );
  NOR2X1 U24781 ( .A(n44293), .B(n1153), .Y(n25332) );
  AND2X1 U24782 ( .A(n44286), .B(u_csr_csr_sr_q_20), .Y(n25331) );
  NAND2X1 U24783 ( .A(n25333), .B(n25334), .Y(n25327) );
  NAND2X1 U24784 ( .A(cpu_id_i[20]), .B(n44288), .Y(n25334) );
  NOR2X1 U24785 ( .A(n24910), .B(n25335), .Y(n25333) );
  NOR2X1 U24786 ( .A(n44291), .B(n37585), .Y(n25335) );
  NOR2X1 U24787 ( .A(n25336), .B(n25337), .Y(n25325) );
  NAND2X1 U24788 ( .A(n25338), .B(n25339), .Y(n25337) );
  NAND2X1 U24789 ( .A(u_csr_csr_mtvec_q[20]), .B(n41738), .Y(n25339) );
  NOR2X1 U24790 ( .A(n25340), .B(n42565), .Y(n25338) );
  AND2X1 U24792 ( .A(n42849), .B(u_csr_csr_mscratch_q[20]), .Y(n25340) );
  NAND2X1 U24793 ( .A(n25342), .B(n25343), .Y(n25336) );
  NOR2X1 U24795 ( .A(n25344), .B(n25345), .Y(n25342) );
  AND2X1 U24796 ( .A(n44079), .B(u_csr_csr_stval_q[20]), .Y(n25345) );
  NOR2X1 U24797 ( .A(n1913), .B(n40682), .Y(n25344) );
  NAND2X1 U24798 ( .A(n25346), .B(n25347), .Y(u_csr_result_r[1]) );
  NOR2X1 U24799 ( .A(n25348), .B(n25349), .Y(n25347) );
  NAND2X1 U24800 ( .A(n25350), .B(n25351), .Y(n25349) );
  NAND2X1 U24801 ( .A(n457), .B(n73417), .Y(n25351) );
  NOR2X1 U24802 ( .A(n25352), .B(n25353), .Y(n25350) );
  NOR2X1 U24803 ( .A(n44295), .B(n37722), .Y(n25353) );
  NOR2X1 U24804 ( .A(n44293), .B(n1154), .Y(n25352) );
  NAND2X1 U24805 ( .A(n25354), .B(n25355), .Y(n25348) );
  NOR2X1 U24806 ( .A(n25356), .B(n25357), .Y(n25355) );
  NOR2X1 U24807 ( .A(n44290), .B(n37343), .Y(n25357) );
  NOR2X1 U24808 ( .A(n25358), .B(n24877), .Y(n25356) );
  NOR2X1 U24809 ( .A(n25359), .B(n25360), .Y(n25358) );
  NAND2X1 U24810 ( .A(n25361), .B(n25362), .Y(n25360) );
  NAND2X1 U24811 ( .A(u_csr_csr_mie_q_1), .B(n73402), .Y(n25362) );
  NAND2X1 U24813 ( .A(n25364), .B(n25365), .Y(n25359) );
  NAND2X1 U24814 ( .A(u_csr_csr_mip_q_1), .B(n73403), .Y(n25365) );
  AND2X1 U24816 ( .A(n25367), .B(n25368), .Y(n25354) );
  NAND2X1 U24817 ( .A(cpu_id_i[1]), .B(n44288), .Y(n25368) );
  NAND2X1 U24818 ( .A(u_csr_csr_sr_q[1]), .B(n458), .Y(n25367) );
  NOR2X1 U24819 ( .A(n25369), .B(n25370), .Y(n25346) );
  NAND2X1 U24820 ( .A(n25371), .B(n25372), .Y(n25370) );
  NAND2X1 U24821 ( .A(n42205), .B(u_csr_csr_mideleg_q[1]), .Y(n25372) );
  NOR2X1 U24822 ( .A(n25373), .B(n25374), .Y(n25371) );
  NOR2X1 U24823 ( .A(n42983), .B(n37713), .Y(n25374) );
  NAND2X1 U24825 ( .A(n25375), .B(n25376), .Y(n25369) );
  NOR2X1 U24826 ( .A(n25377), .B(n25378), .Y(n25376) );
  AND2X1 U24828 ( .A(n44079), .B(u_csr_csr_stval_q[1]), .Y(n25377) );
  NOR2X1 U24829 ( .A(n25379), .B(n25380), .Y(n25375) );
  AND2X1 U24830 ( .A(n73399), .B(u_csr_csr_medeleg_q[1]), .Y(n25380) );
  AND2X1 U24831 ( .A(n42848), .B(u_csr_csr_mscratch_q[1]), .Y(n25379) );
  NAND2X1 U24832 ( .A(n25381), .B(n25382), .Y(u_csr_result_r[19]) );
  NOR2X1 U24833 ( .A(n25383), .B(n25384), .Y(n25382) );
  NAND2X1 U24834 ( .A(n25385), .B(n25386), .Y(n25384) );
  NAND2X1 U24835 ( .A(n457), .B(n73408), .Y(n25386) );
  NOR2X1 U24836 ( .A(n25387), .B(n25388), .Y(n25385) );
  NOR2X1 U24837 ( .A(n44295), .B(n1186), .Y(n25388) );
  NOR2X1 U24838 ( .A(n44293), .B(n1155), .Y(n25387) );
  NAND2X1 U24839 ( .A(n25389), .B(n25390), .Y(n25383) );
  NAND2X1 U24840 ( .A(u_csr_csr_sr_q_19), .B(n44286), .Y(n25390) );
  NOR2X1 U24841 ( .A(n25391), .B(n25392), .Y(n25389) );
  AND2X1 U24842 ( .A(cpu_id_i[19]), .B(n44289), .Y(n25392) );
  NOR2X1 U24843 ( .A(n44290), .B(n37349), .Y(n25391) );
  NOR2X1 U24844 ( .A(n25393), .B(n25394), .Y(n25381) );
  NAND2X1 U24845 ( .A(n25395), .B(n25396), .Y(n25394) );
  NAND2X1 U24847 ( .A(u_csr_csr_mtvec_q[19]), .B(n41738), .Y(n25395) );
  NAND2X1 U24848 ( .A(n25397), .B(n25398), .Y(n25393) );
  NAND2X1 U24849 ( .A(u_csr_csr_mscratch_q[19]), .B(n44080), .Y(n25398) );
  NOR2X1 U24850 ( .A(n25399), .B(n42571), .Y(n25397) );
  AND2X1 U24852 ( .A(n44079), .B(u_csr_csr_stval_q[19]), .Y(n25399) );
  NAND2X1 U24853 ( .A(n25401), .B(n25402), .Y(u_csr_result_r[18]) );
  NOR2X1 U24854 ( .A(n25403), .B(n25404), .Y(n25402) );
  NAND2X1 U24855 ( .A(n25405), .B(n25406), .Y(n25404) );
  NAND2X1 U24856 ( .A(u_csr_csr_stvec_q[18]), .B(n36765), .Y(n25406) );
  NOR2X1 U24857 ( .A(n25407), .B(n25408), .Y(n25405) );
  NOR2X1 U24858 ( .A(n44293), .B(n1156), .Y(n25408) );
  NOR2X1 U24859 ( .A(n8835), .B(n25409), .Y(n25407) );
  NAND2X1 U24860 ( .A(n25410), .B(n25411), .Y(n25403) );
  NAND2X1 U24861 ( .A(cpu_id_i[18]), .B(n44288), .Y(n25411) );
  NOR2X1 U24862 ( .A(n24910), .B(n25412), .Y(n25410) );
  NOR2X1 U24863 ( .A(n44290), .B(n37696), .Y(n25412) );
  NOR2X1 U24864 ( .A(n25413), .B(n25414), .Y(n25401) );
  NAND2X1 U24865 ( .A(n25415), .B(n25416), .Y(n25414) );
  NAND2X1 U24866 ( .A(u_csr_csr_mtvec_q[18]), .B(n41738), .Y(n25416) );
  NOR2X1 U24867 ( .A(n25417), .B(n42566), .Y(n25415) );
  AND2X1 U24869 ( .A(n42849), .B(u_csr_csr_mscratch_q[18]), .Y(n25417) );
  NAND2X1 U24870 ( .A(n25419), .B(n25420), .Y(n25413) );
  NOR2X1 U24872 ( .A(n25421), .B(n25422), .Y(n25419) );
  AND2X1 U24873 ( .A(n44078), .B(u_csr_csr_stval_q[18]), .Y(n25422) );
  NOR2X1 U24874 ( .A(n1916), .B(n40681), .Y(n25421) );
  NAND2X1 U24875 ( .A(n25423), .B(n25424), .Y(u_csr_result_r[17]) );
  NOR2X1 U24876 ( .A(n25425), .B(n25426), .Y(n25424) );
  NAND2X1 U24877 ( .A(n25427), .B(n25428), .Y(n25426) );
  NAND2X1 U24878 ( .A(n457), .B(n73409), .Y(n25428) );
  NOR2X1 U24879 ( .A(n25429), .B(n25430), .Y(n25427) );
  NOR2X1 U24880 ( .A(n44295), .B(n1188), .Y(n25430) );
  NOR2X1 U24881 ( .A(n44293), .B(n1157), .Y(n25429) );
  NAND2X1 U24882 ( .A(n25431), .B(n25432), .Y(n25425) );
  NAND2X1 U24883 ( .A(u_csr_csr_sr_q[17]), .B(n44286), .Y(n25432) );
  NOR2X1 U24884 ( .A(n25433), .B(n25434), .Y(n25431) );
  AND2X1 U24885 ( .A(cpu_id_i[17]), .B(n44289), .Y(n25434) );
  NOR2X1 U24886 ( .A(n44290), .B(n37689), .Y(n25433) );
  NOR2X1 U24887 ( .A(n25435), .B(n25436), .Y(n25423) );
  NAND2X1 U24888 ( .A(n25437), .B(n25438), .Y(n25436) );
  NAND2X1 U24890 ( .A(u_csr_csr_mtvec_q[17]), .B(n41738), .Y(n25437) );
  NAND2X1 U24891 ( .A(n25439), .B(n25440), .Y(n25435) );
  NAND2X1 U24892 ( .A(u_csr_csr_mscratch_q[17]), .B(n44080), .Y(n25440) );
  NOR2X1 U24893 ( .A(n25441), .B(n42572), .Y(n25439) );
  AND2X1 U24895 ( .A(n44078), .B(u_csr_csr_stval_q[17]), .Y(n25441) );
  NAND2X1 U24896 ( .A(n25443), .B(n25444), .Y(u_csr_result_r[16]) );
  NOR2X1 U24897 ( .A(n25445), .B(n25446), .Y(n25444) );
  NAND2X1 U24898 ( .A(n25447), .B(n25448), .Y(n25446) );
  NAND2X1 U24899 ( .A(n457), .B(n73410), .Y(n25448) );
  NOR2X1 U24900 ( .A(n25449), .B(n25450), .Y(n25447) );
  NOR2X1 U24901 ( .A(n44295), .B(n1189), .Y(n25450) );
  NOR2X1 U24902 ( .A(n44294), .B(n1158), .Y(n25449) );
  NAND2X1 U24903 ( .A(n25451), .B(n25452), .Y(n25445) );
  NAND2X1 U24904 ( .A(u_csr_csr_sr_q[16]), .B(n44286), .Y(n25452) );
  NOR2X1 U24905 ( .A(n25453), .B(n25454), .Y(n25451) );
  AND2X1 U24906 ( .A(cpu_id_i[16]), .B(n44289), .Y(n25454) );
  NOR2X1 U24907 ( .A(n44290), .B(n37578), .Y(n25453) );
  NOR2X1 U24908 ( .A(n25455), .B(n25456), .Y(n25443) );
  NAND2X1 U24909 ( .A(n25457), .B(n25458), .Y(n25456) );
  NAND2X1 U24911 ( .A(u_csr_csr_mtvec_q[16]), .B(n41738), .Y(n25457) );
  NAND2X1 U24912 ( .A(n25459), .B(n25460), .Y(n25455) );
  NAND2X1 U24913 ( .A(u_csr_csr_mscratch_q[16]), .B(n44080), .Y(n25460) );
  NOR2X1 U24914 ( .A(n25461), .B(n42573), .Y(n25459) );
  AND2X1 U24916 ( .A(n44078), .B(u_csr_csr_stval_q[16]), .Y(n25461) );
  NAND2X1 U24917 ( .A(n25463), .B(n25464), .Y(u_csr_result_r[15]) );
  NOR2X1 U24918 ( .A(n25465), .B(n25466), .Y(n25464) );
  NAND2X1 U24919 ( .A(n25467), .B(n25468), .Y(n25466) );
  NAND2X1 U24920 ( .A(u_csr_csr_stval_q[15]), .B(n44078), .Y(n25468) );
  NOR2X1 U24921 ( .A(n25469), .B(n25470), .Y(n25467) );
  NOR2X1 U24922 ( .A(n1919), .B(n40682), .Y(n25470) );
  NOR2X1 U24923 ( .A(n44295), .B(n1190), .Y(n25469) );
  NAND2X1 U24924 ( .A(n25471), .B(n25472), .Y(n25465) );
  NOR2X1 U24925 ( .A(n25473), .B(n25474), .Y(n25472) );
  AND2X1 U24926 ( .A(cpu_id_i[15]), .B(n44289), .Y(n25474) );
  NOR2X1 U24927 ( .A(n44290), .B(n37348), .Y(n25473) );
  NOR2X1 U24928 ( .A(n25475), .B(n25476), .Y(n25471) );
  NOR2X1 U24929 ( .A(n44294), .B(n1159), .Y(n25476) );
  AND2X1 U24930 ( .A(n44286), .B(u_csr_csr_sr_q[15]), .Y(n25475) );
  NOR2X1 U24931 ( .A(n25477), .B(n25478), .Y(n25463) );
  NAND2X1 U24932 ( .A(n25479), .B(n25480), .Y(n25478) );
  NAND2X1 U24933 ( .A(u_csr_csr_mideleg_q[15]), .B(n42205), .Y(n25480) );
  NOR2X1 U24934 ( .A(n73497), .B(n25482), .Y(n25479) );
  NOR2X1 U24935 ( .A(n42982), .B(n37719), .Y(n25482) );
  NAND2X1 U24937 ( .A(n25483), .B(n25484), .Y(n25477) );
  NAND2X1 U24938 ( .A(u_csr_csr_medeleg_q[15]), .B(n73399), .Y(n25484) );
  NOR2X1 U24939 ( .A(n73496), .B(n25486), .Y(n25483) );
  AND2X1 U24940 ( .A(n42848), .B(u_csr_csr_mscratch_q[15]), .Y(n25486) );
  NAND2X1 U24942 ( .A(n25487), .B(n25488), .Y(u_csr_result_r[14]) );
  NOR2X1 U24943 ( .A(n25489), .B(n25490), .Y(n25488) );
  NAND2X1 U24944 ( .A(n25491), .B(n25492), .Y(n25490) );
  NAND2X1 U24945 ( .A(u_csr_csr_stval_q[14]), .B(n44078), .Y(n25492) );
  NOR2X1 U24946 ( .A(n25493), .B(n25494), .Y(n25491) );
  NOR2X1 U24947 ( .A(n1920), .B(n40681), .Y(n25494) );
  NOR2X1 U24948 ( .A(n44295), .B(n1191), .Y(n25493) );
  NAND2X1 U24949 ( .A(n25495), .B(n25496), .Y(n25489) );
  NOR2X1 U24950 ( .A(n25497), .B(n25498), .Y(n25496) );
  AND2X1 U24951 ( .A(cpu_id_i[14]), .B(n44288), .Y(n25498) );
  NOR2X1 U24952 ( .A(n44290), .B(n37712), .Y(n25497) );
  NOR2X1 U24953 ( .A(n25499), .B(n25500), .Y(n25495) );
  NOR2X1 U24954 ( .A(n44294), .B(n1160), .Y(n25500) );
  AND2X1 U24955 ( .A(n44286), .B(u_csr_csr_sr_q[14]), .Y(n25499) );
  NOR2X1 U24956 ( .A(n25501), .B(n25502), .Y(n25487) );
  NAND2X1 U24957 ( .A(n25503), .B(n25504), .Y(n25502) );
  NAND2X1 U24958 ( .A(u_csr_csr_mideleg_q[14]), .B(n42205), .Y(n25504) );
  NOR2X1 U24959 ( .A(n73499), .B(n25506), .Y(n25503) );
  NOR2X1 U24960 ( .A(n42982), .B(n37718), .Y(n25506) );
  NAND2X1 U24962 ( .A(n25507), .B(n25508), .Y(n25501) );
  NAND2X1 U24963 ( .A(u_csr_csr_medeleg_q[14]), .B(n73399), .Y(n25508) );
  NOR2X1 U24964 ( .A(n73498), .B(n25510), .Y(n25507) );
  AND2X1 U24965 ( .A(n42849), .B(u_csr_csr_mscratch_q[14]), .Y(n25510) );
  NAND2X1 U24967 ( .A(n25511), .B(n25512), .Y(u_csr_result_r[13]) );
  NOR2X1 U24968 ( .A(n25513), .B(n25514), .Y(n25512) );
  NAND2X1 U24969 ( .A(n25515), .B(n25516), .Y(n25514) );
  NAND2X1 U24970 ( .A(u_csr_csr_stval_q[13]), .B(n44078), .Y(n25516) );
  NOR2X1 U24971 ( .A(n25517), .B(n25518), .Y(n25515) );
  NOR2X1 U24972 ( .A(n1921), .B(n40682), .Y(n25518) );
  NOR2X1 U24973 ( .A(n44295), .B(n1192), .Y(n25517) );
  NAND2X1 U24974 ( .A(n25519), .B(n25520), .Y(n25513) );
  NOR2X1 U24975 ( .A(n25521), .B(n25522), .Y(n25520) );
  AND2X1 U24976 ( .A(cpu_id_i[13]), .B(n44289), .Y(n25522) );
  NOR2X1 U24977 ( .A(n44290), .B(n37692), .Y(n25521) );
  NOR2X1 U24978 ( .A(n25523), .B(n25524), .Y(n25519) );
  NOR2X1 U24979 ( .A(n44294), .B(n1161), .Y(n25524) );
  AND2X1 U24980 ( .A(n44286), .B(u_csr_csr_sr_q[13]), .Y(n25523) );
  NOR2X1 U24981 ( .A(n25525), .B(n25526), .Y(n25511) );
  NAND2X1 U24982 ( .A(n25527), .B(n25528), .Y(n25526) );
  NAND2X1 U24983 ( .A(u_csr_csr_mideleg_q[13]), .B(n42205), .Y(n25528) );
  NOR2X1 U24984 ( .A(n42564), .B(n25530), .Y(n25527) );
  NOR2X1 U24985 ( .A(n42983), .B(n37717), .Y(n25530) );
  NAND2X1 U24987 ( .A(n25531), .B(n25532), .Y(n25525) );
  NAND2X1 U24988 ( .A(u_csr_csr_medeleg_q[13]), .B(n73399), .Y(n25532) );
  NOR2X1 U24989 ( .A(n42569), .B(n25534), .Y(n25531) );
  AND2X1 U24990 ( .A(n42848), .B(u_csr_csr_mscratch_q[13]), .Y(n25534) );
  NAND2X1 U24992 ( .A(n25535), .B(n25536), .Y(u_csr_result_r[12]) );
  NOR2X1 U24993 ( .A(n25537), .B(n25538), .Y(n25536) );
  NAND2X1 U24994 ( .A(n25539), .B(n25540), .Y(n25538) );
  NAND2X1 U24995 ( .A(n457), .B(n73411), .Y(n25540) );
  NOR2X1 U24996 ( .A(n25541), .B(n25542), .Y(n25539) );
  NOR2X1 U24997 ( .A(n44295), .B(n1193), .Y(n25542) );
  NOR2X1 U24998 ( .A(n44294), .B(n1162), .Y(n25541) );
  NAND2X1 U24999 ( .A(n25543), .B(n25544), .Y(n25537) );
  NOR2X1 U25000 ( .A(n24910), .B(n25545), .Y(n25544) );
  NOR2X1 U25001 ( .A(n44290), .B(n37574), .Y(n25545) );
  AND2X1 U25004 ( .A(n25548), .B(n25549), .Y(n25543) );
  NAND2X1 U25005 ( .A(cpu_id_i[12]), .B(n44288), .Y(n25549) );
  NAND2X1 U25006 ( .A(u_csr_csr_sr_q[12]), .B(n44286), .Y(n25548) );
  NOR2X1 U25007 ( .A(n25550), .B(n25551), .Y(n25535) );
  NAND2X1 U25008 ( .A(n25552), .B(n25553), .Y(n25551) );
  NAND2X1 U25009 ( .A(u_csr_csr_mideleg_q[12]), .B(n42205), .Y(n25553) );
  NOR2X1 U25010 ( .A(n73502), .B(n25555), .Y(n25552) );
  NOR2X1 U25011 ( .A(n42982), .B(n37720), .Y(n25555) );
  NAND2X1 U25013 ( .A(n25556), .B(n25557), .Y(n25550) );
  NOR2X1 U25014 ( .A(n25558), .B(n73500), .Y(n25557) );
  AND2X1 U25016 ( .A(n44078), .B(u_csr_csr_stval_q[12]), .Y(n25558) );
  NOR2X1 U25017 ( .A(n25560), .B(n25561), .Y(n25556) );
  AND2X1 U25018 ( .A(n73399), .B(u_csr_csr_medeleg_q[12]), .Y(n25561) );
  AND2X1 U25019 ( .A(n44081), .B(u_csr_csr_mscratch_q[12]), .Y(n25560) );
  NAND2X1 U25020 ( .A(n25562), .B(n25563), .Y(u_csr_result_r[11]) );
  NOR2X1 U25021 ( .A(n25564), .B(n25565), .Y(n25563) );
  NAND2X1 U25022 ( .A(n25566), .B(n25567), .Y(n25565) );
  NAND2X1 U25023 ( .A(n457), .B(n73412), .Y(n25567) );
  NOR2X1 U25024 ( .A(n25568), .B(n25569), .Y(n25566) );
  NOR2X1 U25025 ( .A(n44295), .B(n1225), .Y(n25569) );
  NOR2X1 U25026 ( .A(n44294), .B(n1224), .Y(n25568) );
  NAND2X1 U25027 ( .A(n25570), .B(n25571), .Y(n25564) );
  NOR2X1 U25028 ( .A(n25572), .B(n25573), .Y(n25571) );
  NOR2X1 U25029 ( .A(n44290), .B(n37347), .Y(n25573) );
  NOR2X1 U25031 ( .A(n25575), .B(n25576), .Y(n25574) );
  NOR2X1 U25032 ( .A(n37485), .B(n24942), .Y(n25576) );
  NOR2X1 U25033 ( .A(n37553), .B(n24943), .Y(n25575) );
  AND2X1 U25034 ( .A(n25577), .B(n25578), .Y(n25570) );
  NAND2X1 U25035 ( .A(cpu_id_i[11]), .B(n44288), .Y(n25578) );
  NAND2X1 U25036 ( .A(u_csr_csr_sr_q[11]), .B(n44286), .Y(n25577) );
  NOR2X1 U25037 ( .A(n25579), .B(n25580), .Y(n25562) );
  NAND2X1 U25038 ( .A(n25581), .B(n25582), .Y(n25580) );
  NAND2X1 U25039 ( .A(u_csr_csr_mideleg_q[11]), .B(n42205), .Y(n25582) );
  NOR2X1 U25040 ( .A(n25583), .B(n25584), .Y(n25581) );
  NOR2X1 U25041 ( .A(n42982), .B(n37708), .Y(n25584) );
  NAND2X1 U25043 ( .A(n25585), .B(n25586), .Y(n25579) );
  NOR2X1 U25044 ( .A(n25587), .B(n25588), .Y(n25586) );
  AND2X1 U25046 ( .A(n44078), .B(u_csr_csr_stval_q[11]), .Y(n25587) );
  NOR2X1 U25047 ( .A(n25589), .B(n25590), .Y(n25585) );
  AND2X1 U25048 ( .A(n73399), .B(u_csr_csr_medeleg_q[11]), .Y(n25590) );
  AND2X1 U25049 ( .A(n44081), .B(u_csr_csr_mscratch_q[11]), .Y(n25589) );
  NAND2X1 U25050 ( .A(n25591), .B(n25592), .Y(u_csr_result_r[10]) );
  NOR2X1 U25051 ( .A(n25593), .B(n25594), .Y(n25592) );
  NAND2X1 U25052 ( .A(n25595), .B(n25596), .Y(n25594) );
  NAND2X1 U25053 ( .A(u_csr_csr_stval_q[10]), .B(n44078), .Y(n25596) );
  NOR2X1 U25054 ( .A(n25597), .B(n25598), .Y(n25595) );
  NOR2X1 U25055 ( .A(n1924), .B(n40681), .Y(n25598) );
  NOR2X1 U25056 ( .A(n44295), .B(n1194), .Y(n25597) );
  NAND2X1 U25057 ( .A(n25599), .B(n25600), .Y(n25593) );
  NOR2X1 U25058 ( .A(n25601), .B(n25602), .Y(n25600) );
  AND2X1 U25059 ( .A(cpu_id_i[10]), .B(n44288), .Y(n25602) );
  NOR2X1 U25060 ( .A(n44290), .B(n37711), .Y(n25601) );
  NOR2X1 U25061 ( .A(n25603), .B(n25604), .Y(n25599) );
  NOR2X1 U25062 ( .A(n44294), .B(n1163), .Y(n25604) );
  AND2X1 U25063 ( .A(n44286), .B(u_csr_csr_sr_q[10]), .Y(n25603) );
  NOR2X1 U25064 ( .A(n25605), .B(n25606), .Y(n25591) );
  NAND2X1 U25065 ( .A(n25607), .B(n25608), .Y(n25606) );
  NAND2X1 U25066 ( .A(u_csr_csr_mideleg_q[10]), .B(n42205), .Y(n25608) );
  NOR2X1 U25067 ( .A(n25609), .B(n25610), .Y(n25607) );
  NOR2X1 U25068 ( .A(n42983), .B(n37704), .Y(n25610) );
  NAND2X1 U25070 ( .A(n25611), .B(n25612), .Y(n25605) );
  NAND2X1 U25071 ( .A(u_csr_csr_medeleg_q[10]), .B(n73399), .Y(n25612) );
  NOR2X1 U25072 ( .A(n25613), .B(n25614), .Y(n25611) );
  AND2X1 U25073 ( .A(n44081), .B(u_csr_csr_mscratch_q[10]), .Y(n25614) );
  NAND2X1 U25075 ( .A(n25615), .B(n25616), .Y(u_csr_result_r[0]) );
  NOR2X1 U25076 ( .A(n25617), .B(n25618), .Y(n25616) );
  NAND2X1 U25077 ( .A(n25619), .B(n25620), .Y(n25618) );
  NOR2X1 U25078 ( .A(n25621), .B(n25622), .Y(n25620) );
  NOR2X1 U25079 ( .A(n44294), .B(n1164), .Y(n25622) );
  AND2X1 U25080 ( .A(n458), .B(u_csr_csr_sr_q[0]), .Y(n25621) );
  NOR2X1 U25081 ( .A(n25623), .B(n25624), .Y(n25619) );
  NOR2X1 U25082 ( .A(n1925), .B(n40682), .Y(n25624) );
  NOR2X1 U25083 ( .A(n44295), .B(n37702), .Y(n25623) );
  NAND2X1 U25084 ( .A(n25625), .B(n25626), .Y(n25617) );
  NOR2X1 U25085 ( .A(n25627), .B(n25628), .Y(n25626) );
  AND2X1 U25086 ( .A(n42145), .B(u_csr_csr_mcause_q[0]), .Y(n25628) );
  NOR2X1 U25087 ( .A(n25083), .B(n37727), .Y(n25627) );
  NOR2X1 U25088 ( .A(n25629), .B(n25630), .Y(n25625) );
  AND2X1 U25089 ( .A(cpu_id_i[0]), .B(n44289), .Y(n25630) );
  NOR2X1 U25097 ( .A(n44290), .B(n8886), .Y(n25629) );
  NOR2X1 U25099 ( .A(n25639), .B(n25640), .Y(n25638) );
  NOR2X1 U25105 ( .A(n25643), .B(n25644), .Y(n25615) );
  NAND2X1 U25106 ( .A(n25645), .B(n25646), .Y(n25644) );
  NAND2X1 U25107 ( .A(u_csr_csr_mideleg_q[0]), .B(n42205), .Y(n25646) );
  NOR2X1 U25108 ( .A(n25647), .B(n25648), .Y(n25645) );
  NOR2X1 U25109 ( .A(n42982), .B(n37707), .Y(n25648) );
  NAND2X1 U25111 ( .A(n25649), .B(n25650), .Y(n25643) );
  NOR2X1 U25112 ( .A(n25651), .B(n25652), .Y(n25650) );
  AND2X1 U25114 ( .A(n44079), .B(u_csr_csr_stval_q[0]), .Y(n25651) );
  NOR2X1 U25115 ( .A(n25653), .B(n25654), .Y(n25649) );
  AND2X1 U25116 ( .A(n73399), .B(u_csr_csr_medeleg_q[0]), .Y(n25654) );
  AND2X1 U25117 ( .A(n42848), .B(u_csr_csr_mscratch_q[0]), .Y(n25653) );
  NAND2X1 U25139 ( .A(n25677), .B(n25678), .Y(u_csr_csr_stvec_r[4]) );
  NAND2X1 U25140 ( .A(u_csr_csr_stvec_q[4]), .B(n25679), .Y(n25678) );
  NAND2X1 U25141 ( .A(n25680), .B(n25681), .Y(n25679) );
  NAND2X1 U25143 ( .A(n25683), .B(n25684), .Y(u_csr_csr_stvec_r[3]) );
  NAND2X1 U25144 ( .A(u_csr_csr_stvec_q[3]), .B(n25685), .Y(n25684) );
  NAND2X1 U25145 ( .A(n25680), .B(n25686), .Y(n25685) );
  NAND2X1 U25155 ( .A(n25696), .B(n25697), .Y(u_csr_csr_stvec_r[2]) );
  NAND2X1 U25156 ( .A(u_csr_csr_stvec_q[2]), .B(n25698), .Y(n25697) );
  NAND2X1 U25157 ( .A(n25680), .B(n25699), .Y(n25698) );
  NAND2X1 U25199 ( .A(n25741), .B(n25742), .Y(u_csr_csr_stvec_r[1]) );
  NAND2X1 U25200 ( .A(u_csr_csr_stvec_q[1]), .B(n25743), .Y(n25742) );
  NAND2X1 U25201 ( .A(n25680), .B(n25744), .Y(n25743) );
  NAND2X1 U25245 ( .A(n25788), .B(n25789), .Y(u_csr_csr_stvec_r[0]) );
  NAND2X1 U25246 ( .A(u_csr_csr_stvec_q[0]), .B(n25790), .Y(n25789) );
  NAND2X1 U25247 ( .A(n25680), .B(n25791), .Y(n25790) );
  NOR2X1 U25248 ( .A(n25792), .B(n42302), .Y(n25680) );
  NAND2X1 U25250 ( .A(n25795), .B(n25796), .Y(u_csr_csr_stval_r[9]) );
  NOR2X1 U25251 ( .A(n25797), .B(n25798), .Y(n25796) );
  NOR2X1 U25258 ( .A(n25807), .B(n25808), .Y(n25795) );
  NAND2X1 U25261 ( .A(n25811), .B(n25812), .Y(u_csr_csr_stval_r[8]) );
  NOR2X1 U25262 ( .A(n25813), .B(n25814), .Y(n25812) );
  NOR2X1 U25269 ( .A(n25819), .B(n25820), .Y(n25811) );
  NAND2X1 U25272 ( .A(n25821), .B(n25822), .Y(u_csr_csr_stval_r[7]) );
  NOR2X1 U25273 ( .A(n25823), .B(n25824), .Y(n25822) );
  NOR2X1 U25280 ( .A(n25829), .B(n25830), .Y(n25821) );
  NAND2X1 U25283 ( .A(n25831), .B(n25832), .Y(u_csr_csr_stval_r[6]) );
  NOR2X1 U25284 ( .A(n25833), .B(n25834), .Y(n25832) );
  NOR2X1 U25291 ( .A(n25839), .B(n25840), .Y(n25831) );
  NAND2X1 U25294 ( .A(n25841), .B(n25842), .Y(u_csr_csr_stval_r[5]) );
  NOR2X1 U25295 ( .A(n25843), .B(n25844), .Y(n25842) );
  NOR2X1 U25302 ( .A(n25849), .B(n25850), .Y(n25841) );
  NAND2X1 U25305 ( .A(n25851), .B(n25852), .Y(u_csr_csr_stval_r[4]) );
  NOR2X1 U25306 ( .A(n25853), .B(n25854), .Y(n25852) );
  NAND2X1 U25307 ( .A(n25855), .B(n25856), .Y(n25854) );
  NAND2X1 U25308 ( .A(u_csr_csr_stval_q[4]), .B(n25857), .Y(n25856) );
  NAND2X1 U25309 ( .A(n25858), .B(n25859), .Y(n25857) );
  NAND2X1 U25310 ( .A(n42210), .B(n25860), .Y(n25859) );
  NOR2X1 U25313 ( .A(n25861), .B(n25862), .Y(n25851) );
  NAND2X1 U25316 ( .A(n25864), .B(n25865), .Y(u_csr_csr_stval_r[3]) );
  NOR2X1 U25317 ( .A(n25866), .B(n25867), .Y(n25865) );
  NAND2X1 U25318 ( .A(n25868), .B(n25869), .Y(n25867) );
  NAND2X1 U25319 ( .A(u_csr_csr_stval_q[3]), .B(n25870), .Y(n25869) );
  NAND2X1 U25320 ( .A(n25858), .B(n25871), .Y(n25870) );
  NAND2X1 U25321 ( .A(n42210), .B(n25872), .Y(n25871) );
  NOR2X1 U25324 ( .A(n25873), .B(n25874), .Y(n25864) );
  NAND2X1 U25327 ( .A(n25875), .B(n25876), .Y(u_csr_csr_stval_r[31]) );
  NOR2X1 U25328 ( .A(n25877), .B(n25878), .Y(n25876) );
  NAND2X1 U25338 ( .A(n25885), .B(n25886), .Y(u_csr_csr_stval_r[30]) );
  NOR2X1 U25339 ( .A(n25887), .B(n25888), .Y(n25886) );
  NAND2X1 U25349 ( .A(n25895), .B(n25896), .Y(u_csr_csr_stval_r[2]) );
  NOR2X1 U25350 ( .A(n25897), .B(n25898), .Y(n25896) );
  NAND2X1 U25351 ( .A(n25899), .B(n25900), .Y(n25898) );
  NAND2X1 U25352 ( .A(u_csr_csr_stval_q[2]), .B(n25901), .Y(n25900) );
  NAND2X1 U25353 ( .A(n25858), .B(n25902), .Y(n25901) );
  NAND2X1 U25354 ( .A(n42210), .B(n25903), .Y(n25902) );
  NOR2X1 U25357 ( .A(n25904), .B(n25905), .Y(n25895) );
  NAND2X1 U25360 ( .A(n25906), .B(n25907), .Y(u_csr_csr_stval_r[29]) );
  NOR2X1 U25361 ( .A(n25908), .B(n25909), .Y(n25907) );
  NOR2X1 U25368 ( .A(n25914), .B(n25915), .Y(n25906) );
  NAND2X1 U25371 ( .A(n25916), .B(n25917), .Y(u_csr_csr_stval_r[28]) );
  NOR2X1 U25372 ( .A(n25918), .B(n25919), .Y(n25917) );
  NAND2X1 U25382 ( .A(n25926), .B(n25927), .Y(u_csr_csr_stval_r[27]) );
  NOR2X1 U25383 ( .A(n25928), .B(n25929), .Y(n25927) );
  NAND2X1 U25393 ( .A(n25936), .B(n25937), .Y(u_csr_csr_stval_r[26]) );
  NOR2X1 U25394 ( .A(n25938), .B(n25939), .Y(n25937) );
  NAND2X1 U25404 ( .A(n25946), .B(n25947), .Y(u_csr_csr_stval_r[25]) );
  NOR2X1 U25405 ( .A(n25948), .B(n25949), .Y(n25947) );
  NOR2X1 U25412 ( .A(n25954), .B(n25955), .Y(n25946) );
  NAND2X1 U25415 ( .A(n25956), .B(n25957), .Y(u_csr_csr_stval_r[24]) );
  NOR2X1 U25416 ( .A(n25958), .B(n25959), .Y(n25957) );
  NAND2X1 U25426 ( .A(n25966), .B(n25967), .Y(u_csr_csr_stval_r[23]) );
  NOR2X1 U25427 ( .A(n25968), .B(n25969), .Y(n25967) );
  NAND2X1 U25437 ( .A(n25976), .B(n25977), .Y(u_csr_csr_stval_r[22]) );
  NOR2X1 U25438 ( .A(n25978), .B(n25979), .Y(n25977) );
  NAND2X1 U25448 ( .A(n25986), .B(n25987), .Y(u_csr_csr_stval_r[21]) );
  NOR2X1 U25449 ( .A(n25988), .B(n25989), .Y(n25987) );
  NAND2X1 U25459 ( .A(n25996), .B(n25997), .Y(u_csr_csr_stval_r[20]) );
  NOR2X1 U25460 ( .A(n25998), .B(n25999), .Y(n25997) );
  NOR2X1 U25467 ( .A(n26004), .B(n26005), .Y(n25996) );
  NAND2X1 U25470 ( .A(n26006), .B(n26007), .Y(u_csr_csr_stval_r[1]) );
  NOR2X1 U25471 ( .A(n26008), .B(n26009), .Y(n26007) );
  NAND2X1 U25472 ( .A(n26010), .B(n26011), .Y(n26009) );
  NAND2X1 U25473 ( .A(u_csr_csr_stval_q[1]), .B(n26012), .Y(n26011) );
  NAND2X1 U25474 ( .A(n25858), .B(n26013), .Y(n26012) );
  NAND2X1 U25475 ( .A(n42210), .B(n26014), .Y(n26013) );
  NOR2X1 U25478 ( .A(n26015), .B(n26016), .Y(n26006) );
  NAND2X1 U25481 ( .A(n26017), .B(n26018), .Y(u_csr_csr_stval_r[19]) );
  NOR2X1 U25482 ( .A(n26019), .B(n26020), .Y(n26018) );
  NOR2X1 U25489 ( .A(n26025), .B(n26026), .Y(n26017) );
  NAND2X1 U25492 ( .A(n26027), .B(n26028), .Y(u_csr_csr_stval_r[18]) );
  NOR2X1 U25493 ( .A(n26029), .B(n26030), .Y(n26028) );
  NAND2X1 U25503 ( .A(n26037), .B(n26038), .Y(u_csr_csr_stval_r[17]) );
  NOR2X1 U25504 ( .A(n26039), .B(n26040), .Y(n26038) );
  NAND2X1 U25514 ( .A(n26047), .B(n26048), .Y(u_csr_csr_stval_r[16]) );
  NOR2X1 U25515 ( .A(n26049), .B(n26050), .Y(n26048) );
  NOR2X1 U25522 ( .A(n26055), .B(n26056), .Y(n26047) );
  NAND2X1 U25525 ( .A(n26057), .B(n26058), .Y(u_csr_csr_stval_r[15]) );
  NOR2X1 U25526 ( .A(n26059), .B(n26060), .Y(n26058) );
  NAND2X1 U25536 ( .A(n26067), .B(n26068), .Y(u_csr_csr_stval_r[14]) );
  NOR2X1 U25537 ( .A(n26069), .B(n26070), .Y(n26068) );
  NAND2X1 U25547 ( .A(n26077), .B(n26078), .Y(u_csr_csr_stval_r[13]) );
  NOR2X1 U25548 ( .A(n26079), .B(n26080), .Y(n26078) );
  NAND2X1 U25558 ( .A(n26087), .B(n26088), .Y(u_csr_csr_stval_r[12]) );
  NOR2X1 U25559 ( .A(n26089), .B(n26090), .Y(n26088) );
  NAND2X1 U25569 ( .A(n26097), .B(n26098), .Y(u_csr_csr_stval_r[11]) );
  NOR2X1 U25570 ( .A(n26099), .B(n26100), .Y(n26098) );
  NOR2X1 U25577 ( .A(n26105), .B(n26106), .Y(n26097) );
  NAND2X1 U25580 ( .A(n26107), .B(n26108), .Y(u_csr_csr_stval_r[10]) );
  NOR2X1 U25581 ( .A(n26109), .B(n26110), .Y(n26108) );
  NAND2X1 U25587 ( .A(n973), .B(n44078), .Y(n26116) );
  NOR2X1 U25591 ( .A(n26117), .B(n26118), .Y(n26107) );
  NAND2X1 U25594 ( .A(n26119), .B(n26120), .Y(u_csr_csr_stval_r[0]) );
  NOR2X1 U25595 ( .A(n26121), .B(n26122), .Y(n26120) );
  NAND2X1 U25596 ( .A(n26123), .B(n26124), .Y(n26122) );
  NAND2X1 U25597 ( .A(u_csr_csr_stval_q[0]), .B(n26125), .Y(n26124) );
  NAND2X1 U25598 ( .A(n25858), .B(n26126), .Y(n26125) );
  NAND2X1 U25599 ( .A(n42210), .B(n26127), .Y(n26126) );
  AND2X1 U25601 ( .A(n26115), .B(n26128), .Y(n25858) );
  NAND2X1 U25602 ( .A(n44078), .B(n26129), .Y(n26128) );
  AND2X1 U25603 ( .A(n26130), .B(n26131), .Y(n26115) );
  NOR2X1 U25604 ( .A(n73501), .B(n26132), .Y(n26131) );
  AND2X1 U25605 ( .A(n26133), .B(n42962), .Y(n26132) );
  NOR2X1 U25606 ( .A(n26134), .B(n26135), .Y(n26130) );
  NOR2X1 U25612 ( .A(n26139), .B(n26140), .Y(n26119) );
  NAND2X1 U25636 ( .A(n26159), .B(n26160), .Y(u_csr_csr_sscratch_r[4]) );
  NAND2X1 U25637 ( .A(u_csr_csr_sscratch_q[4]), .B(n26161), .Y(n26160) );
  NAND2X1 U25638 ( .A(n26162), .B(n25681), .Y(n26161) );
  NAND2X1 U25640 ( .A(n26164), .B(n26165), .Y(u_csr_csr_sscratch_r[3]) );
  NAND2X1 U25641 ( .A(u_csr_csr_sscratch_q[3]), .B(n26166), .Y(n26165) );
  NAND2X1 U25642 ( .A(n26162), .B(n25686), .Y(n26166) );
  NAND2X1 U25652 ( .A(n26173), .B(n26174), .Y(u_csr_csr_sscratch_r[2]) );
  NAND2X1 U25653 ( .A(u_csr_csr_sscratch_q[2]), .B(n26175), .Y(n26174) );
  NAND2X1 U25654 ( .A(n26162), .B(n25699), .Y(n26175) );
  NAND2X1 U25696 ( .A(n26206), .B(n26207), .Y(u_csr_csr_sscratch_r[1]) );
  NAND2X1 U25697 ( .A(u_csr_csr_sscratch_q[1]), .B(n26208), .Y(n26207) );
  NAND2X1 U25698 ( .A(n26162), .B(n25744), .Y(n26208) );
  NAND2X1 U25741 ( .A(n26241), .B(n26242), .Y(n25786) );
  NOR2X1 U25742 ( .A(n973), .B(n44081), .Y(n26241) );
  NAND2X1 U25745 ( .A(n26244), .B(n26245), .Y(u_csr_csr_sscratch_r[0]) );
  NAND2X1 U25746 ( .A(u_csr_csr_sscratch_q[0]), .B(n26246), .Y(n26245) );
  NAND2X1 U25747 ( .A(n26162), .B(n25791), .Y(n26246) );
  NAND2X1 U25751 ( .A(n26249), .B(n26242), .Y(n25792) );
  NOR2X1 U25752 ( .A(n26129), .B(n42849), .Y(n26249) );
  NAND2X1 U25754 ( .A(n26250), .B(n26251), .Y(u_csr_csr_sr_r_8) );
  NAND2X1 U25755 ( .A(u_csr_N3161), .B(n26252), .Y(n26251) );
  NOR2X1 U25756 ( .A(n26253), .B(n26254), .Y(n26250) );
  NOR2X1 U25757 ( .A(n26255), .B(n37663), .Y(n26254) );
  NOR2X1 U25758 ( .A(n26256), .B(n26257), .Y(n26255) );
  NAND2X1 U25762 ( .A(n26262), .B(n26263), .Y(u_csr_csr_sr_r_7) );
  NOR2X1 U25763 ( .A(n469), .B(n26264), .Y(n26263) );
  NOR2X1 U25764 ( .A(n26265), .B(n37750), .Y(n26264) );
  NOR2X1 U25765 ( .A(n26266), .B(n26267), .Y(n26265) );
  NAND2X1 U25766 ( .A(n26268), .B(n26269), .Y(n26267) );
  NAND2X1 U25771 ( .A(n26277), .B(n26278), .Y(u_csr_csr_sr_r_5) );
  NOR2X1 U25772 ( .A(n470), .B(n26279), .Y(n26278) );
  NOR2X1 U25773 ( .A(n26280), .B(n37751), .Y(n26279) );
  NOR2X1 U25774 ( .A(n26281), .B(n26282), .Y(n26280) );
  NAND2X1 U25775 ( .A(n26283), .B(n26258), .Y(n26282) );
  NOR2X1 U25777 ( .A(n26286), .B(n26287), .Y(n26277) );
  NOR2X1 U25778 ( .A(n73507), .B(n37540), .Y(n26287) );
  NAND2X1 U25780 ( .A(n26289), .B(n26290), .Y(u_csr_csr_sr_r_3) );
  NOR2X1 U25782 ( .A(n26291), .B(n26292), .Y(n26289) );
  NOR2X1 U25783 ( .A(n37750), .B(n26272), .Y(n26292) );
  NOR2X1 U25784 ( .A(n26293), .B(n37748), .Y(n26291) );
  NOR2X1 U25785 ( .A(n26294), .B(n26295), .Y(n26293) );
  NAND2X1 U25786 ( .A(n26296), .B(n26297), .Y(n26295) );
  NAND2X1 U25787 ( .A(n42144), .B(n26129), .Y(n26296) );
  NAND2X1 U25788 ( .A(n26298), .B(n26299), .Y(u_csr_csr_sr_r_12) );
  NAND2X1 U25789 ( .A(u_csr_N3162), .B(n58246), .Y(n26299) );
  NAND2X1 U25795 ( .A(n26306), .B(n26307), .Y(u_csr_csr_sr_r_11) );
  NAND2X1 U25796 ( .A(u_csr_N3161), .B(n58246), .Y(n26307) );
  NAND2X1 U25801 ( .A(n459), .B(n26269), .Y(n26304) );
  NAND2X1 U25802 ( .A(n973), .B(n42144), .Y(n26269) );
  NAND2X1 U25804 ( .A(n26312), .B(n26268), .Y(n26294) );
  AND2X1 U25805 ( .A(n26313), .B(n73507), .Y(n26268) );
  NOR2X1 U25806 ( .A(n461), .B(n26314), .Y(n26313) );
  NOR2X1 U25807 ( .A(n26315), .B(n42445), .Y(n26312) );
  NAND2X1 U25808 ( .A(n26318), .B(n26319), .Y(u_csr_csr_sr_r_1) );
  NAND2X1 U25809 ( .A(n73509), .B(n26261), .Y(n26319) );
  NOR2X1 U25810 ( .A(n26320), .B(n26321), .Y(n26318) );
  NOR2X1 U25811 ( .A(n37751), .B(n26285), .Y(n26321) );
  NAND2X1 U25812 ( .A(n42445), .B(n42607), .Y(n26285) );
  NOR2X1 U25814 ( .A(n26323), .B(n37540), .Y(n26320) );
  NOR2X1 U25815 ( .A(n411), .B(n26256), .Y(n26323) );
  NAND2X1 U25816 ( .A(n26324), .B(n26283), .Y(n26256) );
  NOR2X1 U25817 ( .A(n26325), .B(n26314), .Y(n26283) );
  NAND2X1 U25818 ( .A(n26326), .B(n26327), .Y(n26314) );
  NAND2X1 U25819 ( .A(n42962), .B(n26328), .Y(n26326) );
  OR2X1 U25820 ( .A(n26329), .B(n58246), .Y(n26325) );
  NOR2X1 U25821 ( .A(n73577), .B(n25409), .Y(n26329) );
  NAND2X1 U25822 ( .A(n42962), .B(n26261), .Y(n25409) );
  NOR2X1 U25823 ( .A(n26315), .B(n42581), .Y(n26324) );
  AND2X1 U25859 ( .A(n26360), .B(n26361), .Y(n26335) );
  NOR2X1 U25860 ( .A(n461), .B(n24877), .Y(n26360) );
  NAND2X1 U26177 ( .A(n26456), .B(n26331), .Y(n26714) );
  NAND2X1 U26312 ( .A(n973), .B(n73501), .Y(n26856) );
  AND2X1 U26343 ( .A(n26456), .B(n26258), .Y(n26373) );
  NAND2X1 U26357 ( .A(n26456), .B(n26906), .Y(n26905) );
  AND2X1 U26358 ( .A(n26855), .B(n26907), .Y(n26456) );
  NAND2X1 U26359 ( .A(n73501), .B(n26129), .Y(n26907) );
  NOR2X1 U26361 ( .A(n26908), .B(n26135), .Y(n26855) );
  NAND2X1 U26362 ( .A(n26909), .B(n26910), .Y(n26135) );
  NOR2X1 U26363 ( .A(n36765), .B(n26911), .Y(n26910) );
  NAND2X1 U26364 ( .A(n40681), .B(n26912), .Y(n26911) );
  NOR2X1 U26367 ( .A(n26913), .B(n26914), .Y(n26909) );
  NAND2X1 U26368 ( .A(n73514), .B(n44294), .Y(n26914) );
  OR2X1 U26371 ( .A(n44078), .B(n26916), .Y(n26908) );
  NOR2X1 U26372 ( .A(n26917), .B(n24877), .Y(n26916) );
  NAND2X1 U26392 ( .A(n26932), .B(n26933), .Y(u_csr_csr_scause_r_31) );
  NAND2X1 U26393 ( .A(u_csr_csr_scause_q_31), .B(n26934), .Y(n26933) );
  NAND2X1 U26394 ( .A(n26935), .B(n26936), .Y(n26934) );
  NOR2X1 U26395 ( .A(n73508), .B(n26937), .Y(n26932) );
  NAND2X1 U26398 ( .A(n26939), .B(n26940), .Y(u_csr_csr_scause_r[3]) );
  NOR2X1 U26399 ( .A(n26941), .B(n26942), .Y(n26940) );
  NAND2X1 U26400 ( .A(n26943), .B(n26944), .Y(n26942) );
  NAND2X1 U26401 ( .A(n42461), .B(n73517), .Y(n26944) );
  NAND2X1 U26402 ( .A(u_csr_csr_scause_q[3]), .B(n26946), .Y(n26943) );
  OR2X1 U26403 ( .A(n26947), .B(n375), .Y(n26946) );
  NOR2X1 U26405 ( .A(n26949), .B(n26950), .Y(n26939) );
  NOR2X1 U26406 ( .A(n1082), .B(n26928), .Y(n26950) );
  NAND2X1 U26408 ( .A(n26952), .B(n26953), .Y(u_csr_csr_scause_r[2]) );
  NOR2X1 U26409 ( .A(n26954), .B(n26955), .Y(n26953) );
  NOR2X1 U26413 ( .A(n26958), .B(n37728), .Y(n26954) );
  NOR2X1 U26414 ( .A(n391), .B(n26947), .Y(n26958) );
  NOR2X1 U26415 ( .A(n26960), .B(n26961), .Y(n26952) );
  NOR2X1 U26417 ( .A(n26962), .B(n26931), .Y(n26960) );
  NAND2X1 U26418 ( .A(n26963), .B(n26964), .Y(u_csr_csr_scause_r[1]) );
  NOR2X1 U26419 ( .A(n26965), .B(n26966), .Y(n26964) );
  NAND2X1 U26420 ( .A(n26967), .B(n26968), .Y(n26966) );
  NAND2X1 U26421 ( .A(n26969), .B(n73508), .Y(n26968) );
  NAND2X1 U26422 ( .A(n26970), .B(n73517), .Y(n26967) );
  AND2X1 U26423 ( .A(n26971), .B(n8810), .Y(n26970) );
  NOR2X1 U26424 ( .A(n26972), .B(n37762), .Y(n26965) );
  NOR2X1 U26425 ( .A(n410), .B(n26947), .Y(n26972) );
  NAND2X1 U26426 ( .A(n26973), .B(n26974), .Y(n26947) );
  NOR2X1 U26427 ( .A(n42145), .B(n466), .Y(n26974) );
  NOR2X1 U26429 ( .A(n26976), .B(n26977), .Y(n26973) );
  NOR2X1 U26430 ( .A(n26979), .B(n26980), .Y(n26963) );
  NAND2X1 U26433 ( .A(n26981), .B(n26982), .Y(u_csr_csr_scause_r[0]) );
  NOR2X1 U26434 ( .A(n26983), .B(n26984), .Y(n26982) );
  NAND2X1 U26435 ( .A(n26985), .B(n26928), .Y(n26984) );
  NAND2X1 U26436 ( .A(n26986), .B(n73517), .Y(n26985) );
  NOR2X1 U26438 ( .A(n26988), .B(n26951), .Y(n26983) );
  NOR2X1 U26440 ( .A(n26989), .B(n26990), .Y(n26981) );
  NOR2X1 U26442 ( .A(n26991), .B(n37727), .Y(n26989) );
  AND2X1 U26443 ( .A(n26992), .B(n26935), .Y(n26991) );
  AND2X1 U26444 ( .A(n26993), .B(n26994), .Y(n26935) );
  NOR2X1 U26445 ( .A(n73516), .B(n26995), .Y(n26994) );
  NOR2X1 U26447 ( .A(n26997), .B(n26998), .Y(n26993) );
  NOR2X1 U26448 ( .A(n73543), .B(n73574), .Y(n26997) );
  NAND2X1 U26471 ( .A(n27019), .B(n25681), .Y(n27018) );
  NAND2X1 U26475 ( .A(n27019), .B(n25686), .Y(n27022) );
  NAND2X1 U26487 ( .A(n27019), .B(n25699), .Y(n27031) );
  NAND2X1 U26531 ( .A(n27019), .B(n25744), .Y(n27064) );
  NAND2X1 U26577 ( .A(n27019), .B(n25791), .Y(n27100) );
  AND2X1 U26578 ( .A(n27095), .B(n73577), .Y(n27019) );
  AND2X1 U26579 ( .A(n27101), .B(n27102), .Y(n27095) );
  NOR2X1 U26580 ( .A(n44080), .B(n24877), .Y(n27102) );
  NOR2X1 U26582 ( .A(n27104), .B(n451), .Y(n27101) );
  NAND2X1 U26604 ( .A(n27122), .B(n27123), .Y(u_csr_csr_mtvec_r[4]) );
  NAND2X1 U26605 ( .A(u_csr_csr_mtvec_q[4]), .B(n27124), .Y(n27123) );
  NAND2X1 U26606 ( .A(n27125), .B(n25681), .Y(n27124) );
  NAND2X1 U26608 ( .A(n27126), .B(n27127), .Y(u_csr_csr_mtvec_r[3]) );
  NAND2X1 U26609 ( .A(u_csr_csr_mtvec_q[3]), .B(n27128), .Y(n27127) );
  NAND2X1 U26610 ( .A(n27125), .B(n25686), .Y(n27128) );
  NAND2X1 U26620 ( .A(n27135), .B(n27136), .Y(u_csr_csr_mtvec_r[2]) );
  NAND2X1 U26621 ( .A(u_csr_csr_mtvec_q[2]), .B(n27137), .Y(n27136) );
  NAND2X1 U26622 ( .A(n27125), .B(n25699), .Y(n27137) );
  NAND2X1 U26664 ( .A(n27168), .B(n27169), .Y(u_csr_csr_mtvec_r[1]) );
  NAND2X1 U26665 ( .A(u_csr_csr_mtvec_q[1]), .B(n27170), .Y(n27169) );
  NAND2X1 U26666 ( .A(n27125), .B(n25744), .Y(n27170) );
  AND2X1 U26708 ( .A(n27096), .B(n27203), .Y(n27201) );
  NAND2X1 U26711 ( .A(n27205), .B(n27206), .Y(u_csr_csr_mtvec_r[0]) );
  NAND2X1 U26712 ( .A(u_csr_csr_mtvec_q[0]), .B(n27207), .Y(n27206) );
  NAND2X1 U26713 ( .A(n27125), .B(n25791), .Y(n27207) );
  AND2X1 U26714 ( .A(n27208), .B(n27203), .Y(n27125) );
  NAND2X1 U26739 ( .A(n27226), .B(n27227), .Y(u_csr_csr_mscratch_r[4]) );
  NAND2X1 U26740 ( .A(u_csr_csr_mscratch_q[4]), .B(n27228), .Y(n27227) );
  NAND2X1 U26741 ( .A(n27229), .B(n25681), .Y(n27228) );
  NAND2X1 U26743 ( .A(n27230), .B(n27231), .Y(u_csr_csr_mscratch_r[3]) );
  NAND2X1 U26744 ( .A(u_csr_csr_mscratch_q[3]), .B(n27232), .Y(n27231) );
  NAND2X1 U26745 ( .A(n27229), .B(n25686), .Y(n27232) );
  NAND2X1 U26746 ( .A(n44082), .B(n25872), .Y(n25686) );
  NAND2X1 U26758 ( .A(n27239), .B(n27240), .Y(u_csr_csr_mscratch_r[2]) );
  NAND2X1 U26759 ( .A(u_csr_csr_mscratch_q[2]), .B(n27241), .Y(n27240) );
  NAND2X1 U26760 ( .A(n27229), .B(n25699), .Y(n27241) );
  NAND2X1 U26809 ( .A(n27272), .B(n27273), .Y(u_csr_csr_mscratch_r[1]) );
  NAND2X1 U26810 ( .A(u_csr_csr_mscratch_q[1]), .B(n27274), .Y(n27273) );
  NAND2X1 U26811 ( .A(n27229), .B(n25744), .Y(n27274) );
  NAND2X1 U26812 ( .A(n44082), .B(n26014), .Y(n25744) );
  NOR2X1 U26855 ( .A(n973), .B(n27104), .Y(n27305) );
  NAND2X1 U26858 ( .A(n27306), .B(n27307), .Y(u_csr_csr_mscratch_r[0]) );
  NAND2X1 U26859 ( .A(u_csr_csr_mscratch_q[0]), .B(n27308), .Y(n27307) );
  NAND2X1 U26860 ( .A(n27229), .B(n25791), .Y(n27308) );
  AND2X1 U26861 ( .A(n27309), .B(n26242), .Y(n27229) );
  AND2X1 U26862 ( .A(n27310), .B(n26917), .Y(n26242) );
  NOR2X1 U26863 ( .A(n26133), .B(n26134), .Y(n26917) );
  NAND2X1 U26864 ( .A(n27311), .B(n27203), .Y(n26134) );
  NOR2X1 U26865 ( .A(n41738), .B(n42131), .Y(n27311) );
  NOR2X1 U26866 ( .A(n73539), .B(n24877), .Y(n27310) );
  NOR2X1 U26867 ( .A(n26129), .B(n27104), .Y(n27309) );
  NAND2X1 U26869 ( .A(n27312), .B(n73514), .Y(n36340) );
  NOR2X1 U26870 ( .A(n27313), .B(n27314), .Y(n27312) );
  NOR2X1 U26871 ( .A(n37749), .B(n26272), .Y(n27314) );
  NAND2X1 U26872 ( .A(n42581), .B(n42607), .Y(n26272) );
  NOR2X1 U26874 ( .A(n27315), .B(n73568), .Y(n27313) );
  NOR2X1 U26875 ( .A(n26315), .B(n73543), .Y(n27315) );
  NOR2X1 U26876 ( .A(n26270), .B(n42607), .Y(n26315) );
  NAND2X1 U26877 ( .A(n27316), .B(n27317), .Y(n36341) );
  NOR2X1 U26878 ( .A(n27318), .B(n27319), .Y(n27317) );
  NOR2X1 U26879 ( .A(n27320), .B(n27321), .Y(n27319) );
  NOR2X1 U26880 ( .A(n27322), .B(n27323), .Y(n27320) );
  NOR2X1 U26883 ( .A(n27324), .B(n27325), .Y(n27316) );
  AND2X1 U26884 ( .A(u_csr_N3161), .B(n27321), .Y(n27324) );
  NAND2X1 U26885 ( .A(n42607), .B(n27326), .Y(n27321) );
  NAND2X1 U26886 ( .A(n27327), .B(n27328), .Y(u_csr_csr_mip_r_9) );
  NAND2X1 U26887 ( .A(intr_i), .B(u_csr_csr_mideleg_q[9]), .Y(n27328) );
  NOR2X1 U26888 ( .A(n27329), .B(n27330), .Y(n27327) );
  NOR2X1 U26889 ( .A(n27331), .B(n37334), .Y(n27330) );
  NAND2X1 U26893 ( .A(n27335), .B(n27336), .Y(u_csr_csr_mip_r_7) );
  NAND2X1 U26895 ( .A(u_csr_csr_mip_q_7), .B(n27338), .Y(n27335) );
  NAND2X1 U26896 ( .A(n27339), .B(n27340), .Y(n27338) );
  NAND2X1 U26898 ( .A(n27343), .B(n27344), .Y(u_csr_csr_mip_r_5) );
  NAND2X1 U26899 ( .A(u_csr_csr_mip_q_5), .B(n27345), .Y(n27344) );
  NAND2X1 U26900 ( .A(n27346), .B(n27347), .Y(n27345) );
  NAND2X1 U26903 ( .A(n27349), .B(n27350), .Y(u_csr_csr_mip_r_3) );
  NAND2X1 U26904 ( .A(u_csr_csr_mip_q_3), .B(n27351), .Y(n27350) );
  NAND2X1 U26905 ( .A(n27340), .B(n27352), .Y(n27351) );
  AND2X1 U26906 ( .A(n27347), .B(n27353), .Y(n27340) );
  NAND2X1 U26908 ( .A(n27355), .B(n27356), .Y(u_csr_csr_mip_r_1) );
  NAND2X1 U26909 ( .A(u_csr_csr_mip_q_1), .B(n27357), .Y(n27356) );
  NAND2X1 U26910 ( .A(n27347), .B(n26978), .Y(n27357) );
  AND2X1 U26911 ( .A(n27358), .B(n889), .Y(n27347) );
  NAND2X1 U26912 ( .A(n73509), .B(n73403), .Y(n27355) );
  NAND2X1 U26913 ( .A(n27359), .B(n27360), .Y(\u_csr_csr_mip_r[11] ) );
  NAND2X1 U26914 ( .A(intr_i), .B(n37531), .Y(n27360) );
  NOR2X1 U26915 ( .A(n27361), .B(n27362), .Y(n27359) );
  NOR2X1 U26916 ( .A(n27363), .B(n37553), .Y(n27362) );
  NOR2X1 U26917 ( .A(n27332), .B(n27364), .Y(n27363) );
  NAND2X1 U26919 ( .A(n43002), .B(n73506), .Y(n27353) );
  NAND2X1 U26920 ( .A(n27367), .B(n27368), .Y(n27332) );
  NOR2X1 U26921 ( .A(n24877), .B(n27369), .Y(n27368) );
  NAND2X1 U26922 ( .A(n27342), .B(n27370), .Y(n27369) );
  NOR2X1 U26923 ( .A(n26261), .B(n27371), .Y(n27367) );
  NAND2X1 U26926 ( .A(n27373), .B(n27374), .Y(u_csr_csr_mie_r_9) );
  NAND2X1 U26929 ( .A(u_csr_csr_mie_q_9), .B(n27376), .Y(n27373) );
  NAND2X1 U26931 ( .A(n27378), .B(n27379), .Y(u_csr_csr_mie_r_7) );
  NAND2X1 U26934 ( .A(u_csr_csr_mie_q_7), .B(n27380), .Y(n27378) );
  NAND2X1 U26936 ( .A(n27382), .B(n27383), .Y(u_csr_csr_mie_r_5) );
  NAND2X1 U26937 ( .A(u_csr_csr_mie_q_5), .B(n27384), .Y(n27383) );
  NAND2X1 U26940 ( .A(n27385), .B(n27386), .Y(u_csr_csr_mie_r_3) );
  NAND2X1 U26941 ( .A(u_csr_csr_mie_q_3), .B(n27387), .Y(n27386) );
  NAND2X1 U26942 ( .A(n27388), .B(n27389), .Y(n27387) );
  NOR2X1 U26943 ( .A(n461), .B(n375), .Y(n27388) );
  NAND2X1 U26945 ( .A(n27391), .B(n27392), .Y(u_csr_csr_mie_r_1) );
  NAND2X1 U26946 ( .A(u_csr_csr_mie_q_1), .B(n27393), .Y(n27392) );
  NAND2X1 U26947 ( .A(n27389), .B(n26978), .Y(n27393) );
  NAND2X1 U26948 ( .A(n73509), .B(n73402), .Y(n27391) );
  NAND2X1 U26949 ( .A(n27394), .B(n27395), .Y(\u_csr_csr_mie_r[11] ) );
  NAND2X1 U26952 ( .A(\u_csr_csr_mie_q[11] ), .B(n27398), .Y(n27394) );
  AND2X1 U26954 ( .A(n27377), .B(n27390), .Y(n27381) );
  NAND2X1 U26955 ( .A(n43004), .B(n73405), .Y(n27390) );
  AND2X1 U26956 ( .A(n27389), .B(n27342), .Y(n27377) );
  AND2X1 U26957 ( .A(n27358), .B(n896), .Y(n27389) );
  AND2X1 U26958 ( .A(n27399), .B(n27400), .Y(n27358) );
  NOR2X1 U26959 ( .A(n884), .B(n27401), .Y(n27400) );
  NOR2X1 U26961 ( .A(n27402), .B(n27403), .Y(n27399) );
  NAND2X1 U26962 ( .A(n887), .B(n73576), .Y(n27403) );
  NAND2X1 U26979 ( .A(n27420), .B(n27421), .Y(u_csr_csr_mideleg_r[5]) );
  NAND2X1 U26980 ( .A(u_csr_csr_mideleg_q[5]), .B(n27422), .Y(n27421) );
  NAND2X1 U26983 ( .A(n27423), .B(n27424), .Y(u_csr_csr_mideleg_r[4]) );
  NAND2X1 U26984 ( .A(u_csr_csr_mideleg_q[4]), .B(n27425), .Y(n27424) );
  NAND2X1 U26985 ( .A(n27426), .B(n27427), .Y(n27425) );
  NAND2X1 U26987 ( .A(n27428), .B(n27429), .Y(u_csr_csr_mideleg_r[3]) );
  NAND2X1 U26988 ( .A(u_csr_csr_mideleg_q[3]), .B(n27430), .Y(n27429) );
  NAND2X1 U26989 ( .A(n27426), .B(n27352), .Y(n27430) );
  NAND2X1 U26991 ( .A(n27431), .B(n27432), .Y(u_csr_csr_mideleg_r[2]) );
  NAND2X1 U26992 ( .A(u_csr_csr_mideleg_q[2]), .B(n27433), .Y(n27432) );
  NAND2X1 U26993 ( .A(n27426), .B(n26959), .Y(n27433) );
  NAND2X1 U26995 ( .A(n27434), .B(n27435), .Y(u_csr_csr_mideleg_r[1]) );
  NAND2X1 U26996 ( .A(u_csr_csr_mideleg_q[1]), .B(n27436), .Y(n27435) );
  NAND2X1 U26997 ( .A(n27426), .B(n26978), .Y(n27436) );
  AND2X1 U27022 ( .A(n27426), .B(n27342), .Y(n27407) );
  NAND2X1 U27025 ( .A(n27461), .B(n27462), .Y(u_csr_csr_mideleg_r[0]) );
  NAND2X1 U27026 ( .A(u_csr_csr_mideleg_q[0]), .B(n27463), .Y(n27462) );
  NAND2X1 U27027 ( .A(n27426), .B(n27464), .Y(n27463) );
  AND2X1 U27028 ( .A(n27465), .B(n27208), .Y(n27426) );
  NAND2X1 U27601 ( .A(n27961), .B(n42131), .Y(n27960) );
  NOR2X1 U27602 ( .A(n73522), .B(n27964), .Y(n27961) );
  AND2X1 U27649 ( .A(n27560), .B(n26258), .Y(n27477) );
  AND2X1 U27667 ( .A(n28010), .B(n28011), .Y(n27560) );
  NOR2X1 U27668 ( .A(n28012), .B(n28013), .Y(n28011) );
  NAND2X1 U27669 ( .A(n28014), .B(n42983), .Y(n28013) );
  NOR2X1 U27670 ( .A(n73577), .B(n42963), .Y(n28012) );
  NOR2X1 U27671 ( .A(n26252), .B(n28015), .Y(n28010) );
  NAND2X1 U27672 ( .A(n462), .B(n27203), .Y(n28015) );
  NOR2X1 U27673 ( .A(n73399), .B(n42205), .Y(n27203) );
  NAND2X1 U27723 ( .A(n28056), .B(n28057), .Y(u_csr_csr_medeleg_r[5]) );
  NAND2X1 U27724 ( .A(u_csr_csr_medeleg_q[5]), .B(n28058), .Y(n28057) );
  NAND2X1 U27729 ( .A(n28059), .B(n28060), .Y(u_csr_csr_medeleg_r[4]) );
  NAND2X1 U27730 ( .A(u_csr_csr_medeleg_q[4]), .B(n28061), .Y(n28060) );
  NAND2X1 U27731 ( .A(n28062), .B(n27427), .Y(n28061) );
  NAND2X1 U27732 ( .A(n43003), .B(n25860), .Y(n27427) );
  NAND2X1 U27735 ( .A(n28064), .B(n28065), .Y(u_csr_csr_medeleg_r[3]) );
  NAND2X1 U27736 ( .A(u_csr_csr_medeleg_q[3]), .B(n28066), .Y(n28065) );
  NAND2X1 U27737 ( .A(n28062), .B(n27352), .Y(n28066) );
  NAND2X1 U27739 ( .A(n28067), .B(n28068), .Y(u_csr_csr_medeleg_r[2]) );
  NAND2X1 U27740 ( .A(u_csr_csr_medeleg_q[2]), .B(n28069), .Y(n28068) );
  NAND2X1 U27741 ( .A(n28062), .B(n26959), .Y(n28069) );
  NAND2X1 U27743 ( .A(n28070), .B(n28071), .Y(u_csr_csr_medeleg_r[1]) );
  NAND2X1 U27744 ( .A(u_csr_csr_medeleg_q[1]), .B(n28072), .Y(n28071) );
  NAND2X1 U27745 ( .A(n28062), .B(n26978), .Y(n28072) );
  AND2X1 U27776 ( .A(n28062), .B(n27342), .Y(n28045) );
  NAND2X1 U27780 ( .A(n28091), .B(n28092), .Y(u_csr_csr_medeleg_r[0]) );
  NAND2X1 U27781 ( .A(u_csr_csr_medeleg_q[0]), .B(n28093), .Y(n28092) );
  NAND2X1 U27782 ( .A(n28062), .B(n27464), .Y(n28093) );
  NAND2X1 U27783 ( .A(n43002), .B(n26127), .Y(n27464) );
  AND2X1 U27784 ( .A(n28094), .B(n27208), .Y(n28062) );
  AND2X1 U27785 ( .A(n27202), .B(n73577), .Y(n27208) );
  AND2X1 U27786 ( .A(n28095), .B(n73503), .Y(n27202) );
  AND2X1 U27787 ( .A(n42963), .B(n28014), .Y(n28095) );
  NAND2X1 U27788 ( .A(n42962), .B(n28096), .Y(n28014) );
  NAND2X1 U27789 ( .A(n28097), .B(n28098), .Y(n28096) );
  NOR2X1 U27792 ( .A(n27104), .B(n26133), .Y(n28097) );
  NAND2X1 U27793 ( .A(n73401), .B(n883), .Y(n26133) );
  NOR2X1 U27797 ( .A(n42205), .B(n41738), .Y(n28094) );
  XNOR2X1 U27801 ( .A(u_csr_csr_mcycle_q[9]), .B(n28100), .Y(
        u_csr_csr_mcycle_r[9]) );
  XNOR2X1 U27802 ( .A(n37571), .B(n28101), .Y(u_csr_csr_mcycle_r[8]) );
  NOR2X1 U27803 ( .A(n37346), .B(n28102), .Y(n28101) );
  XNOR2X1 U27804 ( .A(n37346), .B(n655), .Y(u_csr_csr_mcycle_r[7]) );
  XNOR2X1 U27805 ( .A(n37569), .B(n28103), .Y(u_csr_csr_mcycle_r[6]) );
  AND2X1 U27806 ( .A(u_csr_csr_mcycle_q[5]), .B(n28104), .Y(n28103) );
  XNOR2X1 U27807 ( .A(n37345), .B(n28104), .Y(u_csr_csr_mcycle_r[5]) );
  XNOR2X1 U27808 ( .A(n37721), .B(n28105), .Y(u_csr_csr_mcycle_r[4]) );
  NOR2X1 U27809 ( .A(n37693), .B(n28106), .Y(n28105) );
  XNOR2X1 U27810 ( .A(u_csr_csr_mcycle_q[3]), .B(n28106), .Y(
        u_csr_csr_mcycle_r[3]) );
  XNOR2X1 U27811 ( .A(n37729), .B(n28107), .Y(u_csr_csr_mcycle_r[31]) );
  NOR2X1 U27812 ( .A(n37699), .B(n28108), .Y(n28107) );
  XNOR2X1 U27813 ( .A(u_csr_csr_mcycle_q[30]), .B(n28108), .Y(
        u_csr_csr_mcycle_r[30]) );
  NAND2X1 U27814 ( .A(n28109), .B(u_csr_csr_mcycle_q[29]), .Y(n28108) );
  XNOR2X1 U27815 ( .A(n37563), .B(n28110), .Y(u_csr_csr_mcycle_r[2]) );
  NOR2X1 U27816 ( .A(n37343), .B(n8886), .Y(n28110) );
  XNOR2X1 U27817 ( .A(n37695), .B(n28109), .Y(u_csr_csr_mcycle_r[29]) );
  AND2X1 U27818 ( .A(n28111), .B(n28112), .Y(n28109) );
  NOR2X1 U27819 ( .A(n37598), .B(n37352), .Y(n28111) );
  XNOR2X1 U27820 ( .A(n37598), .B(n28113), .Y(u_csr_csr_mcycle_r[28]) );
  AND2X1 U27821 ( .A(u_csr_csr_mcycle_q[27]), .B(n28112), .Y(n28113) );
  XNOR2X1 U27822 ( .A(n37352), .B(n28112), .Y(u_csr_csr_mcycle_r[27]) );
  NOR2X1 U27823 ( .A(n28114), .B(n28115), .Y(n28112) );
  NAND2X1 U27824 ( .A(u_csr_csr_mcycle_q[26]), .B(u_csr_csr_mcycle_q[25]), .Y(
        n28114) );
  XNOR2X1 U27825 ( .A(n37698), .B(n28116), .Y(u_csr_csr_mcycle_r[26]) );
  NOR2X1 U27826 ( .A(n37691), .B(n28115), .Y(n28116) );
  XNOR2X1 U27827 ( .A(u_csr_csr_mcycle_q[25]), .B(n28115), .Y(
        u_csr_csr_mcycle_r[25]) );
  NAND2X1 U27828 ( .A(n28117), .B(n28118), .Y(n28115) );
  NOR2X1 U27829 ( .A(n37588), .B(n37350), .Y(n28117) );
  XNOR2X1 U27830 ( .A(n37588), .B(n28119), .Y(u_csr_csr_mcycle_r[24]) );
  AND2X1 U27831 ( .A(u_csr_csr_mcycle_q[23]), .B(n28118), .Y(n28119) );
  XNOR2X1 U27832 ( .A(n37350), .B(n28118), .Y(u_csr_csr_mcycle_r[23]) );
  NOR2X1 U27833 ( .A(n28120), .B(n28121), .Y(n28118) );
  NAND2X1 U27834 ( .A(u_csr_csr_mcycle_q[22]), .B(u_csr_csr_mcycle_q[21]), .Y(
        n28120) );
  XNOR2X1 U27835 ( .A(n37697), .B(n28122), .Y(u_csr_csr_mcycle_r[22]) );
  NOR2X1 U27836 ( .A(n37690), .B(n28121), .Y(n28122) );
  XNOR2X1 U27837 ( .A(u_csr_csr_mcycle_q[21]), .B(n28121), .Y(
        u_csr_csr_mcycle_r[21]) );
  NAND2X1 U27838 ( .A(n28123), .B(n28124), .Y(n28121) );
  NOR2X1 U27839 ( .A(n37585), .B(n37349), .Y(n28123) );
  XNOR2X1 U27840 ( .A(n37585), .B(n28125), .Y(u_csr_csr_mcycle_r[20]) );
  AND2X1 U27841 ( .A(u_csr_csr_mcycle_q[19]), .B(n28124), .Y(n28125) );
  XNOR2X1 U27842 ( .A(n8886), .B(u_csr_csr_mcycle_q[1]), .Y(
        u_csr_csr_mcycle_r[1]) );
  XNOR2X1 U27843 ( .A(n37349), .B(n28124), .Y(u_csr_csr_mcycle_r[19]) );
  NOR2X1 U27844 ( .A(n28126), .B(n28127), .Y(n28124) );
  NAND2X1 U27845 ( .A(u_csr_csr_mcycle_q[18]), .B(u_csr_csr_mcycle_q[17]), .Y(
        n28126) );
  XNOR2X1 U27846 ( .A(n37696), .B(n28128), .Y(u_csr_csr_mcycle_r[18]) );
  NOR2X1 U27847 ( .A(n37689), .B(n28127), .Y(n28128) );
  XNOR2X1 U27848 ( .A(u_csr_csr_mcycle_q[17]), .B(n28127), .Y(
        u_csr_csr_mcycle_r[17]) );
  NAND2X1 U27849 ( .A(n28129), .B(n28130), .Y(n28127) );
  NOR2X1 U27850 ( .A(n37578), .B(n37348), .Y(n28129) );
  XNOR2X1 U27851 ( .A(n37578), .B(n28131), .Y(u_csr_csr_mcycle_r[16]) );
  AND2X1 U27852 ( .A(u_csr_csr_mcycle_q[15]), .B(n28130), .Y(n28131) );
  XNOR2X1 U27853 ( .A(n37348), .B(n28130), .Y(u_csr_csr_mcycle_r[15]) );
  NOR2X1 U27854 ( .A(n28132), .B(n28133), .Y(n28130) );
  NAND2X1 U27855 ( .A(u_csr_csr_mcycle_q[14]), .B(u_csr_csr_mcycle_q[13]), .Y(
        n28132) );
  XNOR2X1 U27856 ( .A(n37712), .B(n28134), .Y(u_csr_csr_mcycle_r[14]) );
  NOR2X1 U27857 ( .A(n37692), .B(n28133), .Y(n28134) );
  XNOR2X1 U27858 ( .A(u_csr_csr_mcycle_q[13]), .B(n28133), .Y(
        u_csr_csr_mcycle_r[13]) );
  NAND2X1 U27859 ( .A(n28135), .B(n28136), .Y(n28133) );
  NOR2X1 U27860 ( .A(n37574), .B(n37347), .Y(n28135) );
  XNOR2X1 U27861 ( .A(n37574), .B(n28137), .Y(u_csr_csr_mcycle_r[12]) );
  AND2X1 U27862 ( .A(u_csr_csr_mcycle_q[11]), .B(n28136), .Y(n28137) );
  XNOR2X1 U27863 ( .A(n37347), .B(n28136), .Y(u_csr_csr_mcycle_r[11]) );
  NOR2X1 U27864 ( .A(n28138), .B(n28100), .Y(n28136) );
  NAND2X1 U27865 ( .A(u_csr_csr_mcycle_q[9]), .B(u_csr_csr_mcycle_q[10]), .Y(
        n28138) );
  XNOR2X1 U27866 ( .A(n37711), .B(n28139), .Y(u_csr_csr_mcycle_r[10]) );
  NOR2X1 U27867 ( .A(n37694), .B(n28100), .Y(n28139) );
  NAND2X1 U27868 ( .A(n28140), .B(n655), .Y(n28100) );
  NAND2X1 U27869 ( .A(n28141), .B(n28104), .Y(n28102) );
  NOR2X1 U27870 ( .A(n28142), .B(n28106), .Y(n28104) );
  NAND2X1 U27871 ( .A(n28143), .B(u_csr_csr_mcycle_q[0]), .Y(n28106) );
  NOR2X1 U27872 ( .A(n37563), .B(n37343), .Y(n28143) );
  NAND2X1 U27873 ( .A(u_csr_csr_mcycle_q[4]), .B(u_csr_csr_mcycle_q[3]), .Y(
        n28142) );
  NOR2X1 U27874 ( .A(n37569), .B(n37345), .Y(n28141) );
  NOR2X1 U27875 ( .A(n37571), .B(n37346), .Y(n28140) );
  NAND2X1 U27876 ( .A(n28144), .B(n28145), .Y(u_csr_csr_mcause_r_31) );
  NAND2X1 U27877 ( .A(u_csr_csr_mcause_q_31), .B(n28146), .Y(n28145) );
  NAND2X1 U27878 ( .A(n28147), .B(n26936), .Y(n28146) );
  NAND2X1 U27879 ( .A(n28148), .B(n28149), .Y(n26936) );
  NOR2X1 U27882 ( .A(n73518), .B(n28151), .Y(n28144) );
  NAND2X1 U27886 ( .A(n28153), .B(n28154), .Y(u_csr_csr_mcause_r[3]) );
  NOR2X1 U27887 ( .A(n28155), .B(n28156), .Y(n28154) );
  NAND2X1 U27888 ( .A(n28157), .B(n28158), .Y(n28156) );
  NAND2X1 U27889 ( .A(n42461), .B(n73516), .Y(n28158) );
  NAND2X1 U27892 ( .A(u_csr_csr_mcause_q[3]), .B(n28161), .Y(n28157) );
  NAND2X1 U27893 ( .A(n28162), .B(n27352), .Y(n28161) );
  NAND2X1 U27894 ( .A(n43004), .B(n25872), .Y(n27352) );
  NOR2X1 U27896 ( .A(n28164), .B(n28165), .Y(n28153) );
  NOR2X1 U27897 ( .A(n1082), .B(n28035), .Y(n28165) );
  NAND2X1 U27903 ( .A(n28169), .B(n28170), .Y(u_csr_csr_mcause_r[2]) );
  NOR2X1 U27904 ( .A(n28171), .B(n28172), .Y(n28170) );
  NOR2X1 U27908 ( .A(n1083), .B(n28174), .Y(n26957) );
  NOR2X1 U27909 ( .A(n28176), .B(n37775), .Y(n28171) );
  AND2X1 U27910 ( .A(n26959), .B(n28162), .Y(n28176) );
  NAND2X1 U27911 ( .A(n43003), .B(n25903), .Y(n26959) );
  NOR2X1 U27912 ( .A(n28177), .B(n28178), .Y(n28169) );
  NOR2X1 U27915 ( .A(n26962), .B(n28179), .Y(n28177) );
  AND2X1 U27916 ( .A(n26138), .B(n28180), .Y(n26962) );
  NAND2X1 U27917 ( .A(n73420), .B(n28181), .Y(n28180) );
  NAND2X1 U27918 ( .A(n28182), .B(n28183), .Y(u_csr_csr_mcause_r[1]) );
  NOR2X1 U27919 ( .A(n28184), .B(n28185), .Y(n28183) );
  NAND2X1 U27920 ( .A(n28186), .B(n28187), .Y(n28185) );
  NAND2X1 U27921 ( .A(n26969), .B(n73518), .Y(n28186) );
  NOR2X1 U27922 ( .A(n1085), .B(n28188), .Y(n26969) );
  AND2X1 U27923 ( .A(n28189), .B(n28190), .Y(n28188) );
  NAND2X1 U27924 ( .A(n28191), .B(n28192), .Y(n28190) );
  NAND2X1 U27925 ( .A(n28193), .B(n28194), .Y(n28191) );
  NOR2X1 U27926 ( .A(n28179), .B(n28196), .Y(n28184) );
  NAND2X1 U27927 ( .A(n8810), .B(n26971), .Y(n28196) );
  NAND2X1 U27932 ( .A(n73420), .B(n28203), .Y(n28202) );
  OR2X1 U27933 ( .A(n28204), .B(n73419), .Y(n28203) );
  NOR2X1 U27934 ( .A(n28205), .B(n28206), .Y(n28182) );
  NAND2X1 U27935 ( .A(n28207), .B(n28208), .Y(n28206) );
  NAND2X1 U27936 ( .A(u_csr_csr_mcause_q[1]), .B(n28209), .Y(n28208) );
  NAND2X1 U27937 ( .A(n28162), .B(n26978), .Y(n28209) );
  NAND2X1 U27938 ( .A(n43002), .B(n26014), .Y(n26978) );
  NOR2X1 U27940 ( .A(n28210), .B(n26977), .Y(n28162) );
  NAND2X1 U27941 ( .A(n462), .B(n28211), .Y(n26977) );
  NAND2X1 U27942 ( .A(n42962), .B(n28212), .Y(n28211) );
  NAND2X1 U27943 ( .A(n28213), .B(n883), .Y(n28212) );
  NOR2X1 U27944 ( .A(n73539), .B(n28215), .Y(n28213) );
  NAND2X1 U27945 ( .A(n26270), .B(n26327), .Y(n26913) );
  NAND2X1 U27946 ( .A(n42215), .B(n28031), .Y(n26270) );
  NAND2X1 U27947 ( .A(n25083), .B(n73507), .Y(n28210) );
  NAND2X1 U27952 ( .A(n465), .B(u_csr_N3162), .Y(n28207) );
  NAND2X1 U27958 ( .A(n28220), .B(n28221), .Y(u_csr_csr_mcause_r[0]) );
  NOR2X1 U27959 ( .A(n28222), .B(n28223), .Y(n28221) );
  NAND2X1 U27960 ( .A(n28035), .B(n28187), .Y(n28223) );
  NAND2X1 U27961 ( .A(n28224), .B(n466), .Y(n28187) );
  NOR2X1 U27963 ( .A(n28179), .B(n28225), .Y(n28222) );
  NOR2X1 U27967 ( .A(n28228), .B(n28229), .Y(n28220) );
  NAND2X1 U27968 ( .A(n28230), .B(n28231), .Y(n28229) );
  NAND2X1 U27969 ( .A(u_csr_csr_mcause_q[0]), .B(n28232), .Y(n28231) );
  NAND2X1 U27970 ( .A(n28147), .B(n26992), .Y(n28232) );
  NAND2X1 U27971 ( .A(n28148), .B(n28233), .Y(n26992) );
  NOR2X1 U27972 ( .A(n73575), .B(n73521), .Y(n28233) );
  NOR2X1 U27973 ( .A(n27326), .B(n28235), .Y(n28148) );
  NOR2X1 U27974 ( .A(n28236), .B(n26998), .Y(n28147) );
  NAND2X1 U27975 ( .A(n28237), .B(n474), .Y(n26998) );
  NAND2X1 U27976 ( .A(n28238), .B(n73418), .Y(n28237) );
  NOR2X1 U27977 ( .A(n27318), .B(n28239), .Y(n28238) );
  NOR2X1 U27978 ( .A(n28214), .B(n27402), .Y(n28239) );
  NAND2X1 U27979 ( .A(n28240), .B(n28241), .Y(n27402) );
  NOR2X1 U27982 ( .A(n27326), .B(n28215), .Y(n28240) );
  NAND2X1 U27983 ( .A(n28243), .B(n28244), .Y(n28214) );
  NOR2X1 U27984 ( .A(n884), .B(n73402), .Y(n28244) );
  NOR2X1 U27985 ( .A(n28031), .B(n73543), .Y(n27318) );
  OR2X1 U27986 ( .A(n28245), .B(n28246), .Y(n28236) );
  NOR2X1 U27987 ( .A(n28247), .B(n73516), .Y(n28246) );
  NOR2X1 U27988 ( .A(n73517), .B(n73574), .Y(n28247) );
  NAND2X1 U27991 ( .A(n465), .B(u_csr_N3161), .Y(n28230) );
  NAND2X1 U27993 ( .A(n42215), .B(n28249), .Y(n28032) );
  NAND2X1 U28001 ( .A(n474), .B(n28031), .Y(n28252) );
  NAND2X1 U28008 ( .A(reset_vector_i[31]), .B(n44639), .Y(n28256) );
  NOR2X1 U28011 ( .A(n28262), .B(n28263), .Y(n28259) );
  NOR2X1 U28012 ( .A(n28264), .B(n1172), .Y(n28263) );
  NOR2X1 U28013 ( .A(n44268), .B(n37745), .Y(n28262) );
  NAND2X1 U28017 ( .A(reset_vector_i[30]), .B(n8572), .Y(n28268) );
  NOR2X1 U28020 ( .A(n28272), .B(n28273), .Y(n28270) );
  NOR2X1 U28021 ( .A(n28264), .B(n1173), .Y(n28273) );
  NOR2X1 U28022 ( .A(n44268), .B(n37744), .Y(n28272) );
  NAND2X1 U28026 ( .A(reset_vector_i[29]), .B(n8572), .Y(n28276) );
  NOR2X1 U28029 ( .A(n28280), .B(n28281), .Y(n28278) );
  NOR2X1 U28030 ( .A(n28264), .B(n1175), .Y(n28281) );
  NOR2X1 U28031 ( .A(n44268), .B(n37743), .Y(n28280) );
  NAND2X1 U28035 ( .A(reset_vector_i[28]), .B(n8572), .Y(n28284) );
  NOR2X1 U28038 ( .A(n28288), .B(n28289), .Y(n28286) );
  NOR2X1 U28039 ( .A(n28264), .B(n1176), .Y(n28289) );
  NOR2X1 U28040 ( .A(n44268), .B(n37742), .Y(n28288) );
  NAND2X1 U28044 ( .A(reset_vector_i[27]), .B(n8572), .Y(n28292) );
  NOR2X1 U28047 ( .A(n28296), .B(n28297), .Y(n28294) );
  NOR2X1 U28048 ( .A(n28264), .B(n1177), .Y(n28297) );
  NOR2X1 U28049 ( .A(n44268), .B(n37741), .Y(n28296) );
  NAND2X1 U28053 ( .A(reset_vector_i[26]), .B(n8572), .Y(n28300) );
  NOR2X1 U28056 ( .A(n28304), .B(n28305), .Y(n28302) );
  NOR2X1 U28057 ( .A(n28264), .B(n1178), .Y(n28305) );
  NOR2X1 U28058 ( .A(n44268), .B(n37740), .Y(n28304) );
  NAND2X1 U28062 ( .A(reset_vector_i[25]), .B(n8572), .Y(n28308) );
  NOR2X1 U28065 ( .A(n28312), .B(n28313), .Y(n28310) );
  NOR2X1 U28066 ( .A(n28264), .B(n1179), .Y(n28313) );
  NOR2X1 U28067 ( .A(n44268), .B(n37739), .Y(n28312) );
  NAND2X1 U28071 ( .A(reset_vector_i[24]), .B(n8572), .Y(n28316) );
  NOR2X1 U28074 ( .A(n28320), .B(n28321), .Y(n28318) );
  NOR2X1 U28075 ( .A(n28264), .B(n1180), .Y(n28321) );
  NOR2X1 U28076 ( .A(n44268), .B(n37738), .Y(n28320) );
  NAND2X1 U28080 ( .A(reset_vector_i[23]), .B(n44639), .Y(n28324) );
  NOR2X1 U28083 ( .A(n28328), .B(n28329), .Y(n28326) );
  NOR2X1 U28084 ( .A(n44270), .B(n1181), .Y(n28329) );
  NOR2X1 U28085 ( .A(n44267), .B(n37737), .Y(n28328) );
  NAND2X1 U28089 ( .A(reset_vector_i[22]), .B(n44639), .Y(n28332) );
  NOR2X1 U28092 ( .A(n28336), .B(n28337), .Y(n28334) );
  NOR2X1 U28093 ( .A(n44270), .B(n1182), .Y(n28337) );
  NOR2X1 U28094 ( .A(n44267), .B(n37736), .Y(n28336) );
  NAND2X1 U28098 ( .A(reset_vector_i[21]), .B(n44639), .Y(n28340) );
  NOR2X1 U28101 ( .A(n28344), .B(n28345), .Y(n28342) );
  NOR2X1 U28102 ( .A(n44270), .B(n1183), .Y(n28345) );
  NOR2X1 U28103 ( .A(n44267), .B(n37735), .Y(n28344) );
  NAND2X1 U28107 ( .A(reset_vector_i[20]), .B(n44639), .Y(n28348) );
  NOR2X1 U28110 ( .A(n28352), .B(n28353), .Y(n28350) );
  NOR2X1 U28111 ( .A(n44270), .B(n1184), .Y(n28353) );
  NOR2X1 U28112 ( .A(n44267), .B(n37734), .Y(n28352) );
  NAND2X1 U28116 ( .A(reset_vector_i[19]), .B(n44639), .Y(n28356) );
  NOR2X1 U28119 ( .A(n28360), .B(n28361), .Y(n28358) );
  NOR2X1 U28120 ( .A(n44270), .B(n1186), .Y(n28361) );
  NOR2X1 U28121 ( .A(n44267), .B(n37733), .Y(n28360) );
  NAND2X1 U28125 ( .A(reset_vector_i[18]), .B(n44639), .Y(n28364) );
  NOR2X1 U28128 ( .A(n28368), .B(n28369), .Y(n28366) );
  NOR2X1 U28129 ( .A(n44270), .B(n1187), .Y(n28369) );
  NOR2X1 U28130 ( .A(n44267), .B(n37732), .Y(n28368) );
  NAND2X1 U28134 ( .A(reset_vector_i[17]), .B(n44639), .Y(n28372) );
  NOR2X1 U28137 ( .A(n28376), .B(n28377), .Y(n28374) );
  NOR2X1 U28138 ( .A(n44270), .B(n1188), .Y(n28377) );
  NOR2X1 U28139 ( .A(n44267), .B(n37731), .Y(n28376) );
  NAND2X1 U28143 ( .A(reset_vector_i[16]), .B(n44639), .Y(n28380) );
  NOR2X1 U28146 ( .A(n28384), .B(n28385), .Y(n28382) );
  NOR2X1 U28147 ( .A(n44270), .B(n1189), .Y(n28385) );
  NOR2X1 U28148 ( .A(n44267), .B(n37730), .Y(n28384) );
  NAND2X1 U28152 ( .A(reset_vector_i[15]), .B(n44639), .Y(n28388) );
  NOR2X1 U28155 ( .A(n28392), .B(n28393), .Y(n28390) );
  NOR2X1 U28156 ( .A(n44270), .B(n1190), .Y(n28393) );
  NOR2X1 U28157 ( .A(n44267), .B(n37719), .Y(n28392) );
  NAND2X1 U28161 ( .A(reset_vector_i[14]), .B(n44639), .Y(n28396) );
  NOR2X1 U28164 ( .A(n28400), .B(n28401), .Y(n28398) );
  NOR2X1 U28165 ( .A(n44270), .B(n1191), .Y(n28401) );
  NOR2X1 U28166 ( .A(n44267), .B(n37718), .Y(n28400) );
  NAND2X1 U28170 ( .A(reset_vector_i[13]), .B(n44640), .Y(n28404) );
  NOR2X1 U28173 ( .A(n28408), .B(n28409), .Y(n28406) );
  NOR2X1 U28174 ( .A(n44270), .B(n1192), .Y(n28409) );
  NOR2X1 U28175 ( .A(n44267), .B(n37717), .Y(n28408) );
  NAND2X1 U28179 ( .A(reset_vector_i[12]), .B(n44640), .Y(n28412) );
  NOR2X1 U28182 ( .A(n28416), .B(n28417), .Y(n28414) );
  NOR2X1 U28183 ( .A(n44270), .B(n1193), .Y(n28417) );
  NOR2X1 U28184 ( .A(n44267), .B(n37720), .Y(n28416) );
  NAND2X1 U28188 ( .A(reset_vector_i[11]), .B(n44640), .Y(n28420) );
  NOR2X1 U28191 ( .A(n28424), .B(n28425), .Y(n28422) );
  NOR2X1 U28192 ( .A(n44269), .B(n1225), .Y(n28425) );
  NOR2X1 U28193 ( .A(n44266), .B(n37708), .Y(n28424) );
  NAND2X1 U28197 ( .A(reset_vector_i[10]), .B(n44640), .Y(n28428) );
  NOR2X1 U28200 ( .A(n28432), .B(n28433), .Y(n28430) );
  NOR2X1 U28201 ( .A(n44269), .B(n1194), .Y(n28433) );
  NOR2X1 U28202 ( .A(n44266), .B(n37704), .Y(n28432) );
  NAND2X1 U28206 ( .A(reset_vector_i[9]), .B(n44640), .Y(n28436) );
  NOR2X1 U28209 ( .A(n28440), .B(n28441), .Y(n28438) );
  NOR2X1 U28210 ( .A(n44269), .B(n1165), .Y(n28441) );
  NOR2X1 U28211 ( .A(n44266), .B(n37716), .Y(n28440) );
  NAND2X1 U28215 ( .A(reset_vector_i[8]), .B(n44640), .Y(n28444) );
  NOR2X1 U28218 ( .A(n28448), .B(n28449), .Y(n28446) );
  NOR2X1 U28219 ( .A(n44269), .B(n1166), .Y(n28449) );
  NOR2X1 U28220 ( .A(n44266), .B(n37710), .Y(n28448) );
  NAND2X1 U28224 ( .A(reset_vector_i[7]), .B(n44640), .Y(n28452) );
  NOR2X1 U28227 ( .A(n28456), .B(n28457), .Y(n28454) );
  NOR2X1 U28228 ( .A(n44269), .B(n1167), .Y(n28457) );
  NOR2X1 U28229 ( .A(n44266), .B(n37715), .Y(n28456) );
  NAND2X1 U28233 ( .A(reset_vector_i[6]), .B(n44640), .Y(n28460) );
  NOR2X1 U28236 ( .A(n28464), .B(n28465), .Y(n28462) );
  NOR2X1 U28237 ( .A(n44269), .B(n1168), .Y(n28465) );
  NOR2X1 U28238 ( .A(n44266), .B(n37706), .Y(n28464) );
  NAND2X1 U28242 ( .A(reset_vector_i[5]), .B(n44640), .Y(n28468) );
  NOR2X1 U28245 ( .A(n28472), .B(n28473), .Y(n28470) );
  NOR2X1 U28246 ( .A(n44269), .B(n1169), .Y(n28473) );
  NOR2X1 U28247 ( .A(n44266), .B(n37714), .Y(n28472) );
  NAND2X1 U28251 ( .A(reset_vector_i[4]), .B(n44640), .Y(n28476) );
  NOR2X1 U28254 ( .A(n28480), .B(n28481), .Y(n28478) );
  NOR2X1 U28255 ( .A(n44269), .B(n37701), .Y(n28481) );
  NOR2X1 U28256 ( .A(n44266), .B(n37705), .Y(n28480) );
  NAND2X1 U28260 ( .A(reset_vector_i[3]), .B(n44640), .Y(n28484) );
  NOR2X1 U28263 ( .A(n28488), .B(n28489), .Y(n28486) );
  NOR2X1 U28264 ( .A(n44269), .B(n37723), .Y(n28489) );
  NOR2X1 U28265 ( .A(n44266), .B(n37700), .Y(n28488) );
  NAND2X1 U28269 ( .A(reset_vector_i[2]), .B(n44640), .Y(n28492) );
  NOR2X1 U28272 ( .A(n28496), .B(n28497), .Y(n28494) );
  NOR2X1 U28273 ( .A(n44269), .B(n37703), .Y(n28497) );
  NOR2X1 U28274 ( .A(n44266), .B(n37709), .Y(n28496) );
  NAND2X1 U28278 ( .A(reset_vector_i[1]), .B(n1751), .Y(n28500) );
  NOR2X1 U28281 ( .A(n28504), .B(n28505), .Y(n28502) );
  NOR2X1 U28282 ( .A(n44269), .B(n37722), .Y(n28505) );
  NOR2X1 U28283 ( .A(n44266), .B(n37713), .Y(n28504) );
  NAND2X1 U28289 ( .A(reset_vector_i[0]), .B(n1751), .Y(n28508) );
  NOR2X1 U28294 ( .A(n971), .B(n28515), .Y(n28510) );
  NOR2X1 U28295 ( .A(n28516), .B(n28517), .Y(n28512) );
  NOR2X1 U28296 ( .A(n44269), .B(n37702), .Y(n28517) );
  AND2X1 U28297 ( .A(n28518), .B(n28519), .Y(n28264) );
  NAND2X1 U28298 ( .A(n463), .B(n73574), .Y(n28519) );
  NAND2X1 U28299 ( .A(n8805), .B(n26920), .Y(n28518) );
  NOR2X1 U28302 ( .A(n44266), .B(n37707), .Y(n28516) );
  NAND2X1 U28304 ( .A(n28523), .B(n463), .Y(n28522) );
  NAND2X1 U28305 ( .A(n8805), .B(n73576), .Y(n28515) );
  NOR2X1 U28306 ( .A(n73574), .B(n28524), .Y(n28523) );
  NAND2X1 U28307 ( .A(n73568), .B(n28525), .Y(n28249) );
  NAND2X1 U28308 ( .A(n28526), .B(n28527), .Y(n28525) );
  NAND2X1 U28309 ( .A(n73544), .B(n28528), .Y(n28527) );
  NAND2X1 U28310 ( .A(n28529), .B(n28530), .Y(n28528) );
  NAND2X1 U28312 ( .A(n28532), .B(n28533), .Y(n28531) );
  NAND2X1 U28313 ( .A(u_csr_csr_medeleg_q[8]), .B(n73569), .Y(n28533) );
  NAND2X1 U28314 ( .A(u_csr_csr_medeleg_q[9]), .B(u_csr_N3161), .Y(n28532) );
  NAND2X1 U28316 ( .A(n8805), .B(n26976), .Y(n28521) );
  AND2X1 U28323 ( .A(n28537), .B(n28538), .Y(n28526) );
  NOR2X1 U28324 ( .A(n28539), .B(n28540), .Y(n28538) );
  NAND2X1 U28325 ( .A(n28541), .B(n28542), .Y(n28540) );
  NAND2X1 U28326 ( .A(n28543), .B(u_csr_csr_medeleg_q[5]), .Y(n28542) );
  NOR2X1 U28327 ( .A(n28544), .B(n575), .Y(n28543) );
  NAND2X1 U28328 ( .A(n73419), .B(u_csr_csr_medeleg_q[1]), .Y(n28541) );
  NOR2X1 U28329 ( .A(n37566), .B(n28204), .Y(n28539) );
  NOR2X1 U28330 ( .A(n28536), .B(n28545), .Y(n28537) );
  NAND2X1 U28331 ( .A(n28546), .B(n28547), .Y(n28545) );
  NAND2X1 U28332 ( .A(n73520), .B(u_csr_csr_medeleg_q[12]), .Y(n28547) );
  NAND2X1 U28333 ( .A(u_csr_csr_medeleg_q[2]), .B(n28227), .Y(n28546) );
  NOR2X1 U28335 ( .A(n28550), .B(n28551), .Y(n28549) );
  NAND2X1 U28349 ( .A(n28561), .B(n28562), .Y(n28560) );
  NOR2X1 U28350 ( .A(n24367), .B(n28563), .Y(n28562) );
  NOR2X1 U28352 ( .A(n27964), .B(n971), .Y(n28561) );
  NAND2X1 U28375 ( .A(n28578), .B(n28579), .Y(u_csr_N2391) );
  NAND2X1 U28378 ( .A(n28582), .B(n37776), .Y(n28578) );
  AND2X1 U28420 ( .A(n26361), .B(n28607), .Y(n28567) );
  NAND2X1 U28421 ( .A(n73405), .B(n28234), .Y(n28607) );
  NOR2X1 U28422 ( .A(n26328), .B(n973), .Y(n26361) );
  NAND2X1 U28423 ( .A(n28608), .B(n28234), .Y(n27096) );
  NAND2X1 U28424 ( .A(n73577), .B(n27964), .Y(n28234) );
  NAND2X1 U28425 ( .A(n73522), .B(n73577), .Y(n28608) );
  NAND2X1 U28428 ( .A(n28610), .B(n28611), .Y(u_csr_N2377) );
  NAND2X1 U28429 ( .A(u_csr_csr_sr_q[4]), .B(n28612), .Y(n28611) );
  NAND2X1 U28430 ( .A(n28613), .B(n25681), .Y(n28612) );
  NAND2X1 U28431 ( .A(n44082), .B(n25860), .Y(n25681) );
  NAND2X1 U28432 ( .A(n73404), .B(n73504), .Y(n28610) );
  NAND2X1 U28436 ( .A(n28616), .B(n28617), .Y(u_csr_N2375) );
  NAND2X1 U28437 ( .A(n37567), .B(n73505), .Y(n28617) );
  NAND2X1 U28439 ( .A(u_csr_csr_sr_q[2]), .B(n28618), .Y(n28616) );
  NAND2X1 U28440 ( .A(n28619), .B(n28613), .Y(n28618) );
  NOR2X1 U28441 ( .A(n388), .B(n28620), .Y(n28619) );
  NOR2X1 U28442 ( .A(n27964), .B(n28621), .Y(n28620) );
  NAND2X1 U28443 ( .A(n44082), .B(n25903), .Y(n25699) );
  NAND2X1 U28447 ( .A(n28624), .B(n28625), .Y(u_csr_N2373) );
  NAND2X1 U28448 ( .A(u_csr_csr_sr_q[0]), .B(n28626), .Y(n28625) );
  NAND2X1 U28449 ( .A(n28613), .B(n25791), .Y(n28626) );
  NAND2X1 U28450 ( .A(n44082), .B(n26127), .Y(n25791) );
  NOR2X1 U28451 ( .A(n26328), .B(n26129), .Y(n28613) );
  NAND2X1 U28452 ( .A(n28627), .B(n885), .Y(n26328) );
  NOR2X1 U28453 ( .A(n884), .B(n73403), .Y(n28627) );
  NAND2X1 U28454 ( .A(n28243), .B(n885), .Y(n27370) );
  NAND2X1 U28455 ( .A(n28628), .B(n28629), .Y(n27371) );
  NOR2X1 U28460 ( .A(n73402), .B(n28215), .Y(n28628) );
  NAND2X1 U28461 ( .A(n28632), .B(n28633), .Y(n28215) );
  NOR2X1 U28467 ( .A(n28636), .B(n27104), .Y(n28632) );
  NOR2X1 U28478 ( .A(n26261), .B(n73403), .Y(n28243) );
  NAND2X1 U28485 ( .A(n73404), .B(n73521), .Y(n28624) );
  NOR2X1 U28676 ( .A(mem_d_accept_i), .B(n28734), .Y(n8558) );
  NOR2X1 U28677 ( .A(n28735), .B(n28736), .Y(n28734) );
  OR2X1 U28678 ( .A(mem_d_wr_o[0]), .B(u_arb_read_hold_q), .Y(n28736) );
  NAND2X1 U28679 ( .A(n28737), .B(n28738), .Y(n8557) );
  NAND2X1 U28680 ( .A(u_arb_src_mmu_q), .B(n28739), .Y(n28738) );
  NAND2X1 U28681 ( .A(n440), .B(n28740), .Y(n28739) );
  NAND2X1 U28682 ( .A(n28741), .B(n692), .Y(n28740) );
  NAND2X1 U28683 ( .A(n28742), .B(n28743), .Y(n28735) );
  NOR2X1 U28684 ( .A(mem_d_rd_o), .B(mem_d_wr_o[3]), .Y(n28743) );
  NAND2X1 U28685 ( .A(n28744), .B(n28745), .Y(mem_d_rd_o) );
  NOR2X1 U28694 ( .A(mem_d_wr_o[2]), .B(mem_d_wr_o[1]), .Y(n28742) );
  NAND2X1 U28700 ( .A(n44257), .B(n440), .Y(n28737) );
  NAND2X1 U28717 ( .A(n28776), .B(n28777), .Y(n8550) );
  NAND2X1 U28718 ( .A(mem_d_data_rd_i[22]), .B(n42978), .Y(n28777) );
  NAND2X1 U28719 ( .A(u_mmu_pte_entry_q[24]), .B(n73538), .Y(n28776) );
  NAND2X1 U28720 ( .A(n28778), .B(n28779), .Y(n8549) );
  NAND2X1 U28721 ( .A(mem_d_data_rd_i[23]), .B(n42979), .Y(n28779) );
  NAND2X1 U28722 ( .A(u_mmu_pte_entry_q[25]), .B(n73538), .Y(n28778) );
  NAND2X1 U28723 ( .A(n28780), .B(n28781), .Y(n8548) );
  NAND2X1 U28724 ( .A(mem_d_data_rd_i[24]), .B(n42978), .Y(n28781) );
  NAND2X1 U28725 ( .A(u_mmu_pte_entry_q[26]), .B(n73538), .Y(n28780) );
  NAND2X1 U28726 ( .A(n28782), .B(n28783), .Y(n8547) );
  NAND2X1 U28727 ( .A(mem_d_data_rd_i[25]), .B(n42979), .Y(n28783) );
  NAND2X1 U28728 ( .A(u_mmu_pte_entry_q[27]), .B(n73538), .Y(n28782) );
  NAND2X1 U28729 ( .A(n28784), .B(n28785), .Y(n8546) );
  NAND2X1 U28730 ( .A(mem_d_data_rd_i[26]), .B(n42978), .Y(n28785) );
  NAND2X1 U28731 ( .A(u_mmu_pte_entry_q[28]), .B(n73538), .Y(n28784) );
  NAND2X1 U28732 ( .A(n28786), .B(n28787), .Y(n8545) );
  NAND2X1 U28733 ( .A(mem_d_data_rd_i[27]), .B(n42979), .Y(n28787) );
  NAND2X1 U28734 ( .A(u_mmu_pte_entry_q[29]), .B(n73538), .Y(n28786) );
  NAND2X1 U28735 ( .A(n28788), .B(n28789), .Y(n8544) );
  NAND2X1 U28736 ( .A(mem_d_data_rd_i[28]), .B(n42978), .Y(n28789) );
  NAND2X1 U28737 ( .A(u_mmu_pte_entry_q[30]), .B(n73538), .Y(n28788) );
  NAND2X1 U28738 ( .A(n28790), .B(n28791), .Y(n8543) );
  NAND2X1 U28739 ( .A(mem_d_data_rd_i[29]), .B(n42979), .Y(n28791) );
  NAND2X1 U28745 ( .A(u_mmu_pte_entry_q[31]), .B(n73538), .Y(n28790) );
  NAND2X1 U28767 ( .A(n28813), .B(n28814), .Y(n8536) );
  NAND2X1 U28768 ( .A(u_muldiv_q_mask_q[31]), .B(n44624), .Y(n28814) );
  NAND2X1 U28769 ( .A(n28815), .B(n28816), .Y(n8535) );
  NAND2X1 U28770 ( .A(u_muldiv_q_mask_q[18]), .B(n44616), .Y(n28816) );
  NAND2X1 U28771 ( .A(u_muldiv_q_mask_q[17]), .B(n441), .Y(n28815) );
  NAND2X1 U28772 ( .A(n28817), .B(n28818), .Y(n8534) );
  NAND2X1 U28773 ( .A(u_muldiv_q_mask_q[19]), .B(n44616), .Y(n28818) );
  NAND2X1 U28774 ( .A(u_muldiv_q_mask_q[18]), .B(n441), .Y(n28817) );
  NAND2X1 U28775 ( .A(n28819), .B(n28820), .Y(n8533) );
  NAND2X1 U28776 ( .A(u_muldiv_q_mask_q[20]), .B(n44614), .Y(n28820) );
  NAND2X1 U28777 ( .A(u_muldiv_q_mask_q[19]), .B(n441), .Y(n28819) );
  NAND2X1 U28778 ( .A(n28821), .B(n28822), .Y(n8532) );
  NAND2X1 U28779 ( .A(u_muldiv_q_mask_q[21]), .B(n44614), .Y(n28822) );
  NAND2X1 U28780 ( .A(u_muldiv_q_mask_q[20]), .B(n441), .Y(n28821) );
  NAND2X1 U28781 ( .A(n28823), .B(n28824), .Y(n8531) );
  NAND2X1 U28782 ( .A(u_muldiv_q_mask_q[22]), .B(n44614), .Y(n28824) );
  NAND2X1 U28783 ( .A(u_muldiv_q_mask_q[21]), .B(n441), .Y(n28823) );
  NAND2X1 U28784 ( .A(n28825), .B(n28826), .Y(n8530) );
  NAND2X1 U28785 ( .A(u_muldiv_q_mask_q[23]), .B(n44614), .Y(n28826) );
  NAND2X1 U28786 ( .A(u_muldiv_q_mask_q[22]), .B(n441), .Y(n28825) );
  NAND2X1 U28787 ( .A(n28827), .B(n28828), .Y(n8529) );
  NAND2X1 U28788 ( .A(u_muldiv_q_mask_q[24]), .B(n44614), .Y(n28828) );
  NAND2X1 U28789 ( .A(u_muldiv_q_mask_q[23]), .B(n441), .Y(n28827) );
  NAND2X1 U28790 ( .A(n28829), .B(n28830), .Y(n8528) );
  NAND2X1 U28791 ( .A(u_muldiv_q_mask_q[25]), .B(n44614), .Y(n28830) );
  NAND2X1 U28792 ( .A(u_muldiv_q_mask_q[24]), .B(n441), .Y(n28829) );
  NAND2X1 U28793 ( .A(n28831), .B(n28832), .Y(n8527) );
  NAND2X1 U28794 ( .A(u_muldiv_q_mask_q[26]), .B(n44614), .Y(n28832) );
  NAND2X1 U28795 ( .A(u_muldiv_q_mask_q[25]), .B(n441), .Y(n28831) );
  NAND2X1 U28796 ( .A(n28833), .B(n28834), .Y(n8526) );
  NAND2X1 U28797 ( .A(u_muldiv_q_mask_q[27]), .B(n44614), .Y(n28834) );
  NAND2X1 U28798 ( .A(u_muldiv_q_mask_q[26]), .B(n441), .Y(n28833) );
  NAND2X1 U28799 ( .A(n28835), .B(n28836), .Y(n8525) );
  NAND2X1 U28800 ( .A(u_muldiv_q_mask_q[28]), .B(n44614), .Y(n28836) );
  NAND2X1 U28801 ( .A(u_muldiv_q_mask_q[27]), .B(n441), .Y(n28835) );
  NAND2X1 U28802 ( .A(n28837), .B(n28838), .Y(n8524) );
  NAND2X1 U28803 ( .A(u_muldiv_q_mask_q[29]), .B(n44615), .Y(n28838) );
  NAND2X1 U28804 ( .A(u_muldiv_q_mask_q[28]), .B(n441), .Y(n28837) );
  NAND2X1 U28805 ( .A(n28839), .B(n28840), .Y(n8523) );
  NAND2X1 U28806 ( .A(u_muldiv_q_mask_q[30]), .B(n44615), .Y(n28840) );
  NAND2X1 U28807 ( .A(u_muldiv_q_mask_q[29]), .B(n441), .Y(n28839) );
  NAND2X1 U28808 ( .A(n28841), .B(n28842), .Y(n8522) );
  NAND2X1 U28809 ( .A(u_muldiv_q_mask_q[31]), .B(n44615), .Y(n28842) );
  NAND2X1 U28810 ( .A(u_muldiv_q_mask_q[30]), .B(n441), .Y(n28841) );
  NAND2X1 U28811 ( .A(n28843), .B(n28844), .Y(n8521) );
  NAND2X1 U28812 ( .A(n73428), .B(n28845), .Y(n28844) );
  NAND2X1 U28814 ( .A(n44822), .B(n28813), .Y(n28843) );
  NAND2X1 U28815 ( .A(n28846), .B(n28847), .Y(n8520) );
  NAND2X1 U28816 ( .A(n73428), .B(n28848), .Y(n28847) );
  NAND2X1 U28852 ( .A(u_muldiv_invert_res_q), .B(n28813), .Y(n28846) );
  NAND2X1 U28913 ( .A(u_muldiv_rd_q[0]), .B(u_muldiv_div_busy_q), .Y(n28905)
         );
  NAND2X1 U28914 ( .A(n28907), .B(n28908), .Y(n8509) );
  NAND2X1 U28916 ( .A(u_muldiv_rd_q[1]), .B(u_muldiv_div_busy_q), .Y(n28907)
         );
  NAND2X1 U28917 ( .A(n28909), .B(n28910), .Y(n8508) );
  NAND2X1 U28919 ( .A(u_muldiv_rd_q[2]), .B(u_muldiv_div_busy_q), .Y(n28909)
         );
  NAND2X1 U28922 ( .A(u_muldiv_rd_q[3]), .B(u_muldiv_div_busy_q), .Y(n28911)
         );
  NAND2X1 U28928 ( .A(u_muldiv_rd_q[4]), .B(u_muldiv_div_busy_q), .Y(n28913)
         );
  NAND2X1 U28954 ( .A(n28932), .B(n28933), .Y(n8498) );
  OR2X1 U28955 ( .A(n28934), .B(n1883), .Y(n28933) );
  NAND2X1 U28969 ( .A(n28941), .B(n28942), .Y(n8496) );
  NAND2X1 U28970 ( .A(n28943), .B(n28934), .Y(n28942) );
  OR2X1 U28972 ( .A(n28934), .B(n1884), .Y(n28941) );
  NAND2X1 U28973 ( .A(n28944), .B(n28945), .Y(n8495) );
  NAND2X1 U28974 ( .A(n28946), .B(n28934), .Y(n28945) );
  OR2X1 U28976 ( .A(n28934), .B(n1885), .Y(n28944) );
  NAND2X1 U28977 ( .A(n28947), .B(n28948), .Y(n8494) );
  NAND2X1 U28978 ( .A(n28949), .B(n28934), .Y(n28948) );
  OR2X1 U28980 ( .A(n28934), .B(n1886), .Y(n28947) );
  NAND2X1 U29025 ( .A(u_mmu_dtlb_va_addr_q[25]), .B(n28953), .Y(n28982) );
  NAND2X1 U29046 ( .A(u_mmu_dtlb_va_addr_q[29]), .B(n28953), .Y(n28996) );
  NAND2X1 U29086 ( .A(n29026), .B(n29027), .Y(n17305) );
  NAND2X1 U29087 ( .A(challenge[97]), .B(n44854), .Y(n29026) );
  NAND2X1 U29088 ( .A(n29028), .B(n29027), .Y(n17304) );
  NAND2X1 U29089 ( .A(n29029), .B(n44862), .Y(n29027) );
  NAND2X1 U29090 ( .A(n29030), .B(n538), .Y(n29029) );
  NOR2X1 U29091 ( .A(n18691), .B(n18688), .Y(n29030) );
  NOR2X1 U29092 ( .A(n29031), .B(n29032), .Y(n18688) );
  NAND2X1 U29093 ( .A(n1062), .B(n538), .Y(n29031) );
  NOR2X1 U29094 ( .A(n29034), .B(n24252), .Y(n18691) );
  NAND2X1 U29095 ( .A(n29035), .B(n29036), .Y(n24252) );
  OR2X1 U29096 ( .A(n29037), .B(n29033), .Y(n29034) );
  NAND2X1 U29097 ( .A(n24256), .B(n44582), .Y(n29033) );
  NOR2X1 U29100 ( .A(n29040), .B(n29032), .Y(n29037) );
  NAND2X1 U29101 ( .A(challenge[96]), .B(n44854), .Y(n29028) );
  NAND2X1 U29102 ( .A(n29041), .B(n29042), .Y(n17303) );
  NAND2X1 U29103 ( .A(challenge[95]), .B(n44854), .Y(n29041) );
  NAND2X1 U29104 ( .A(n29043), .B(n29042), .Y(n17302) );
  NAND2X1 U29105 ( .A(n29044), .B(n44862), .Y(n29042) );
  NAND2X1 U29106 ( .A(n29045), .B(n546), .Y(n29044) );
  AND2X1 U29107 ( .A(n44348), .B(n44357), .Y(n29045) );
  NAND2X1 U29110 ( .A(n29036), .B(n29049), .Y(n24184) );
  OR2X1 U29111 ( .A(n29046), .B(n29047), .Y(n29048) );
  NAND2X1 U29112 ( .A(n24188), .B(n44351), .Y(n29047) );
  NOR2X1 U29115 ( .A(n29053), .B(n29032), .Y(n29046) );
  NAND2X1 U29116 ( .A(challenge[94]), .B(n44854), .Y(n29043) );
  NAND2X1 U29117 ( .A(n29054), .B(n29055), .Y(n17301) );
  NAND2X1 U29118 ( .A(challenge[93]), .B(n44854), .Y(n29054) );
  NAND2X1 U29119 ( .A(n29056), .B(n29055), .Y(n17300) );
  NAND2X1 U29120 ( .A(n29057), .B(n44861), .Y(n29055) );
  NAND2X1 U29121 ( .A(n29058), .B(n564), .Y(n29057) );
  AND2X1 U29122 ( .A(n44588), .B(n44597), .Y(n29058) );
  NOR2X1 U29124 ( .A(n29059), .B(n29061), .Y(n29060) );
  NAND2X1 U29126 ( .A(n29063), .B(n29036), .Y(n24243) );
  OR2X1 U29127 ( .A(n29064), .B(n29059), .Y(n29062) );
  NAND2X1 U29128 ( .A(n24247), .B(n44591), .Y(n29059) );
  NOR2X1 U29131 ( .A(n29061), .B(n29040), .Y(n29064) );
  NAND2X1 U29132 ( .A(challenge[92]), .B(n44854), .Y(n29056) );
  NAND2X1 U29133 ( .A(n29067), .B(n29068), .Y(n17299) );
  NAND2X1 U29134 ( .A(challenge[91]), .B(n44853), .Y(n29067) );
  NAND2X1 U29135 ( .A(n29069), .B(n29068), .Y(n17298) );
  NAND2X1 U29136 ( .A(n29070), .B(n44861), .Y(n29068) );
  NAND2X1 U29137 ( .A(n29071), .B(n550), .Y(n29070) );
  AND2X1 U29138 ( .A(n44336), .B(n44345), .Y(n29071) );
  NAND2X1 U29141 ( .A(n29075), .B(n29076), .Y(n24200) );
  OR2X1 U29142 ( .A(n29072), .B(n29073), .Y(n29074) );
  NAND2X1 U29143 ( .A(n24203), .B(n44339), .Y(n29073) );
  NOR2X1 U29145 ( .A(n29053), .B(n29079), .Y(n29072) );
  NAND2X1 U29146 ( .A(challenge[90]), .B(n44853), .Y(n29069) );
  NAND2X1 U29147 ( .A(n29080), .B(n29081), .Y(n17297) );
  NAND2X1 U29148 ( .A(challenge[89]), .B(n44853), .Y(n29080) );
  NAND2X1 U29149 ( .A(n29082), .B(n29081), .Y(n17296) );
  NAND2X1 U29150 ( .A(n29083), .B(n44861), .Y(n29081) );
  NAND2X1 U29151 ( .A(n29084), .B(n523), .Y(n29083) );
  NOR2X1 U29152 ( .A(n18299), .B(n18295), .Y(n29084) );
  NOR2X1 U29153 ( .A(n29086), .B(n29087), .Y(n18295) );
  OR2X1 U29154 ( .A(n29053), .B(n29085), .Y(n29086) );
  NOR2X1 U29155 ( .A(n29088), .B(n24235), .Y(n18299) );
  NAND2X1 U29156 ( .A(n29049), .B(n29089), .Y(n24235) );
  OR2X1 U29157 ( .A(n29090), .B(n29085), .Y(n29088) );
  NAND2X1 U29158 ( .A(n18296), .B(n44600), .Y(n29085) );
  NOR2X1 U29160 ( .A(n29053), .B(n29087), .Y(n29090) );
  NAND2X1 U29161 ( .A(challenge[88]), .B(n44853), .Y(n29082) );
  NAND2X1 U29162 ( .A(n29093), .B(n29094), .Y(n17295) );
  NAND2X1 U29163 ( .A(challenge[87]), .B(n44853), .Y(n29093) );
  NAND2X1 U29164 ( .A(n29095), .B(n29094), .Y(n17294) );
  NAND2X1 U29165 ( .A(n29096), .B(n44860), .Y(n29094) );
  NAND2X1 U29166 ( .A(n29097), .B(n548), .Y(n29096) );
  AND2X1 U29167 ( .A(n44324), .B(n44333), .Y(n29097) );
  NAND2X1 U29170 ( .A(n29075), .B(n29049), .Y(n24207) );
  OR2X1 U29171 ( .A(n29098), .B(n29099), .Y(n29100) );
  NAND2X1 U29172 ( .A(n24210), .B(n44327), .Y(n29099) );
  NOR2X1 U29175 ( .A(n29053), .B(n29101), .Y(n29098) );
  NAND2X1 U29176 ( .A(challenge[86]), .B(n44853), .Y(n29095) );
  NAND2X1 U29177 ( .A(n29102), .B(n29103), .Y(n17293) );
  NAND2X1 U29178 ( .A(challenge[85]), .B(n44853), .Y(n29102) );
  NAND2X1 U29179 ( .A(n29104), .B(n29103), .Y(n17292) );
  NAND2X1 U29180 ( .A(n29105), .B(n44860), .Y(n29103) );
  NAND2X1 U29181 ( .A(n29106), .B(n517), .Y(n29105) );
  NOR2X1 U29182 ( .A(n24104), .B(n24100), .Y(n29106) );
  NOR2X1 U29183 ( .A(n29108), .B(n29109), .Y(n24100) );
  OR2X1 U29184 ( .A(n29107), .B(n29053), .Y(n29108) );
  NOR2X1 U29185 ( .A(n29110), .B(n24228), .Y(n24104) );
  NAND2X1 U29186 ( .A(n29076), .B(n29089), .Y(n24228) );
  OR2X1 U29187 ( .A(n29111), .B(n29107), .Y(n29110) );
  NAND2X1 U29188 ( .A(n24101), .B(n44606), .Y(n29107) );
  NOR2X1 U29191 ( .A(n29053), .B(n29109), .Y(n29111) );
  NAND2X1 U29192 ( .A(challenge[84]), .B(n44853), .Y(n29104) );
  NAND2X1 U29193 ( .A(n29112), .B(n29113), .Y(n17291) );
  NAND2X1 U29194 ( .A(challenge[83]), .B(n44853), .Y(n29112) );
  NAND2X1 U29195 ( .A(n29114), .B(n29113), .Y(n17290) );
  NAND2X1 U29196 ( .A(n29115), .B(n44860), .Y(n29113) );
  NAND2X1 U29197 ( .A(n29116), .B(n551), .Y(n29115) );
  AND2X1 U29198 ( .A(n44312), .B(n44321), .Y(n29116) );
  NAND2X1 U29201 ( .A(n29120), .B(n29076), .Y(n24214) );
  OR2X1 U29202 ( .A(n29117), .B(n29118), .Y(n29119) );
  NAND2X1 U29203 ( .A(n24217), .B(n44315), .Y(n29118) );
  NOR2X1 U29205 ( .A(n29053), .B(n29122), .Y(n29117) );
  NAND2X1 U29206 ( .A(challenge[82]), .B(n44853), .Y(n29114) );
  NAND2X1 U29207 ( .A(n29123), .B(n29124), .Y(n17289) );
  NAND2X1 U29208 ( .A(challenge[81]), .B(n44853), .Y(n29123) );
  NAND2X1 U29209 ( .A(n29125), .B(n29124), .Y(n17288) );
  NAND2X1 U29210 ( .A(n29126), .B(n44857), .Y(n29124) );
  NAND2X1 U29211 ( .A(n29127), .B(n544), .Y(n29126) );
  AND2X1 U29212 ( .A(n44300), .B(n44309), .Y(n29127) );
  NAND2X1 U29215 ( .A(n29120), .B(n29049), .Y(n24221) );
  OR2X1 U29216 ( .A(n29128), .B(n29129), .Y(n29130) );
  NAND2X1 U29217 ( .A(n24224), .B(n44303), .Y(n29129) );
  NOR2X1 U29220 ( .A(n29053), .B(n29132), .Y(n29128) );
  NAND2X1 U29221 ( .A(challenge[80]), .B(n44853), .Y(n29125) );
  NAND2X1 U29222 ( .A(n29133), .B(n29134), .Y(n17287) );
  NAND2X1 U29223 ( .A(challenge[79]), .B(n44852), .Y(n29133) );
  NAND2X1 U29224 ( .A(n29135), .B(n29134), .Y(n17286) );
  NAND2X1 U29225 ( .A(n29136), .B(n44863), .Y(n29134) );
  NAND2X1 U29226 ( .A(n29137), .B(n554), .Y(n29136) );
  AND2X1 U29227 ( .A(n44360), .B(n44369), .Y(n29137) );
  NAND2X1 U29230 ( .A(n29036), .B(n29076), .Y(n24175) );
  AND2X1 U29231 ( .A(n29141), .B(writeback_muldiv_idx_w[2]), .Y(n29036) );
  NOR2X1 U29232 ( .A(n37339), .B(n37541), .Y(n29141) );
  OR2X1 U29233 ( .A(n29138), .B(n29139), .Y(n29140) );
  NAND2X1 U29234 ( .A(n24179), .B(n44363), .Y(n29139) );
  NOR2X1 U29237 ( .A(n29053), .B(n29061), .Y(n29138) );
  NAND2X1 U29238 ( .A(n37482), .B(n29144), .Y(n29053) );
  NAND2X1 U29239 ( .A(challenge[78]), .B(n44852), .Y(n29135) );
  NAND2X1 U29240 ( .A(n29145), .B(n29146), .Y(n17285) );
  NAND2X1 U29241 ( .A(challenge[77]), .B(n44852), .Y(n29145) );
  NAND2X1 U29242 ( .A(n29147), .B(n29146), .Y(n17284) );
  NAND2X1 U29243 ( .A(n29148), .B(n44856), .Y(n29146) );
  NAND2X1 U29244 ( .A(n29149), .B(n37472), .Y(n29148) );
  AND2X1 U29245 ( .A(n44372), .B(n44375), .Y(n29149) );
  NOR2X1 U29247 ( .A(n29152), .B(n24274), .Y(n29151) );
  NAND2X1 U29248 ( .A(n29153), .B(n29063), .Y(n24274) );
  NOR2X1 U29252 ( .A(n29109), .B(n1065), .Y(n29152) );
  NAND2X1 U29253 ( .A(challenge[76]), .B(n44852), .Y(n29147) );
  NAND2X1 U29254 ( .A(n29156), .B(n29157), .Y(n17283) );
  NAND2X1 U29255 ( .A(challenge[75]), .B(n44852), .Y(n29156) );
  NAND2X1 U29256 ( .A(n29158), .B(n29157), .Y(n17282) );
  NAND2X1 U29257 ( .A(n29159), .B(n44859), .Y(n29157) );
  NAND2X1 U29258 ( .A(n29160), .B(n526), .Y(n29159) );
  AND2X1 U29259 ( .A(n44378), .B(n44387), .Y(n29160) );
  NAND2X1 U29262 ( .A(n29164), .B(n29035), .Y(n24192) );
  OR2X1 U29263 ( .A(n29161), .B(n29162), .Y(n29163) );
  NAND2X1 U29264 ( .A(n24196), .B(n44381), .Y(n29162) );
  NOR2X1 U29266 ( .A(n29132), .B(n1065), .Y(n29161) );
  NAND2X1 U29267 ( .A(challenge[74]), .B(n44852), .Y(n29158) );
  NAND2X1 U29268 ( .A(n29167), .B(n29168), .Y(n17281) );
  NAND2X1 U29269 ( .A(challenge[73]), .B(n44852), .Y(n29167) );
  NAND2X1 U29270 ( .A(n29169), .B(n29168), .Y(n17280) );
  NAND2X1 U29271 ( .A(n29170), .B(n44859), .Y(n29168) );
  NAND2X1 U29272 ( .A(n29171), .B(n566), .Y(n29170) );
  AND2X1 U29273 ( .A(n44390), .B(n44399), .Y(n29171) );
  NAND2X1 U29276 ( .A(n29164), .B(n29063), .Y(n24166) );
  OR2X1 U29277 ( .A(n29172), .B(n29173), .Y(n29174) );
  NAND2X1 U29278 ( .A(n24170), .B(n44393), .Y(n29173) );
  NOR2X1 U29281 ( .A(n29122), .B(n1065), .Y(n29172) );
  NAND2X1 U29282 ( .A(challenge[72]), .B(n44852), .Y(n29169) );
  NAND2X1 U29283 ( .A(n29176), .B(n29177), .Y(n17279) );
  NAND2X1 U29284 ( .A(challenge[71]), .B(n44852), .Y(n29176) );
  NAND2X1 U29285 ( .A(n29178), .B(n29177), .Y(n17278) );
  NAND2X1 U29286 ( .A(n29179), .B(n44859), .Y(n29177) );
  NAND2X1 U29287 ( .A(n29180), .B(n528), .Y(n29179) );
  AND2X1 U29288 ( .A(n44402), .B(n44411), .Y(n29180) );
  NAND2X1 U29291 ( .A(n29184), .B(n29035), .Y(n24158) );
  OR2X1 U29292 ( .A(n29181), .B(n29182), .Y(n29183) );
  NAND2X1 U29293 ( .A(n24161), .B(n44405), .Y(n29182) );
  NOR2X1 U29296 ( .A(n29101), .B(n1065), .Y(n29181) );
  NAND2X1 U29297 ( .A(challenge[70]), .B(n44852), .Y(n29178) );
  NAND2X1 U29298 ( .A(n29187), .B(n29188), .Y(n17277) );
  NAND2X1 U29299 ( .A(challenge[69]), .B(n44852), .Y(n29187) );
  NAND2X1 U29300 ( .A(n29189), .B(n29188), .Y(n17276) );
  NAND2X1 U29301 ( .A(n29190), .B(n44862), .Y(n29188) );
  NAND2X1 U29302 ( .A(n29191), .B(n572), .Y(n29190) );
  AND2X1 U29303 ( .A(n44414), .B(n44423), .Y(n29191) );
  NAND2X1 U29306 ( .A(n29184), .B(n29063), .Y(n24149) );
  OR2X1 U29307 ( .A(n29192), .B(n29193), .Y(n29194) );
  NAND2X1 U29308 ( .A(n24153), .B(n44417), .Y(n29193) );
  NOR2X1 U29311 ( .A(n29079), .B(n1065), .Y(n29192) );
  NAND2X1 U29312 ( .A(challenge[68]), .B(n44852), .Y(n29189) );
  NAND2X1 U29313 ( .A(n29197), .B(n29198), .Y(n17275) );
  NAND2X1 U29314 ( .A(challenge[67]), .B(wm_select), .Y(n29197) );
  NAND2X1 U29315 ( .A(n29199), .B(n29198), .Y(n17274) );
  NAND2X1 U29316 ( .A(n29200), .B(n44861), .Y(n29198) );
  NAND2X1 U29317 ( .A(n29201), .B(n530), .Y(n29200) );
  AND2X1 U29318 ( .A(n44426), .B(n44435), .Y(n29201) );
  NAND2X1 U29321 ( .A(n29205), .B(n29035), .Y(n24140) );
  OR2X1 U29322 ( .A(n29202), .B(n29203), .Y(n29204) );
  NAND2X1 U29323 ( .A(n24144), .B(n44429), .Y(n29203) );
  NOR2X1 U29325 ( .A(n29032), .B(n1065), .Y(n29202) );
  NAND2X1 U29326 ( .A(challenge[66]), .B(wm_select), .Y(n29199) );
  NAND2X1 U29327 ( .A(n29207), .B(n29208), .Y(n17273) );
  NAND2X1 U29328 ( .A(challenge[65]), .B(n44846), .Y(n29207) );
  NAND2X1 U29329 ( .A(n29209), .B(n29208), .Y(n17272) );
  NAND2X1 U29330 ( .A(n29210), .B(n44857), .Y(n29208) );
  NAND2X1 U29331 ( .A(n29211), .B(n570), .Y(n29210) );
  AND2X1 U29332 ( .A(n44438), .B(n44447), .Y(n29211) );
  NOR2X1 U29334 ( .A(n29061), .B(n29212), .Y(n29213) );
  NAND2X1 U29336 ( .A(n29205), .B(n29063), .Y(n24129) );
  OR2X1 U29337 ( .A(n29216), .B(n29212), .Y(n29215) );
  NAND2X1 U29338 ( .A(n24134), .B(n44441), .Y(n29212) );
  NOR2X1 U29341 ( .A(n29061), .B(n1065), .Y(n29216) );
  NOR2X1 U29342 ( .A(n29144), .B(n37482), .Y(n29214) );
  NAND2X1 U29343 ( .A(challenge[64]), .B(wm_select), .Y(n29209) );
  NAND2X1 U29344 ( .A(n29217), .B(n29218), .Y(n17271) );
  NAND2X1 U29345 ( .A(challenge[63]), .B(wm_select), .Y(n29217) );
  NAND2X1 U29346 ( .A(n29219), .B(n29218), .Y(n17270) );
  NAND2X1 U29347 ( .A(n29220), .B(n44858), .Y(n29218) );
  NAND2X1 U29348 ( .A(n29221), .B(n73406), .Y(n29220) );
  AND2X1 U29349 ( .A(n44450), .B(n44453), .Y(n29221) );
  NAND2X1 U29352 ( .A(n29153), .B(n29049), .Y(n24122) );
  OR2X1 U29353 ( .A(n29222), .B(n29223), .Y(n29224) );
  NOR2X1 U29356 ( .A(n29087), .B(n1063), .Y(n29222) );
  NAND2X1 U29357 ( .A(challenge[62]), .B(n44846), .Y(n29219) );
  NAND2X1 U29358 ( .A(n29225), .B(n29226), .Y(n17269) );
  NAND2X1 U29359 ( .A(challenge[61]), .B(wm_select), .Y(n29225) );
  NAND2X1 U29360 ( .A(n29227), .B(n29226), .Y(n17268) );
  NAND2X1 U29361 ( .A(n29228), .B(n44858), .Y(n29226) );
  NAND2X1 U29362 ( .A(n29229), .B(n491), .Y(n29228) );
  AND2X1 U29363 ( .A(n44456), .B(n44465), .Y(n29229) );
  NAND2X1 U29366 ( .A(n29153), .B(n29076), .Y(n24115) );
  AND2X1 U29367 ( .A(n29233), .B(n37541), .Y(n29153) );
  OR2X1 U29368 ( .A(n29230), .B(n29231), .Y(n29232) );
  NAND2X1 U29369 ( .A(n21240), .B(n44459), .Y(n29231) );
  NOR2X1 U29372 ( .A(n29109), .B(n1063), .Y(n29230) );
  NAND2X1 U29373 ( .A(challenge[60]), .B(n44846), .Y(n29227) );
  NAND2X1 U29374 ( .A(n29234), .B(n29235), .Y(n17267) );
  NAND2X1 U29375 ( .A(challenge[59]), .B(wm_select), .Y(n29234) );
  NAND2X1 U29376 ( .A(n29236), .B(n29235), .Y(n17266) );
  NAND2X1 U29377 ( .A(n29237), .B(n44860), .Y(n29235) );
  NAND2X1 U29378 ( .A(n29238), .B(n502), .Y(n29237) );
  AND2X1 U29379 ( .A(n44468), .B(n44477), .Y(n29238) );
  NAND2X1 U29382 ( .A(n29164), .B(n29049), .Y(n24357) );
  OR2X1 U29383 ( .A(n29239), .B(n29240), .Y(n29241) );
  NAND2X1 U29384 ( .A(n24361), .B(n44471), .Y(n29240) );
  NOR2X1 U29386 ( .A(n29132), .B(n1063), .Y(n29239) );
  NAND2X1 U29387 ( .A(challenge[58]), .B(n44846), .Y(n29236) );
  NAND2X1 U29388 ( .A(n29242), .B(n29243), .Y(n17265) );
  NAND2X1 U29389 ( .A(challenge[57]), .B(wm_select), .Y(n29242) );
  NAND2X1 U29390 ( .A(n29244), .B(n29243), .Y(n17264) );
  NAND2X1 U29391 ( .A(n29245), .B(n44859), .Y(n29243) );
  NAND2X1 U29392 ( .A(n29246), .B(n494), .Y(n29245) );
  AND2X1 U29393 ( .A(n44480), .B(n44489), .Y(n29246) );
  NAND2X1 U29396 ( .A(n29164), .B(n29076), .Y(n24349) );
  AND2X1 U29397 ( .A(n29233), .B(writeback_muldiv_idx_w[1]), .Y(n29164) );
  NOR2X1 U29398 ( .A(writeback_muldiv_idx_w[4]), .B(writeback_muldiv_idx_w[2]), 
        .Y(n29233) );
  OR2X1 U29399 ( .A(n29247), .B(n29248), .Y(n29249) );
  NAND2X1 U29400 ( .A(n24353), .B(n44483), .Y(n29248) );
  NOR2X1 U29403 ( .A(n29122), .B(n1063), .Y(n29247) );
  NAND2X1 U29404 ( .A(challenge[56]), .B(n44851), .Y(n29244) );
  NAND2X1 U29405 ( .A(n29250), .B(n29251), .Y(n17263) );
  NAND2X1 U29406 ( .A(challenge[55]), .B(n44851), .Y(n29250) );
  NAND2X1 U29407 ( .A(n29252), .B(n29251), .Y(n17262) );
  NAND2X1 U29408 ( .A(n29253), .B(n44859), .Y(n29251) );
  NAND2X1 U29409 ( .A(n29254), .B(n73407), .Y(n29253) );
  AND2X1 U29410 ( .A(n44492), .B(n44495), .Y(n29254) );
  NAND2X1 U29413 ( .A(n29184), .B(n29049), .Y(n24341) );
  OR2X1 U29414 ( .A(n29255), .B(n29256), .Y(n29257) );
  NOR2X1 U29417 ( .A(n29101), .B(n1063), .Y(n29255) );
  NAND2X1 U29418 ( .A(challenge[54]), .B(n44851), .Y(n29252) );
  NAND2X1 U29419 ( .A(n29258), .B(n29259), .Y(n17261) );
  NAND2X1 U29420 ( .A(challenge[53]), .B(n44851), .Y(n29258) );
  NAND2X1 U29421 ( .A(n29260), .B(n29259), .Y(n17260) );
  NAND2X1 U29422 ( .A(n29261), .B(n44858), .Y(n29259) );
  NAND2X1 U29423 ( .A(n29262), .B(n498), .Y(n29261) );
  AND2X1 U29424 ( .A(n44498), .B(n44507), .Y(n29262) );
  NAND2X1 U29427 ( .A(n29184), .B(n29076), .Y(n24333) );
  AND2X1 U29428 ( .A(n29266), .B(writeback_muldiv_idx_w[2]), .Y(n29184) );
  NOR2X1 U29429 ( .A(writeback_muldiv_idx_w[4]), .B(writeback_muldiv_idx_w[1]), 
        .Y(n29266) );
  OR2X1 U29430 ( .A(n29263), .B(n29264), .Y(n29265) );
  NAND2X1 U29431 ( .A(n24336), .B(n44501), .Y(n29264) );
  NOR2X1 U29434 ( .A(n29079), .B(n1063), .Y(n29263) );
  NAND2X1 U29435 ( .A(challenge[52]), .B(n44851), .Y(n29260) );
  NAND2X1 U29436 ( .A(n29267), .B(n29268), .Y(n17259) );
  NAND2X1 U29437 ( .A(challenge[51]), .B(n44851), .Y(n29267) );
  NAND2X1 U29438 ( .A(n29269), .B(n29268), .Y(n17258) );
  NAND2X1 U29439 ( .A(n29270), .B(n44847), .Y(n29268) );
  NAND2X1 U29440 ( .A(n29271), .B(n504), .Y(n29270) );
  AND2X1 U29441 ( .A(n44510), .B(n44519), .Y(n29271) );
  NAND2X1 U29444 ( .A(n29205), .B(n29049), .Y(n24323) );
  NOR2X1 U29445 ( .A(n37542), .B(writeback_muldiv_idx_w[0]), .Y(n29049) );
  OR2X1 U29446 ( .A(n29272), .B(n29273), .Y(n29274) );
  NAND2X1 U29447 ( .A(n24328), .B(n44513), .Y(n29273) );
  NOR2X1 U29450 ( .A(n29032), .B(n1063), .Y(n29272) );
  NAND2X1 U29451 ( .A(n37337), .B(n29275), .Y(n29032) );
  NAND2X1 U29452 ( .A(challenge[50]), .B(n44851), .Y(n29269) );
  NAND2X1 U29453 ( .A(n29276), .B(n29277), .Y(n17257) );
  NAND2X1 U29454 ( .A(challenge[49]), .B(n44851), .Y(n29276) );
  NAND2X1 U29455 ( .A(n29278), .B(n29277), .Y(n17256) );
  NAND2X1 U29456 ( .A(n29279), .B(n44858), .Y(n29277) );
  NAND2X1 U29457 ( .A(n29280), .B(n496), .Y(n29279) );
  AND2X1 U29458 ( .A(n44522), .B(n44531), .Y(n29280) );
  NOR2X1 U29460 ( .A(n29061), .B(n29281), .Y(n29282) );
  NAND2X1 U29462 ( .A(n29205), .B(n29076), .Y(n24312) );
  NOR2X1 U29463 ( .A(n37542), .B(n37338), .Y(n29076) );
  AND2X1 U29464 ( .A(n29285), .B(writeback_muldiv_idx_w[2]), .Y(n29205) );
  NOR2X1 U29465 ( .A(writeback_muldiv_idx_w[4]), .B(n37541), .Y(n29285) );
  OR2X1 U29466 ( .A(n29286), .B(n29281), .Y(n29284) );
  NAND2X1 U29467 ( .A(n24316), .B(n44525), .Y(n29281) );
  NOR2X1 U29472 ( .A(n29061), .B(n1063), .Y(n29286) );
  NOR2X1 U29473 ( .A(n1064), .B(n37482), .Y(n29283) );
  NAND2X1 U29474 ( .A(n29287), .B(u_csr_writeback_idx_q[1]), .Y(n29061) );
  NOR2X1 U29475 ( .A(n1053), .B(n1057), .Y(n29287) );
  NAND2X1 U29476 ( .A(challenge[48]), .B(n44851), .Y(n29278) );
  NAND2X1 U29477 ( .A(n29288), .B(n29289), .Y(n17255) );
  NAND2X1 U29478 ( .A(challenge[47]), .B(n44851), .Y(n29288) );
  NAND2X1 U29479 ( .A(n29290), .B(n29289), .Y(n17254) );
  NAND2X1 U29480 ( .A(n29291), .B(n44847), .Y(n29289) );
  NAND2X1 U29481 ( .A(n29292), .B(n512), .Y(n29291) );
  AND2X1 U29482 ( .A(n44534), .B(n44543), .Y(n29292) );
  NAND2X1 U29485 ( .A(n29035), .B(n29089), .Y(n24302) );
  OR2X1 U29486 ( .A(n29293), .B(n29294), .Y(n29295) );
  NAND2X1 U29487 ( .A(n19867), .B(n44537), .Y(n29294) );
  NOR2X1 U29490 ( .A(n29087), .B(n29040), .Y(n29293) );
  NAND2X1 U29491 ( .A(n36767), .B(n1057), .Y(n29087) );
  NAND2X1 U29492 ( .A(challenge[46]), .B(n44851), .Y(n29290) );
  NAND2X1 U29493 ( .A(n29298), .B(n29299), .Y(n17253) );
  NAND2X1 U29494 ( .A(challenge[45]), .B(n44851), .Y(n29298) );
  NAND2X1 U29495 ( .A(n29300), .B(n29299), .Y(n17252) );
  NAND2X1 U29496 ( .A(n29301), .B(n44863), .Y(n29299) );
  NAND2X1 U29497 ( .A(n29302), .B(n519), .Y(n29301) );
  AND2X1 U29498 ( .A(n44546), .B(n44555), .Y(n29302) );
  NAND2X1 U29501 ( .A(n29063), .B(n29089), .Y(n24294) );
  AND2X1 U29502 ( .A(n29306), .B(n37541), .Y(n29089) );
  OR2X1 U29503 ( .A(n29303), .B(n29304), .Y(n29305) );
  NAND2X1 U29504 ( .A(n19670), .B(n44549), .Y(n29304) );
  NOR2X1 U29507 ( .A(n29109), .B(n29040), .Y(n29303) );
  NAND2X1 U29508 ( .A(n29308), .B(n29309), .Y(n29109) );
  NOR2X1 U29509 ( .A(u_csr_writeback_idx_q[1]), .B(n29275), .Y(n29308) );
  NAND2X1 U29510 ( .A(challenge[44]), .B(n44850), .Y(n29300) );
  NAND2X1 U29511 ( .A(n29310), .B(n29311), .Y(n17251) );
  NAND2X1 U29512 ( .A(challenge[43]), .B(n44850), .Y(n29310) );
  NAND2X1 U29513 ( .A(n29312), .B(n29311), .Y(n17250) );
  NAND2X1 U29514 ( .A(n29313), .B(n44862), .Y(n29311) );
  NAND2X1 U29515 ( .A(n29314), .B(n542), .Y(n29313) );
  NOR2X1 U29516 ( .A(n19475), .B(n19472), .Y(n29314) );
  NOR2X1 U29517 ( .A(n29315), .B(n29132), .Y(n19472) );
  NAND2X1 U29518 ( .A(n1062), .B(n542), .Y(n29315) );
  NOR2X1 U29519 ( .A(n29317), .B(n24287), .Y(n19475) );
  NAND2X1 U29520 ( .A(n29120), .B(n29035), .Y(n24287) );
  OR2X1 U29521 ( .A(n29318), .B(n29316), .Y(n29317) );
  NAND2X1 U29522 ( .A(n24290), .B(n44558), .Y(n29316) );
  NOR2X1 U29526 ( .A(n29040), .B(n29132), .Y(n29318) );
  NAND2X1 U29527 ( .A(n29320), .B(n37337), .Y(n29132) );
  NOR2X1 U29529 ( .A(n29275), .B(n29321), .Y(n29320) );
  NAND2X1 U29530 ( .A(challenge[42]), .B(n44850), .Y(n29312) );
  NAND2X1 U29531 ( .A(n29322), .B(n29323), .Y(n17249) );
  NAND2X1 U29532 ( .A(challenge[41]), .B(n44850), .Y(n29322) );
  NAND2X1 U29533 ( .A(n29324), .B(n29323), .Y(n17248) );
  NAND2X1 U29534 ( .A(n29325), .B(n44860), .Y(n29323) );
  NAND2X1 U29535 ( .A(n29326), .B(n562), .Y(n29325) );
  NOR2X1 U29536 ( .A(n19279), .B(n19276), .Y(n29326) );
  NOR2X1 U29537 ( .A(n29327), .B(n29122), .Y(n19276) );
  NAND2X1 U29538 ( .A(n1062), .B(n562), .Y(n29327) );
  NOR2X1 U29539 ( .A(n29329), .B(n24280), .Y(n19279) );
  NAND2X1 U29540 ( .A(n29120), .B(n29063), .Y(n24280) );
  AND2X1 U29541 ( .A(writeback_muldiv_idx_w[1]), .B(n29306), .Y(n29120) );
  NOR2X1 U29542 ( .A(n37339), .B(writeback_muldiv_idx_w[2]), .Y(n29306) );
  OR2X1 U29543 ( .A(n29330), .B(n29328), .Y(n29329) );
  NAND2X1 U29544 ( .A(n24283), .B(n44564), .Y(n29328) );
  NOR2X1 U29548 ( .A(n29040), .B(n29122), .Y(n29330) );
  NAND2X1 U29549 ( .A(n29332), .B(u_csr_writeback_idx_q[1]), .Y(n29122) );
  NOR2X1 U29550 ( .A(n29275), .B(n1053), .Y(n29332) );
  NAND2X1 U29551 ( .A(challenge[40]), .B(n44850), .Y(n29324) );
  NAND2X1 U29552 ( .A(n29333), .B(n29334), .Y(n17247) );
  NAND2X1 U29553 ( .A(challenge[39]), .B(n44850), .Y(n29333) );
  NAND2X1 U29554 ( .A(n29335), .B(n29334), .Y(n17246) );
  NAND2X1 U29555 ( .A(n29336), .B(n44857), .Y(n29334) );
  NAND2X1 U29556 ( .A(n29337), .B(n534), .Y(n29336) );
  NOR2X1 U29557 ( .A(n19083), .B(n19080), .Y(n29337) );
  NOR2X1 U29558 ( .A(n29338), .B(n29101), .Y(n19080) );
  NAND2X1 U29559 ( .A(n1062), .B(n534), .Y(n29338) );
  NOR2X1 U29560 ( .A(n29340), .B(n24267), .Y(n19083) );
  NAND2X1 U29561 ( .A(n29075), .B(n29035), .Y(n24267) );
  NOR2X1 U29562 ( .A(writeback_muldiv_idx_w[0]), .B(writeback_muldiv_idx_w[3]), 
        .Y(n29035) );
  OR2X1 U29563 ( .A(n29341), .B(n29339), .Y(n29340) );
  NAND2X1 U29564 ( .A(n24270), .B(n44570), .Y(n29339) );
  NOR2X1 U29567 ( .A(n29040), .B(n29101), .Y(n29341) );
  NAND2X1 U29568 ( .A(n29275), .B(n36767), .Y(n29101) );
  NAND2X1 U29570 ( .A(challenge[38]), .B(n44850), .Y(n29335) );
  NAND2X1 U29571 ( .A(n29343), .B(n29344), .Y(n17245) );
  NAND2X1 U29572 ( .A(challenge[37]), .B(n44850), .Y(n29343) );
  NAND2X1 U29573 ( .A(n29345), .B(n29344), .Y(n17244) );
  NAND2X1 U29574 ( .A(n29346), .B(n44859), .Y(n29344) );
  NAND2X1 U29575 ( .A(n29347), .B(n558), .Y(n29346) );
  NOR2X1 U29576 ( .A(n18887), .B(n18884), .Y(n29347) );
  NOR2X1 U29577 ( .A(n29348), .B(n29079), .Y(n18884) );
  NAND2X1 U29578 ( .A(n1062), .B(n558), .Y(n29348) );
  NOR2X1 U29579 ( .A(n29350), .B(n24260), .Y(n18887) );
  NAND2X1 U29580 ( .A(n29075), .B(n29063), .Y(n24260) );
  NOR2X1 U29581 ( .A(n37338), .B(writeback_muldiv_idx_w[3]), .Y(n29063) );
  AND2X1 U29582 ( .A(n29351), .B(writeback_muldiv_idx_w[2]), .Y(n29075) );
  NOR2X1 U29583 ( .A(writeback_muldiv_idx_w[1]), .B(n37339), .Y(n29351) );
  OR2X1 U29584 ( .A(n29352), .B(n29349), .Y(n29350) );
  NAND2X1 U29585 ( .A(n24263), .B(n44576), .Y(n29349) );
  NOR2X1 U29590 ( .A(n29040), .B(n29079), .Y(n29352) );
  NAND2X1 U29591 ( .A(n29354), .B(n29275), .Y(n29079) );
  NOR2X1 U29592 ( .A(n37483), .B(n29321), .Y(n29275) );
  NOR2X1 U29593 ( .A(u_csr_writeback_idx_q[1]), .B(n1053), .Y(n29354) );
  NAND2X1 U29595 ( .A(n37482), .B(n1064), .Y(n29040) );
  NAND2X1 U29599 ( .A(challenge[36]), .B(n44850), .Y(n29345) );
  NAND2X1 U29626 ( .A(n29371), .B(n29372), .Y(n17236) );
  NAND2X1 U29627 ( .A(challenge[28]), .B(n44850), .Y(n29371) );
  NAND2X1 U29628 ( .A(n29373), .B(n29372), .Y(n17235) );
  NAND2X1 U29629 ( .A(challenge[27]), .B(n44850), .Y(n29373) );
  NAND2X1 U29630 ( .A(n29374), .B(n29372), .Y(n17234) );
  NAND2X1 U29631 ( .A(challenge[26]), .B(n44850), .Y(n29374) );
  NAND2X1 U29632 ( .A(n29375), .B(n29372), .Y(n17233) );
  NAND2X1 U29633 ( .A(n29376), .B(n44861), .Y(n29372) );
  NAND2X1 U29634 ( .A(n28813), .B(n29377), .Y(n29376) );
  NAND2X1 U29635 ( .A(n29378), .B(n29379), .Y(n29377) );
  NOR2X1 U29636 ( .A(n29380), .B(n29381), .Y(n29379) );
  NAND2X1 U29637 ( .A(n29382), .B(n29383), .Y(n29381) );
  NOR2X1 U29638 ( .A(n29384), .B(n29385), .Y(n29383) );
  OR2X1 U29639 ( .A(u_muldiv_divisor_q[50]), .B(u_muldiv_divisor_q[51]), .Y(
        n29385) );
  OR2X1 U29640 ( .A(u_muldiv_divisor_q[52]), .B(u_muldiv_divisor_q[53]), .Y(
        n29384) );
  NOR2X1 U29641 ( .A(n29386), .B(n29387), .Y(n29382) );
  OR2X1 U29642 ( .A(u_muldiv_divisor_q[46]), .B(u_muldiv_divisor_q[47]), .Y(
        n29387) );
  OR2X1 U29643 ( .A(u_muldiv_divisor_q[48]), .B(u_muldiv_divisor_q[49]), .Y(
        n29386) );
  NAND2X1 U29644 ( .A(n29388), .B(n29389), .Y(n29380) );
  NOR2X1 U29645 ( .A(n29390), .B(n29391), .Y(n29389) );
  OR2X1 U29646 ( .A(u_muldiv_divisor_q[58]), .B(u_muldiv_divisor_q[59]), .Y(
        n29391) );
  NAND2X1 U29647 ( .A(n29392), .B(n1629), .Y(n29390) );
  NOR2X1 U29648 ( .A(u_muldiv_divisor_q[62]), .B(u_muldiv_divisor_q[61]), .Y(
        n29392) );
  NOR2X1 U29649 ( .A(n29393), .B(n29394), .Y(n29388) );
  OR2X1 U29650 ( .A(u_muldiv_divisor_q[54]), .B(u_muldiv_divisor_q[55]), .Y(
        n29394) );
  OR2X1 U29651 ( .A(u_muldiv_divisor_q[56]), .B(u_muldiv_divisor_q[57]), .Y(
        n29393) );
  NOR2X1 U29652 ( .A(n29395), .B(n29396), .Y(n29378) );
  NAND2X1 U29653 ( .A(n29397), .B(n29398), .Y(n29396) );
  NOR2X1 U29654 ( .A(n29399), .B(n29400), .Y(n29398) );
  OR2X1 U29655 ( .A(u_muldiv_divisor_q[33]), .B(u_muldiv_divisor_q[34]), .Y(
        n29400) );
  OR2X1 U29656 ( .A(u_muldiv_divisor_q[35]), .B(u_muldiv_divisor_q[36]), .Y(
        n29399) );
  NOR2X1 U29657 ( .A(n29401), .B(n29402), .Y(n29397) );
  NAND2X1 U29658 ( .A(n44612), .B(n29403), .Y(n29402) );
  OR2X1 U29659 ( .A(n29404), .B(u_muldiv_dividend_q[31]), .Y(n29403) );
  NAND2X1 U29660 ( .A(n29405), .B(n37591), .Y(n29401) );
  NAND2X1 U29661 ( .A(u_muldiv_divisor_q[31]), .B(n29406), .Y(n29405) );
  NAND2X1 U29662 ( .A(u_muldiv_dividend_q[31]), .B(n29404), .Y(n29406) );
  NAND2X1 U29663 ( .A(n14474), .B(n29407), .Y(n29404) );
  NAND2X1 U29664 ( .A(n29408), .B(n29409), .Y(n29407) );
  NAND2X1 U29665 ( .A(n29410), .B(n1630), .Y(n29409) );
  NOR2X1 U29666 ( .A(n14461), .B(n29411), .Y(n29408) );
  NOR2X1 U29667 ( .A(n29412), .B(n37583), .Y(n29411) );
  NOR2X1 U29668 ( .A(n29410), .B(n1630), .Y(n29412) );
  AND2X1 U29669 ( .A(n29413), .B(n29414), .Y(n29410) );
  NAND2X1 U29670 ( .A(n29415), .B(n29416), .Y(n29414) );
  NAND2X1 U29671 ( .A(u_muldiv_divisor_q[28]), .B(n805), .Y(n29416) );
  NOR2X1 U29672 ( .A(n29417), .B(n29418), .Y(n29415) );
  AND2X1 U29673 ( .A(n1561), .B(n29419), .Y(n29418) );
  NOR2X1 U29674 ( .A(n29420), .B(n37573), .Y(n29417) );
  NOR2X1 U29675 ( .A(n1561), .B(n29419), .Y(n29420) );
  NAND2X1 U29676 ( .A(n29421), .B(n29422), .Y(n29419) );
  NAND2X1 U29679 ( .A(n29424), .B(n1511), .Y(n29421) );
  NAND2X1 U29680 ( .A(n29425), .B(n29426), .Y(n29424) );
  NAND2X1 U29681 ( .A(u_muldiv_divisor_q[25]), .B(n29427), .Y(n29426) );
  NAND2X1 U29682 ( .A(u_muldiv_dividend_q[25]), .B(n29428), .Y(n29427) );
  OR2X1 U29683 ( .A(n29428), .B(u_muldiv_dividend_q[25]), .Y(n29425) );
  NAND2X1 U29684 ( .A(n29429), .B(n29430), .Y(n29428) );
  NAND2X1 U29685 ( .A(n29431), .B(n29432), .Y(n29430) );
  NAND2X1 U29686 ( .A(u_muldiv_divisor_q[24]), .B(n1582), .Y(n29432) );
  NOR2X1 U29687 ( .A(n29433), .B(n29434), .Y(n29431) );
  AND2X1 U29688 ( .A(n1459), .B(n29435), .Y(n29434) );
  NOR2X1 U29689 ( .A(n29436), .B(n37557), .Y(n29433) );
  NOR2X1 U29690 ( .A(n1459), .B(n29435), .Y(n29436) );
  NAND2X1 U29691 ( .A(n29437), .B(n29438), .Y(n29435) );
  NAND2X1 U29694 ( .A(n29440), .B(n1471), .Y(n29437) );
  NAND2X1 U29695 ( .A(n29441), .B(n29442), .Y(n29440) );
  NAND2X1 U29696 ( .A(u_muldiv_divisor_q[21]), .B(n29443), .Y(n29442) );
  NAND2X1 U29697 ( .A(u_muldiv_dividend_q[21]), .B(n29444), .Y(n29443) );
  OR2X1 U29698 ( .A(n29444), .B(u_muldiv_dividend_q[21]), .Y(n29441) );
  NAND2X1 U29699 ( .A(n29445), .B(n29446), .Y(n29444) );
  NAND2X1 U29700 ( .A(n29447), .B(n29448), .Y(n29446) );
  NAND2X1 U29701 ( .A(u_muldiv_divisor_q[20]), .B(n1439), .Y(n29448) );
  NOR2X1 U29702 ( .A(n29449), .B(n29450), .Y(n29447) );
  AND2X1 U29703 ( .A(n1409), .B(n29451), .Y(n29450) );
  NOR2X1 U29704 ( .A(n29452), .B(n37538), .Y(n29449) );
  NOR2X1 U29705 ( .A(n1409), .B(n29451), .Y(n29452) );
  NAND2X1 U29706 ( .A(n29453), .B(n29454), .Y(n29451) );
  NAND2X1 U29709 ( .A(n29456), .B(n37461), .Y(n29453) );
  NAND2X1 U29710 ( .A(n29457), .B(n29458), .Y(n29456) );
  NAND2X1 U29711 ( .A(u_muldiv_divisor_q[17]), .B(n29459), .Y(n29458) );
  NAND2X1 U29712 ( .A(u_muldiv_dividend_q[17]), .B(n29460), .Y(n29459) );
  OR2X1 U29713 ( .A(n29460), .B(u_muldiv_dividend_q[17]), .Y(n29457) );
  NAND2X1 U29714 ( .A(n29461), .B(n29462), .Y(n29460) );
  NAND2X1 U29715 ( .A(n29463), .B(n29464), .Y(n29462) );
  NAND2X1 U29716 ( .A(u_muldiv_divisor_q[16]), .B(n37451), .Y(n29464) );
  NOR2X1 U29717 ( .A(n29465), .B(n29466), .Y(n29463) );
  AND2X1 U29718 ( .A(n37446), .B(n29467), .Y(n29466) );
  NOR2X1 U29719 ( .A(n29468), .B(n37447), .Y(n29465) );
  NOR2X1 U29720 ( .A(n37446), .B(n29467), .Y(n29468) );
  NAND2X1 U29721 ( .A(n29469), .B(n29470), .Y(n29467) );
  NAND2X1 U29724 ( .A(n29472), .B(n37445), .Y(n29469) );
  NAND2X1 U29725 ( .A(n29473), .B(n29474), .Y(n29472) );
  NAND2X1 U29726 ( .A(u_muldiv_divisor_q[13]), .B(n29475), .Y(n29474) );
  NAND2X1 U29727 ( .A(u_muldiv_dividend_q[13]), .B(n29476), .Y(n29475) );
  OR2X1 U29728 ( .A(n29476), .B(u_muldiv_dividend_q[13]), .Y(n29473) );
  NAND2X1 U29729 ( .A(n29477), .B(n29478), .Y(n29476) );
  NAND2X1 U29730 ( .A(n29479), .B(n29480), .Y(n29478) );
  NAND2X1 U29731 ( .A(u_muldiv_divisor_q[12]), .B(n37441), .Y(n29480) );
  NOR2X1 U29732 ( .A(n29481), .B(n29482), .Y(n29479) );
  AND2X1 U29733 ( .A(n37439), .B(n29483), .Y(n29482) );
  NOR2X1 U29734 ( .A(n29484), .B(n37440), .Y(n29481) );
  NOR2X1 U29735 ( .A(n37439), .B(n29483), .Y(n29484) );
  NAND2X1 U29736 ( .A(n29485), .B(n29486), .Y(n29483) );
  NAND2X1 U29739 ( .A(n29488), .B(n37437), .Y(n29485) );
  NAND2X1 U29740 ( .A(n29489), .B(n29490), .Y(n29488) );
  NAND2X1 U29741 ( .A(u_muldiv_divisor_q[9]), .B(n29491), .Y(n29490) );
  NAND2X1 U29742 ( .A(u_muldiv_dividend_q[9]), .B(n29492), .Y(n29491) );
  OR2X1 U29743 ( .A(n29492), .B(u_muldiv_dividend_q[9]), .Y(n29489) );
  NAND2X1 U29744 ( .A(n29493), .B(n29494), .Y(n29492) );
  NAND2X1 U29745 ( .A(n29495), .B(n29496), .Y(n29494) );
  NAND2X1 U29746 ( .A(u_muldiv_divisor_q[8]), .B(n37428), .Y(n29496) );
  NOR2X1 U29747 ( .A(n29497), .B(n29498), .Y(n29495) );
  AND2X1 U29748 ( .A(n37426), .B(n29499), .Y(n29498) );
  NOR2X1 U29749 ( .A(n29500), .B(n37427), .Y(n29497) );
  NOR2X1 U29750 ( .A(n37426), .B(n29499), .Y(n29500) );
  NAND2X1 U29751 ( .A(n29501), .B(n29502), .Y(n29499) );
  NAND2X1 U29752 ( .A(u_muldiv_divisor_q[6]), .B(n29503), .Y(n29502) );
  OR2X1 U29753 ( .A(n29504), .B(n37423), .Y(n29503) );
  NAND2X1 U29754 ( .A(n29504), .B(n37423), .Y(n29501) );
  NAND2X1 U29755 ( .A(n29505), .B(n29506), .Y(n29504) );
  NAND2X1 U29756 ( .A(u_muldiv_divisor_q[5]), .B(n29507), .Y(n29506) );
  NAND2X1 U29757 ( .A(u_muldiv_dividend_q[5]), .B(n29508), .Y(n29507) );
  OR2X1 U29758 ( .A(n29508), .B(u_muldiv_dividend_q[5]), .Y(n29505) );
  NAND2X1 U29759 ( .A(n29509), .B(n29510), .Y(n29508) );
  NAND2X1 U29760 ( .A(n29511), .B(n29512), .Y(n29510) );
  NAND2X1 U29761 ( .A(u_muldiv_divisor_q[4]), .B(n37420), .Y(n29512) );
  NOR2X1 U29762 ( .A(n29513), .B(n29514), .Y(n29511) );
  NOR2X1 U29763 ( .A(u_muldiv_dividend_q[3]), .B(n37438), .Y(n29514) );
  NOR2X1 U29764 ( .A(n14835), .B(n29515), .Y(n29513) );
  NOR2X1 U29765 ( .A(n29516), .B(n29517), .Y(n29515) );
  NOR2X1 U29766 ( .A(u_muldiv_dividend_q[2]), .B(n37435), .Y(n29517) );
  NOR2X1 U29767 ( .A(n14854), .B(n14857), .Y(n29516) );
  NAND2X1 U29768 ( .A(n29518), .B(n29519), .Y(n14857) );
  NAND2X1 U29769 ( .A(n29520), .B(n37419), .Y(n29519) );
  OR2X1 U29770 ( .A(n14881), .B(u_muldiv_dividend_q[1]), .Y(n29520) );
  NAND2X1 U29771 ( .A(u_muldiv_dividend_q[1]), .B(n14881), .Y(n29518) );
  OR2X1 U29772 ( .A(n37418), .B(u_muldiv_dividend_q[0]), .Y(n14881) );
  NOR2X1 U29773 ( .A(n37325), .B(u_muldiv_divisor_q[2]), .Y(n14854) );
  NOR2X1 U29774 ( .A(n37326), .B(u_muldiv_divisor_q[3]), .Y(n14835) );
  NAND2X1 U29775 ( .A(u_muldiv_dividend_q[4]), .B(n37421), .Y(n29509) );
  NAND2X1 U29776 ( .A(u_muldiv_dividend_q[8]), .B(n37429), .Y(n29493) );
  NAND2X1 U29777 ( .A(u_muldiv_dividend_q[12]), .B(n37442), .Y(n29477) );
  NAND2X1 U29778 ( .A(u_muldiv_dividend_q[16]), .B(n37452), .Y(n29461) );
  NAND2X1 U29779 ( .A(u_muldiv_dividend_q[20]), .B(n37543), .Y(n29445) );
  NAND2X1 U29780 ( .A(u_muldiv_dividend_q[24]), .B(n37559), .Y(n29429) );
  NAND2X1 U29781 ( .A(u_muldiv_dividend_q[28]), .B(n37576), .Y(n29413) );
  NOR2X1 U29782 ( .A(n37582), .B(u_muldiv_dividend_q[30]), .Y(n14461) );
  NAND2X1 U29783 ( .A(u_muldiv_dividend_q[30]), .B(n37582), .Y(n14474) );
  NAND2X1 U29784 ( .A(n29521), .B(n29522), .Y(n29395) );
  NOR2X1 U29785 ( .A(n29523), .B(n29524), .Y(n29522) );
  OR2X1 U29786 ( .A(u_muldiv_divisor_q[41]), .B(u_muldiv_divisor_q[42]), .Y(
        n29524) );
  NAND2X1 U29787 ( .A(n29525), .B(n37590), .Y(n29523) );
  NOR2X1 U29788 ( .A(u_muldiv_divisor_q[45]), .B(u_muldiv_divisor_q[44]), .Y(
        n29525) );
  NOR2X1 U29789 ( .A(n29526), .B(n29527), .Y(n29521) );
  OR2X1 U29790 ( .A(u_muldiv_divisor_q[37]), .B(u_muldiv_divisor_q[38]), .Y(
        n29527) );
  OR2X1 U29791 ( .A(u_muldiv_divisor_q[39]), .B(u_muldiv_divisor_q[40]), .Y(
        n29526) );
  NAND2X1 U29792 ( .A(challenge[25]), .B(n44849), .Y(n29375) );
  NAND2X1 U29793 ( .A(n29528), .B(n29529), .Y(n17232) );
  NAND2X1 U29794 ( .A(challenge[24]), .B(n44849), .Y(n29528) );
  NAND2X1 U29795 ( .A(n29530), .B(n29529), .Y(n17231) );
  NAND2X1 U29796 ( .A(challenge[23]), .B(n44849), .Y(n29530) );
  NAND2X1 U29797 ( .A(n29531), .B(n29529), .Y(n17230) );
  NAND2X1 U29798 ( .A(challenge[22]), .B(n44849), .Y(n29531) );
  NAND2X1 U29799 ( .A(n29532), .B(n29529), .Y(n17229) );
  NAND2X1 U29800 ( .A(challenge[21]), .B(n44849), .Y(n29532) );
  NAND2X1 U29801 ( .A(n29533), .B(n29529), .Y(n17228) );
  NAND2X1 U29802 ( .A(u_muldiv_N264), .B(n44847), .Y(n29529) );
  NAND2X1 U29803 ( .A(n28813), .B(n44624), .Y(u_muldiv_N264) );
  NOR2X1 U29806 ( .A(n29536), .B(n29537), .Y(n29535) );
  NAND2X1 U29807 ( .A(n29538), .B(n29539), .Y(n29537) );
  NAND2X1 U29814 ( .A(n29544), .B(n29545), .Y(n29536) );
  NOR2X1 U29815 ( .A(n29546), .B(n29547), .Y(n29545) );
  OR2X1 U29816 ( .A(u_muldiv_q_mask_q[5]), .B(u_muldiv_q_mask_q[6]), .Y(n29547) );
  NOR2X1 U29819 ( .A(n29549), .B(n29550), .Y(n29544) );
  OR2X1 U29820 ( .A(u_muldiv_q_mask_q[30]), .B(u_muldiv_q_mask_q[31]), .Y(
        n29550) );
  OR2X1 U29821 ( .A(u_muldiv_q_mask_q[3]), .B(u_muldiv_q_mask_q[4]), .Y(n29549) );
  NOR2X1 U29822 ( .A(n29551), .B(n29552), .Y(n29534) );
  NAND2X1 U29823 ( .A(n29553), .B(n29554), .Y(n29552) );
  NOR2X1 U29824 ( .A(n29555), .B(n29556), .Y(n29554) );
  OR2X1 U29825 ( .A(u_muldiv_q_mask_q[12]), .B(u_muldiv_q_mask_q[13]), .Y(
        n29556) );
  OR2X1 U29826 ( .A(u_muldiv_q_mask_q[14]), .B(u_muldiv_q_mask_q[15]), .Y(
        n29555) );
  NOR2X1 U29827 ( .A(n29557), .B(n29558), .Y(n29553) );
  OR2X1 U29828 ( .A(n37436), .B(u_muldiv_q_mask_q[0]), .Y(n29558) );
  OR2X1 U29829 ( .A(u_muldiv_q_mask_q[10]), .B(u_muldiv_q_mask_q[11]), .Y(
        n29557) );
  NAND2X1 U29830 ( .A(n29559), .B(n29560), .Y(n29551) );
  NOR2X1 U29831 ( .A(n29561), .B(n29562), .Y(n29560) );
  OR2X1 U29832 ( .A(u_muldiv_q_mask_q[1]), .B(u_muldiv_q_mask_q[20]), .Y(
        n29562) );
  OR2X1 U29833 ( .A(u_muldiv_q_mask_q[21]), .B(u_muldiv_q_mask_q[22]), .Y(
        n29561) );
  NOR2X1 U29834 ( .A(n29563), .B(n29564), .Y(n29559) );
  OR2X1 U29835 ( .A(u_muldiv_q_mask_q[16]), .B(u_muldiv_q_mask_q[17]), .Y(
        n29564) );
  OR2X1 U29836 ( .A(u_muldiv_q_mask_q[18]), .B(u_muldiv_q_mask_q[19]), .Y(
        n29563) );
  NAND2X1 U29839 ( .A(challenge[20]), .B(n44849), .Y(n29533) );
  NAND2X1 U29840 ( .A(n29567), .B(n29568), .Y(n17227) );
  NAND2X1 U29841 ( .A(n42962), .B(n44857), .Y(n29568) );
  AND2X1 U29843 ( .A(n26327), .B(n73543), .Y(n29569) );
  NAND2X1 U29844 ( .A(n29570), .B(n73576), .Y(n26327) );
  NAND2X1 U29845 ( .A(n73418), .B(n28558), .Y(n27325) );
  NOR2X1 U29849 ( .A(n28034), .B(n29574), .Y(n29571) );
  NAND2X1 U29850 ( .A(n73532), .B(n29575), .Y(n29574) );
  NAND2X1 U29851 ( .A(n29576), .B(n28166), .Y(n29575) );
  NOR2X1 U29852 ( .A(n28174), .B(n28175), .Y(n28166) );
  NAND2X1 U29853 ( .A(n28194), .B(n28192), .Y(n28175) );
  NAND2X1 U29854 ( .A(n29577), .B(n29578), .Y(n28192) );
  NOR2X1 U29855 ( .A(n1086), .B(n29579), .Y(n29578) );
  AND2X1 U29856 ( .A(n73519), .B(u_csr_csr_mideleg_q[5]), .Y(n29579) );
  NOR2X1 U29857 ( .A(n37331), .B(n37546), .Y(n29577) );
  NAND2X1 U29858 ( .A(n29580), .B(n29581), .Y(n28194) );
  NOR2X1 U29859 ( .A(n1086), .B(n29582), .Y(n29581) );
  AND2X1 U29860 ( .A(n73519), .B(u_csr_csr_mideleg_q[7]), .Y(n29582) );
  NOR2X1 U29861 ( .A(n37330), .B(n37545), .Y(n29580) );
  NAND2X1 U29862 ( .A(n28189), .B(n28195), .Y(n28174) );
  NAND2X1 U29863 ( .A(n29583), .B(n29584), .Y(n28195) );
  NOR2X1 U29864 ( .A(n1086), .B(n29585), .Y(n29584) );
  AND2X1 U29865 ( .A(n73519), .B(u_csr_csr_mideleg_q[1]), .Y(n29585) );
  AND2X1 U29866 ( .A(u_csr_csr_mie_q_1), .B(u_csr_csr_mip_q_1), .Y(n29583) );
  NAND2X1 U29867 ( .A(n29586), .B(n29587), .Y(n28189) );
  NOR2X1 U29868 ( .A(n1086), .B(n29588), .Y(n29587) );
  NOR2X1 U29869 ( .A(n28520), .B(n37533), .Y(n29588) );
  NOR2X1 U29870 ( .A(n37544), .B(n37335), .Y(n29586) );
  NOR2X1 U29871 ( .A(n28193), .B(n29589), .Y(n29576) );
  NOR2X1 U29872 ( .A(n37553), .B(n29590), .Y(n29589) );
  NAND2X1 U29873 ( .A(\u_csr_csr_mie_q[11] ), .B(n29591), .Y(n29590) );
  AND2X1 U29874 ( .A(n29592), .B(n29593), .Y(n28193) );
  NOR2X1 U29875 ( .A(n1086), .B(n29594), .Y(n29593) );
  NOR2X1 U29876 ( .A(n28520), .B(n37531), .Y(n29594) );
  NAND2X1 U29877 ( .A(n28520), .B(n29595), .Y(n29591) );
  NAND2X1 U29878 ( .A(n73568), .B(n29596), .Y(n29595) );
  NAND2X1 U29879 ( .A(n37540), .B(u_csr_N3161), .Y(n29596) );
  NAND2X1 U29881 ( .A(n29599), .B(u_csr_N3162), .Y(n29598) );
  NOR2X1 U29882 ( .A(u_csr_csr_sr_q[3]), .B(n73569), .Y(n29599) );
  NAND2X1 U29883 ( .A(n29600), .B(n29601), .Y(n29597) );
  NOR2X1 U29884 ( .A(n29602), .B(n29603), .Y(n29601) );
  NAND2X1 U29885 ( .A(n29604), .B(n29605), .Y(n29603) );
  NAND2X1 U29886 ( .A(n29606), .B(\u_csr_csr_mip_q[11] ), .Y(n29605) );
  NOR2X1 U29887 ( .A(u_csr_csr_mideleg_q[11]), .B(n37485), .Y(n29606) );
  NAND2X1 U29888 ( .A(n29607), .B(u_csr_csr_mip_q_1), .Y(n29604) );
  NOR2X1 U29890 ( .A(n37335), .B(n29608), .Y(n29602) );
  NAND2X1 U29891 ( .A(u_csr_csr_mie_q_3), .B(n37533), .Y(n29608) );
  NOR2X1 U29892 ( .A(n29609), .B(n29610), .Y(n29600) );
  NAND2X1 U29893 ( .A(n29611), .B(n29612), .Y(n29610) );
  NAND2X1 U29894 ( .A(n29613), .B(u_csr_csr_mip_q_5), .Y(n29612) );
  NOR2X1 U29895 ( .A(u_csr_csr_mideleg_q[5]), .B(n37331), .Y(n29613) );
  NAND2X1 U29896 ( .A(n29614), .B(u_csr_csr_mip_q_7), .Y(n29611) );
  NOR2X1 U29897 ( .A(u_csr_csr_mideleg_q[7]), .B(n37330), .Y(n29614) );
  NOR2X1 U29898 ( .A(n37334), .B(n29615), .Y(n29609) );
  NAND2X1 U29899 ( .A(u_csr_csr_mie_q_9), .B(n37531), .Y(n29615) );
  NOR2X1 U29900 ( .A(n37549), .B(n37334), .Y(n29592) );
  NAND2X1 U29908 ( .A(n28204), .B(n26138), .Y(n29620) );
  NAND2X1 U29910 ( .A(n29621), .B(n29622), .Y(n28204) );
  NOR2X1 U29911 ( .A(mem_d_resp_tag_i[9]), .B(n487), .Y(n29622) );
  NOR2X1 U29912 ( .A(n29623), .B(n575), .Y(n29621) );
  NAND2X1 U29918 ( .A(n73543), .B(n29628), .Y(n29627) );
  NAND2X1 U29919 ( .A(n29629), .B(n29630), .Y(n29628) );
  NOR2X1 U29921 ( .A(n29631), .B(n29632), .Y(n29629) );
  NOR2X1 U29922 ( .A(n29633), .B(n25635), .Y(n29632) );
  NAND2X1 U29932 ( .A(n26129), .B(n44083), .Y(n29640) );
  NOR2X1 U29936 ( .A(n29634), .B(n24367), .Y(n26129) );
  NAND2X1 U29940 ( .A(challenge[19]), .B(n44849), .Y(n29567) );
  NAND2X1 U29941 ( .A(n29643), .B(n29644), .Y(n17226) );
  NAND2X1 U29942 ( .A(challenge[18]), .B(n44849), .Y(n29643) );
  NAND2X1 U29943 ( .A(n29645), .B(n29644), .Y(n17225) );
  NAND2X1 U29944 ( .A(challenge[17]), .B(n44849), .Y(n29645) );
  NAND2X1 U29945 ( .A(n29646), .B(n29644), .Y(n17224) );
  NAND2X1 U29946 ( .A(challenge[16]), .B(n44849), .Y(n29646) );
  NAND2X1 U29947 ( .A(n29647), .B(n29644), .Y(n17223) );
  NAND2X1 U29951 ( .A(challenge[15]), .B(n44849), .Y(n29647) );
  NAND2X1 U29952 ( .A(n29649), .B(n29650), .Y(n17222) );
  NAND2X1 U29953 ( .A(challenge[14]), .B(n44849), .Y(n29649) );
  NAND2X1 U29954 ( .A(n29651), .B(n29650), .Y(n17221) );
  NAND2X1 U29955 ( .A(challenge[13]), .B(n44848), .Y(n29651) );
  NAND2X1 U29956 ( .A(n29652), .B(n29650), .Y(n17220) );
  NAND2X1 U29957 ( .A(challenge[12]), .B(n44848), .Y(n29652) );
  NAND2X1 U29958 ( .A(n29653), .B(n29650), .Y(n17219) );
  NAND2X1 U29959 ( .A(challenge[11]), .B(n44848), .Y(n29653) );
  NAND2X1 U29960 ( .A(n29654), .B(n29650), .Y(n17218) );
  NAND2X1 U29961 ( .A(n28934), .B(n44861), .Y(n29650) );
  NAND2X1 U29962 ( .A(challenge[10]), .B(n44848), .Y(n29654) );
  NAND2X1 U29964 ( .A(challenge[9]), .B(n44848), .Y(n29655) );
  NAND2X1 U29967 ( .A(challenge[8]), .B(n44848), .Y(n29657) );
  NAND2X1 U29977 ( .A(n29664), .B(n29665), .Y(n17212) );
  NAND2X1 U29978 ( .A(n28797), .B(n44857), .Y(n29665) );
  NAND2X1 U29983 ( .A(challenge[4]), .B(n44848), .Y(n29664) );
  NAND2X1 U29984 ( .A(n29669), .B(n29670), .Y(n17211) );
  NAND2X1 U29985 ( .A(challenge[3]), .B(n44848), .Y(n29669) );
  NAND2X1 U29986 ( .A(n29671), .B(n29670), .Y(n17210) );
  NAND2X1 U29987 ( .A(n37548), .B(n44857), .Y(n29670) );
  NAND2X1 U29990 ( .A(challenge[2]), .B(n44848), .Y(n29671) );
  NAND2X1 U29991 ( .A(n29673), .B(n29674), .Y(n17209) );
  NAND2X1 U29992 ( .A(challenge[1]), .B(n44848), .Y(n29673) );
  NAND2X1 U29993 ( .A(n29675), .B(n29674), .Y(n17208) );
  NAND2X1 U29994 ( .A(n73429), .B(n44858), .Y(n29674) );
  NAND2X1 U29997 ( .A(challenge[0]), .B(n44846), .Y(n29675) );
  NOR2X1 U29998 ( .A(n29677), .B(n29013), .Y(mem_i_rd_o) );
  NOR2X1 U30002 ( .A(n29681), .B(n29682), .Y(n29680) );
  NOR2X1 U30003 ( .A(u_mmu_itlb_entry_q_4), .B(u_csr_N3161), .Y(n29682) );
  XNOR2X1 U30011 ( .A(n29691), .B(n29692), .Y(n29690) );
  XOR2X1 U30017 ( .A(n29692), .B(n29702), .Y(n29701) );
  NAND2X1 U30018 ( .A(n29703), .B(n29704), .Y(n29692) );
  XNOR2X1 U30028 ( .A(n29713), .B(n29714), .Y(n29712) );
  XOR2X1 U30034 ( .A(n29714), .B(n29723), .Y(n29722) );
  NAND2X1 U30035 ( .A(n29724), .B(n29725), .Y(n29714) );
  XNOR2X1 U30045 ( .A(n29734), .B(n29735), .Y(n29733) );
  XOR2X1 U30051 ( .A(n29735), .B(n29744), .Y(n29743) );
  NAND2X1 U30052 ( .A(n29745), .B(n29746), .Y(n29735) );
  XNOR2X1 U30062 ( .A(n29755), .B(n29756), .Y(n29754) );
  XOR2X1 U30068 ( .A(n29756), .B(n29765), .Y(n29764) );
  NAND2X1 U30069 ( .A(n29766), .B(n29767), .Y(n29756) );
  NAND2X1 U30086 ( .A(n29787), .B(n29788), .Y(n29777) );
  XNOR2X1 U30244 ( .A(n29930), .B(n29931), .Y(n29929) );
  XOR2X1 U30250 ( .A(n29931), .B(n29940), .Y(n29939) );
  NAND2X1 U30251 ( .A(n29941), .B(n29942), .Y(n29931) );
  NAND2X1 U30281 ( .A(n1885), .B(n44263), .Y(mem_d_req_tag_o[9]) );
  NAND2X1 U30282 ( .A(n1884), .B(n44261), .Y(mem_d_req_tag_o[8]) );
  NAND2X1 U30283 ( .A(n36758), .B(n8255), .Y(mem_d_req_tag_o[7]) );
  NOR2X1 U30284 ( .A(n1883), .B(n44258), .Y(mem_d_req_tag_o[6]) );
  NOR2X1 U30285 ( .A(n1882), .B(n44258), .Y(mem_d_req_tag_o[5]) );
  NOR2X1 U30288 ( .A(n1879), .B(n44258), .Y(mem_d_req_tag_o[2]) );
  NOR2X1 U30289 ( .A(n1878), .B(n44258), .Y(mem_d_req_tag_o[1]) );
  NOR2X1 U30290 ( .A(n1886), .B(n44258), .Y(mem_d_req_tag_o[10]) );
  NOR2X1 U30292 ( .A(n8647), .B(n44258), .Y(mem_d_invalidate_o) );
  NOR2X1 U30293 ( .A(n8954), .B(n44258), .Y(mem_d_flush_o) );
  NOR2X1 U30294 ( .A(n2752), .B(n44258), .Y(mem_d_data_wr_o[9]) );
  NOR2X1 U30295 ( .A(n2950), .B(n44258), .Y(mem_d_data_wr_o[8]) );
  NOR2X1 U30296 ( .A(n2613), .B(n44258), .Y(mem_d_data_wr_o[7]) );
  NOR2X1 U30297 ( .A(n2348), .B(n44258), .Y(mem_d_data_wr_o[6]) );
  NOR2X1 U30298 ( .A(n2946), .B(n44259), .Y(mem_d_data_wr_o[5]) );
  NOR2X1 U30299 ( .A(n2748), .B(n44259), .Y(mem_d_data_wr_o[4]) );
  NOR2X1 U30300 ( .A(n2416), .B(n44259), .Y(mem_d_data_wr_o[3]) );
  NOR2X1 U30301 ( .A(n2616), .B(n44259), .Y(mem_d_data_wr_o[31]) );
  NOR2X1 U30302 ( .A(n3043), .B(n44259), .Y(mem_d_data_wr_o[30]) );
  NOR2X1 U30303 ( .A(n2349), .B(n44259), .Y(mem_d_data_wr_o[2]) );
  NOR2X1 U30304 ( .A(n3012), .B(n44259), .Y(mem_d_data_wr_o[29]) );
  NOR2X1 U30305 ( .A(n2953), .B(n44259), .Y(mem_d_data_wr_o[28]) );
  NOR2X1 U30306 ( .A(n2816), .B(n44259), .Y(mem_d_data_wr_o[27]) );
  NOR2X1 U30307 ( .A(n2649), .B(n44259), .Y(mem_d_data_wr_o[26]) );
  NOR2X1 U30308 ( .A(n2849), .B(n44259), .Y(mem_d_data_wr_o[25]) );
  NOR2X1 U30309 ( .A(n2952), .B(n44259), .Y(mem_d_data_wr_o[24]) );
  NOR2X1 U30310 ( .A(n2615), .B(n44259), .Y(mem_d_data_wr_o[23]) );
  NOR2X1 U30311 ( .A(n2515), .B(n44259), .Y(mem_d_data_wr_o[22]) );
  NOR2X1 U30312 ( .A(n2948), .B(n44260), .Y(mem_d_data_wr_o[21]) );
  NOR2X1 U30313 ( .A(n2750), .B(n44260), .Y(mem_d_data_wr_o[20]) );
  NOR2X1 U30314 ( .A(n2751), .B(n44260), .Y(mem_d_data_wr_o[1]) );
  NOR2X1 U30315 ( .A(n2418), .B(n44260), .Y(mem_d_data_wr_o[19]) );
  NOR2X1 U30316 ( .A(n2682), .B(n44260), .Y(mem_d_data_wr_o[18]) );
  NOR2X1 U30317 ( .A(n2915), .B(n44260), .Y(mem_d_data_wr_o[17]) );
  NOR2X1 U30318 ( .A(n2951), .B(n44260), .Y(mem_d_data_wr_o[16]) );
  NOR2X1 U30319 ( .A(n2614), .B(n44260), .Y(mem_d_data_wr_o[15]) );
  NOR2X1 U30320 ( .A(n3042), .B(n44260), .Y(mem_d_data_wr_o[14]) );
  NOR2X1 U30321 ( .A(n2947), .B(n44260), .Y(mem_d_data_wr_o[13]) );
  NOR2X1 U30322 ( .A(n2749), .B(n44260), .Y(mem_d_data_wr_o[12]) );
  NOR2X1 U30323 ( .A(n2417), .B(n44260), .Y(mem_d_data_wr_o[11]) );
  NOR2X1 U30324 ( .A(n2382), .B(n44260), .Y(mem_d_data_wr_o[10]) );
  NOR2X1 U30325 ( .A(n2949), .B(n44260), .Y(mem_d_data_wr_o[0]) );
  NOR2X1 U30326 ( .A(n29963), .B(n29964), .Y(mem_d_cacheable_o) );
  NAND2X1 U30327 ( .A(mem_d_addr_o[31]), .B(n697), .Y(n29964) );
  OR2X1 U30328 ( .A(mem_d_addr_o[29]), .B(mem_d_addr_o[30]), .Y(n29963) );
  NAND2X1 U30329 ( .A(n29965), .B(n29966), .Y(mem_d_addr_o[9]) );
  NOR2X1 U30331 ( .A(n29967), .B(n29968), .Y(n29965) );
  NAND2X1 U30334 ( .A(n29971), .B(n29972), .Y(mem_d_addr_o[8]) );
  NOR2X1 U30336 ( .A(n29973), .B(n29974), .Y(n29971) );
  NAND2X1 U30339 ( .A(n29975), .B(n29976), .Y(mem_d_addr_o[7]) );
  NOR2X1 U30341 ( .A(n29977), .B(n29978), .Y(n29975) );
  NAND2X1 U30344 ( .A(n29979), .B(n29980), .Y(mem_d_addr_o[6]) );
  NOR2X1 U30346 ( .A(n29981), .B(n29982), .Y(n29979) );
  NAND2X1 U30349 ( .A(n29983), .B(n29984), .Y(mem_d_addr_o[5]) );
  NOR2X1 U30351 ( .A(n29985), .B(n29986), .Y(n29983) );
  NAND2X1 U30354 ( .A(n29987), .B(n29988), .Y(mem_d_addr_o[4]) );
  NOR2X1 U30356 ( .A(n29989), .B(n29990), .Y(n29987) );
  NAND2X1 U30359 ( .A(n29991), .B(n29992), .Y(mem_d_addr_o[3]) );
  NOR2X1 U30361 ( .A(n29993), .B(n29994), .Y(n29991) );
  NAND2X1 U30364 ( .A(n29995), .B(n29996), .Y(mem_d_addr_o[31]) );
  NOR2X1 U30365 ( .A(n29997), .B(n29998), .Y(n29996) );
  NOR2X1 U30367 ( .A(n42974), .B(n1844), .Y(n29997) );
  NAND2X1 U30371 ( .A(n30003), .B(n30004), .Y(mem_d_addr_o[30]) );
  NOR2X1 U30374 ( .A(n42975), .B(n1843), .Y(n30005) );
  NOR2X1 U30375 ( .A(n30007), .B(n30008), .Y(n30003) );
  NAND2X1 U30378 ( .A(n30009), .B(n30010), .Y(mem_d_addr_o[2]) );
  NOR2X1 U30380 ( .A(n30011), .B(n30012), .Y(n30009) );
  NAND2X1 U30383 ( .A(n30013), .B(n30014), .Y(mem_d_addr_o[29]) );
  NOR2X1 U30384 ( .A(n30015), .B(n30016), .Y(n30014) );
  NOR2X1 U30386 ( .A(n42974), .B(n1842), .Y(n30015) );
  NOR2X1 U30387 ( .A(n30017), .B(n30018), .Y(n30013) );
  NAND2X1 U30390 ( .A(n30019), .B(n30020), .Y(mem_d_addr_o[28]) );
  NOR2X1 U30393 ( .A(n42976), .B(n1841), .Y(n30021) );
  NOR2X1 U30394 ( .A(n30023), .B(n30024), .Y(n30019) );
  NAND2X1 U30397 ( .A(n30025), .B(n30026), .Y(mem_d_addr_o[27]) );
  NOR2X1 U30398 ( .A(n30027), .B(n30028), .Y(n30026) );
  NOR2X1 U30400 ( .A(n42976), .B(n1840), .Y(n30027) );
  NAND2X1 U30404 ( .A(n30031), .B(n30032), .Y(mem_d_addr_o[26]) );
  NOR2X1 U30405 ( .A(n30033), .B(n30034), .Y(n30032) );
  NOR2X1 U30407 ( .A(n42974), .B(n1839), .Y(n30033) );
  NAND2X1 U30411 ( .A(n30037), .B(n30038), .Y(mem_d_addr_o[25]) );
  NOR2X1 U30412 ( .A(n30039), .B(n30040), .Y(n30038) );
  NOR2X1 U30414 ( .A(n42976), .B(n1838), .Y(n30039) );
  NOR2X1 U30415 ( .A(n30041), .B(n30042), .Y(n30037) );
  NAND2X1 U30418 ( .A(n30043), .B(n30044), .Y(mem_d_addr_o[24]) );
  NOR2X1 U30421 ( .A(n42975), .B(n1847), .Y(n30045) );
  NOR2X1 U30422 ( .A(n30047), .B(n30048), .Y(n30043) );
  NAND2X1 U30425 ( .A(n30049), .B(n30050), .Y(mem_d_addr_o[23]) );
  NOR2X1 U30428 ( .A(n42975), .B(n1846), .Y(n30051) );
  NOR2X1 U30429 ( .A(n30053), .B(n30054), .Y(n30049) );
  NAND2X1 U30432 ( .A(n30055), .B(n30056), .Y(mem_d_addr_o[22]) );
  NOR2X1 U30435 ( .A(n42976), .B(n1845), .Y(n30057) );
  NAND2X1 U30439 ( .A(n30061), .B(n30062), .Y(mem_d_addr_o[21]) );
  NOR2X1 U30440 ( .A(n30063), .B(n30064), .Y(n30062) );
  NOR2X1 U30442 ( .A(n42976), .B(n2550), .Y(n30063) );
  NAND2X1 U30446 ( .A(n30067), .B(n30068), .Y(mem_d_addr_o[20]) );
  NOR2X1 U30447 ( .A(n30069), .B(n30070), .Y(n30068) );
  NOR2X1 U30449 ( .A(n42974), .B(n2385), .Y(n30069) );
  NOR2X1 U30450 ( .A(n30071), .B(n30072), .Y(n30067) );
  NAND2X1 U30453 ( .A(n30073), .B(n30074), .Y(mem_d_addr_o[1]) );
  NAND2X1 U30456 ( .A(n30075), .B(n30076), .Y(mem_d_addr_o[19]) );
  NOR2X1 U30457 ( .A(n30077), .B(n30078), .Y(n30076) );
  NOR2X1 U30459 ( .A(n42975), .B(n2285), .Y(n30077) );
  NOR2X1 U30460 ( .A(n30079), .B(n30080), .Y(n30075) );
  NAND2X1 U30463 ( .A(n30081), .B(n30082), .Y(mem_d_addr_o[18]) );
  NOR2X1 U30467 ( .A(n30085), .B(n30086), .Y(n30081) );
  NAND2X1 U30470 ( .A(n30087), .B(n30088), .Y(mem_d_addr_o[17]) );
  NAND2X1 U30477 ( .A(n30093), .B(n30094), .Y(mem_d_addr_o[16]) );
  NOR2X1 U30478 ( .A(n30095), .B(n30096), .Y(n30094) );
  NOR2X1 U30480 ( .A(n42974), .B(n2518), .Y(n30095) );
  NOR2X1 U30481 ( .A(n30097), .B(n30098), .Y(n30093) );
  NAND2X1 U30484 ( .A(n30099), .B(n30100), .Y(mem_d_addr_o[15]) );
  NAND2X1 U30491 ( .A(n30105), .B(n30106), .Y(mem_d_addr_o[14]) );
  NOR2X1 U30495 ( .A(n30109), .B(n30110), .Y(n30105) );
  NAND2X1 U30498 ( .A(n30111), .B(n30112), .Y(mem_d_addr_o[13]) );
  NOR2X1 U30499 ( .A(n30113), .B(n30114), .Y(n30112) );
  NOR2X1 U30501 ( .A(n42974), .B(n2754), .Y(n30113) );
  NAND2X1 U30505 ( .A(n30117), .B(n30118), .Y(mem_d_addr_o[12]) );
  NAND2X1 U30516 ( .A(n30123), .B(n30124), .Y(mem_d_addr_o[11]) );
  NOR2X1 U30518 ( .A(n30125), .B(n30126), .Y(n30123) );
  NAND2X1 U30521 ( .A(n30127), .B(n30128), .Y(mem_d_addr_o[10]) );
  NOR2X1 U30523 ( .A(n30129), .B(n30130), .Y(n30127) );
  NAND2X1 U30526 ( .A(n30131), .B(n30132), .Y(mem_d_addr_o[0]) );
  NAND2X1 U30719 ( .A(n30271), .B(n30272), .Y(n28765) );
  NOR2X1 U30720 ( .A(n576), .B(n487), .Y(n30271) );
  AND2X1 U30722 ( .A(n30274), .B(n438), .Y(n28796) );
  NOR2X1 U30723 ( .A(mem_d_data_rd_i[3]), .B(mem_d_data_rd_i[2]), .Y(n30274)
         );
  NOR2X1 U30724 ( .A(mem_d_error_i), .B(n73554), .Y(n30273) );
  XNOR2X1 U30768 ( .A(n30318), .B(n30319), .Y(n30317) );
  XOR2X1 U30774 ( .A(n30319), .B(n30328), .Y(n30327) );
  NAND2X1 U30775 ( .A(n30329), .B(n30330), .Y(n30319) );
  NOR2X1 U30867 ( .A(n42437), .B(n30429), .Y(n30426) );
  NOR2X1 U30873 ( .A(n30429), .B(n30436), .Y(n30435) );
  XNOR2X1 U30905 ( .A(n30470), .B(n30471), .Y(n30469) );
  XOR2X1 U30911 ( .A(n30471), .B(n30480), .Y(n30479) );
  NAND2X1 U30912 ( .A(n30481), .B(n30482), .Y(n30471) );
  NAND2X1 U30925 ( .A(n30494), .B(n30495), .Y(n30493) );
  NAND2X1 U30933 ( .A(n30505), .B(n30494), .Y(n30504) );
  XNOR2X1 U30947 ( .A(n30514), .B(n30515), .Y(n30513) );
  XOR2X1 U30953 ( .A(n30515), .B(n30524), .Y(n30523) );
  NAND2X1 U30954 ( .A(n30525), .B(n30526), .Y(n30515) );
  NAND2X1 U30971 ( .A(n30456), .B(n30445), .Y(n30544) );
  NAND2X1 U30973 ( .A(n30414), .B(n30403), .Y(n30545) );
  NAND2X1 U30975 ( .A(n30548), .B(n30549), .Y(n30547) );
  NAND2X1 U30983 ( .A(n30455), .B(n30456), .Y(n30558) );
  NAND2X1 U30986 ( .A(n30413), .B(n30414), .Y(n30559) );
  NAND2X1 U30989 ( .A(n30561), .B(n30548), .Y(n30560) );
  XNOR2X1 U31005 ( .A(n30549), .B(n30570), .Y(n30569) );
  NAND2X1 U31006 ( .A(n30330), .B(n30571), .Y(n30549) );
  NAND2X1 U31007 ( .A(n30329), .B(n30318), .Y(n30571) );
  NAND2X1 U31008 ( .A(n30572), .B(n30573), .Y(n30318) );
  NAND2X1 U31009 ( .A(n30574), .B(n30575), .Y(n30573) );
  XOR2X1 U31015 ( .A(n30570), .B(n30561), .Y(n30583) );
  NAND2X1 U31016 ( .A(n30330), .B(n30584), .Y(n30561) );
  NAND2X1 U31017 ( .A(n30328), .B(n30329), .Y(n30584) );
  NAND2X1 U31019 ( .A(n30572), .B(n30585), .Y(n30328) );
  NAND2X1 U31020 ( .A(n30586), .B(n30574), .Y(n30585) );
  NAND2X1 U31022 ( .A(n30548), .B(n30546), .Y(n30570) );
  XNOR2X1 U31035 ( .A(n30595), .B(n30596), .Y(n30594) );
  XOR2X1 U31041 ( .A(n30596), .B(n30605), .Y(n30604) );
  NAND2X1 U31042 ( .A(n30606), .B(n30607), .Y(n30596) );
  XNOR2X1 U31054 ( .A(n30575), .B(n30617), .Y(n30616) );
  NAND2X1 U31055 ( .A(n30526), .B(n30618), .Y(n30575) );
  NAND2X1 U31056 ( .A(n30525), .B(n30514), .Y(n30618) );
  NAND2X1 U31057 ( .A(n30482), .B(n30619), .Y(n30514) );
  NAND2X1 U31058 ( .A(n30481), .B(n30470), .Y(n30619) );
  NAND2X1 U31059 ( .A(n30607), .B(n30620), .Y(n30470) );
  NAND2X1 U31060 ( .A(n30606), .B(n30595), .Y(n30620) );
  NAND2X1 U31061 ( .A(n30621), .B(n30622), .Y(n30595) );
  NAND2X1 U31062 ( .A(n30623), .B(n30624), .Y(n30622) );
  XOR2X1 U31068 ( .A(n30617), .B(n30586), .Y(n30632) );
  NAND2X1 U31069 ( .A(n30526), .B(n30633), .Y(n30586) );
  NAND2X1 U31070 ( .A(n30524), .B(n30525), .Y(n30633) );
  NAND2X1 U31072 ( .A(n30482), .B(n30634), .Y(n30524) );
  NAND2X1 U31073 ( .A(n30480), .B(n30481), .Y(n30634) );
  NAND2X1 U31075 ( .A(n30607), .B(n30635), .Y(n30480) );
  NAND2X1 U31076 ( .A(n30605), .B(n30606), .Y(n30635) );
  NAND2X1 U31078 ( .A(n30621), .B(n30636), .Y(n30605) );
  NAND2X1 U31079 ( .A(n30637), .B(n30623), .Y(n30636) );
  NAND2X1 U31083 ( .A(n30574), .B(n30572), .Y(n30617) );
  XNOR2X1 U31157 ( .A(n30624), .B(n30709), .Y(n30708) );
  NAND2X1 U31158 ( .A(n30710), .B(n30711), .Y(n30624) );
  NAND2X1 U31188 ( .A(n30623), .B(n30621), .Y(n30709) );
  NAND2X1 U31228 ( .A(n29941), .B(n29930), .Y(n30771) );
  NAND2X1 U31229 ( .A(n29704), .B(n30772), .Y(n29930) );
  NAND2X1 U31230 ( .A(n29703), .B(n29691), .Y(n30772) );
  NAND2X1 U31231 ( .A(n29725), .B(n30773), .Y(n29691) );
  NAND2X1 U31232 ( .A(n29724), .B(n29713), .Y(n30773) );
  NAND2X1 U31233 ( .A(n29746), .B(n30774), .Y(n29713) );
  NAND2X1 U31234 ( .A(n29745), .B(n29734), .Y(n30774) );
  NAND2X1 U31235 ( .A(n29767), .B(n30775), .Y(n29734) );
  NAND2X1 U31236 ( .A(n29766), .B(n29755), .Y(n30775) );
  NAND2X1 U31237 ( .A(n29788), .B(n30776), .Y(n29755) );
  NAND2X1 U31238 ( .A(n29787), .B(n29776), .Y(n30776) );
  NAND2X1 U31284 ( .A(n29940), .B(n29941), .Y(n30820) );
  NAND2X1 U31286 ( .A(n29704), .B(n30821), .Y(n29940) );
  NAND2X1 U31287 ( .A(n29702), .B(n29703), .Y(n30821) );
  NAND2X1 U31289 ( .A(n29725), .B(n30822), .Y(n29702) );
  NAND2X1 U31290 ( .A(n29723), .B(n29724), .Y(n30822) );
  NAND2X1 U31292 ( .A(n29746), .B(n30823), .Y(n29723) );
  NAND2X1 U31293 ( .A(n29744), .B(n29745), .Y(n30823) );
  NAND2X1 U31295 ( .A(n29767), .B(n30824), .Y(n29744) );
  NAND2X1 U31296 ( .A(n29765), .B(n29766), .Y(n30824) );
  NAND2X1 U31298 ( .A(n29788), .B(n30825), .Y(n29765) );
  NAND2X1 U31299 ( .A(n29786), .B(n29787), .Y(n30825) );
  NOR2X1 U31666 ( .A(n31128), .B(n31129), .Y(n31124) );
  NOR2X1 U31670 ( .A(n31132), .B(n31133), .Y(n31128) );
  NAND2X1 U31671 ( .A(n31134), .B(n31135), .Y(n31133) );
  NAND2X1 U31672 ( .A(n31136), .B(n31137), .Y(n31135) );
  NAND2X1 U31673 ( .A(n31138), .B(n31139), .Y(n31137) );
  NOR2X1 U31680 ( .A(n31144), .B(n31145), .Y(n31136) );
  NOR2X1 U31681 ( .A(n31146), .B(n31147), .Y(n31145) );
  NOR2X1 U31682 ( .A(n31148), .B(n31149), .Y(n31147) );
  NAND2X1 U31683 ( .A(n31150), .B(n31151), .Y(n31149) );
  NAND2X1 U31685 ( .A(n31153), .B(n31154), .Y(n31150) );
  NAND2X1 U31686 ( .A(n31155), .B(n31156), .Y(n31154) );
  NOR2X1 U31688 ( .A(n31158), .B(n31159), .Y(n31155) );
  NOR2X1 U31689 ( .A(n31160), .B(n31161), .Y(n31159) );
  NOR2X1 U31690 ( .A(n31162), .B(n31163), .Y(n31161) );
  NAND2X1 U31691 ( .A(n31164), .B(n31165), .Y(n31163) );
  NOR2X1 U31707 ( .A(n31176), .B(n31177), .Y(n31160) );
  NAND2X1 U31708 ( .A(n31178), .B(n31179), .Y(n31177) );
  NOR2X1 U31714 ( .A(n31182), .B(n31183), .Y(n31176) );
  NOR2X1 U31715 ( .A(n31184), .B(n31185), .Y(n31183) );
  NAND2X1 U31716 ( .A(n31186), .B(n31187), .Y(n31185) );
  NOR2X1 U31732 ( .A(n31198), .B(n31199), .Y(n31182) );
  NAND2X1 U31733 ( .A(n31200), .B(n31201), .Y(n31199) );
  NOR2X1 U31740 ( .A(n31204), .B(n31205), .Y(n31198) );
  NOR2X1 U31741 ( .A(n31206), .B(n31207), .Y(n31205) );
  NAND2X1 U31742 ( .A(n31208), .B(n31209), .Y(n31207) );
  NOR2X1 U31758 ( .A(n31220), .B(n31221), .Y(n31204) );
  NAND2X1 U31759 ( .A(n31222), .B(n31223), .Y(n31221) );
  NOR2X1 U31766 ( .A(n31226), .B(n31227), .Y(n31220) );
  NOR2X1 U31767 ( .A(n31228), .B(n31229), .Y(n31227) );
  NAND2X1 U31768 ( .A(n31230), .B(n31231), .Y(n31229) );
  NOR2X1 U31784 ( .A(n31242), .B(n31243), .Y(n31226) );
  NAND2X1 U31785 ( .A(n31244), .B(n31245), .Y(n31243) );
  NOR2X1 U31791 ( .A(n31248), .B(n31249), .Y(n31242) );
  NOR2X1 U31792 ( .A(n31250), .B(n31251), .Y(n31249) );
  NAND2X1 U31793 ( .A(n31252), .B(n31253), .Y(n31251) );
  NOR2X1 U31809 ( .A(n31264), .B(n31265), .Y(n31248) );
  NAND2X1 U31810 ( .A(n31266), .B(n31267), .Y(n31265) );
  NAND2X1 U31811 ( .A(n31268), .B(n31269), .Y(n31267) );
  NAND2X1 U31812 ( .A(n31270), .B(n31271), .Y(n31269) );
  NAND2X1 U31813 ( .A(n31272), .B(n31273), .Y(n31271) );
  NAND2X1 U31814 ( .A(n31274), .B(n31275), .Y(n31273) );
  NAND2X1 U31815 ( .A(n31276), .B(n31277), .Y(n31275) );
  NAND2X1 U31816 ( .A(n31278), .B(n31279), .Y(n31277) );
  NAND2X1 U31817 ( .A(n31280), .B(n31281), .Y(n31279) );
  NAND2X1 U31818 ( .A(n31282), .B(n31283), .Y(n31281) );
  AND2X1 U31837 ( .A(n31302), .B(n31303), .Y(n31289) );
  NOR2X1 U31845 ( .A(n31308), .B(n31309), .Y(n31302) );
  NAND2X1 U31854 ( .A(n31316), .B(n31317), .Y(n31280) );
  NOR2X1 U31862 ( .A(n31322), .B(n31323), .Y(n31316) );
  NOR2X1 U31871 ( .A(n31330), .B(n31331), .Y(n31278) );
  NAND2X1 U31878 ( .A(n31337), .B(n31338), .Y(n31276) );
  NOR2X1 U31886 ( .A(n31343), .B(n31344), .Y(n31337) );
  NOR2X1 U31895 ( .A(n31351), .B(n31352), .Y(n31274) );
  NAND2X1 U31900 ( .A(n31357), .B(n31358), .Y(n31272) );
  NOR2X1 U31908 ( .A(n31363), .B(n31364), .Y(n31357) );
  NOR2X1 U31917 ( .A(n31371), .B(n31372), .Y(n31270) );
  NAND2X1 U31923 ( .A(n31377), .B(n31378), .Y(n31268) );
  NOR2X1 U31931 ( .A(n31383), .B(n31384), .Y(n31377) );
  NAND2X1 U31943 ( .A(n31394), .B(n31395), .Y(n31153) );
  NOR2X1 U31951 ( .A(n31400), .B(n31401), .Y(n31394) );
  NOR2X1 U31961 ( .A(n31409), .B(n31410), .Y(n31146) );
  NAND2X1 U31962 ( .A(n31411), .B(n31412), .Y(n31410) );
  NAND2X1 U31978 ( .A(n31423), .B(n31424), .Y(n31134) );
  NOR2X1 U32003 ( .A(n31444), .B(n31445), .Y(n31132) );
  NAND2X1 U32011 ( .A(n31450), .B(n31451), .Y(n31444) );
  NAND2X1 U32024 ( .A(n31462), .B(n31463), .Y(n31461) );
  NOR2X1 U32025 ( .A(n31464), .B(n31465), .Y(n31463) );
  NAND2X1 U32165 ( .A(n31653), .B(n31654), .Y(n31464) );
  NOR2X1 U32306 ( .A(n31786), .B(n31787), .Y(n31462) );
  NOR2X1 U32443 ( .A(n31923), .B(n395), .Y(n31922) );
  NOR2X1 U32532 ( .A(n32009), .B(n430), .Y(n32008) );
  NOR2X1 U32533 ( .A(n581), .B(n73552), .Y(n32007) );
  NOR2X1 U32535 ( .A(n577), .B(n438), .Y(n32011) );
  AND2X1 U32536 ( .A(n583), .B(mem_d_data_rd_i[25]), .Y(n32010) );
  NAND2X1 U32728 ( .A(n32196), .B(n32197), .Y(n31460) );
  NOR2X1 U32729 ( .A(n32198), .B(n32199), .Y(n32197) );
  NOR2X1 U32869 ( .A(n47178), .B(n430), .Y(n32333) );
  NAND2X1 U32871 ( .A(n73435), .B(n32335), .Y(n32198) );
  NOR2X1 U33012 ( .A(n32467), .B(n32468), .Y(n32196) );
  NAND2X1 U33024 ( .A(n32473), .B(n32474), .Y(n32472) );
  NOR2X1 U33025 ( .A(n32475), .B(n32476), .Y(n32474) );
  NAND2X1 U33026 ( .A(n32477), .B(n73434), .Y(n32476) );
  NOR2X1 U33030 ( .A(n31408), .B(n31391), .Y(n32477) );
  NOR2X1 U33168 ( .A(n31923), .B(n384), .Y(n32610) );
  NOR2X1 U33305 ( .A(n31923), .B(n373), .Y(n32743) );
  NAND2X1 U33309 ( .A(n32744), .B(n73436), .Y(n32475) );
  NOR2X1 U33313 ( .A(n31152), .B(n31393), .Y(n32744) );
  NOR2X1 U33856 ( .A(n33270), .B(n33271), .Y(n32473) );
  AND2X1 U34128 ( .A(n584), .B(mem_d_data_rd_i[12]), .Y(n33540) );
  NOR2X1 U34129 ( .A(n581), .B(n73549), .Y(n33539) );
  NOR2X1 U34131 ( .A(n33543), .B(n373), .Y(n33542) );
  NOR2X1 U34132 ( .A(n577), .B(n432), .Y(n33541) );
  NAND2X1 U34268 ( .A(mem_d_data_rd_i[5]), .B(n33678), .Y(n33677) );
  NAND2X1 U34269 ( .A(mem_d_data_rd_i[29]), .B(n583), .Y(n33676) );
  NAND2X1 U34271 ( .A(mem_d_data_rd_i[21]), .B(n33681), .Y(n33680) );
  NAND2X1 U34272 ( .A(mem_d_data_rd_i[13]), .B(n584), .Y(n33679) );
  AND2X1 U34680 ( .A(n584), .B(mem_d_data_rd_i[11]), .Y(n34081) );
  NOR2X1 U34681 ( .A(n581), .B(n73550), .Y(n34080) );
  NOR2X1 U34683 ( .A(n33543), .B(n384), .Y(n34083) );
  NOR2X1 U34684 ( .A(n577), .B(n436), .Y(n34082) );
  NAND2X1 U34686 ( .A(n34084), .B(n34085), .Y(n32471) );
  NOR2X1 U34687 ( .A(n34086), .B(n34087), .Y(n34085) );
  AND2X1 U34824 ( .A(n73578), .B(mem_d_data_rd_i[29]), .Y(n34221) );
  AND2X1 U34963 ( .A(n73578), .B(mem_d_data_rd_i[30]), .Y(n34356) );
  NAND2X1 U35100 ( .A(n34491), .B(n34492), .Y(n34086) );
  NOR2X1 U35238 ( .A(n47178), .B(n431), .Y(n34625) );
  NAND2X1 U35374 ( .A(mem_d_data_rd_i[6]), .B(n33678), .Y(n34759) );
  NAND2X1 U35375 ( .A(mem_d_data_rd_i[30]), .B(n583), .Y(n34758) );
  NAND2X1 U35377 ( .A(mem_d_data_rd_i[22]), .B(n33681), .Y(n34761) );
  NAND2X1 U35378 ( .A(mem_d_data_rd_i[14]), .B(n584), .Y(n34760) );
  NOR2X1 U35650 ( .A(n429), .B(n32009), .Y(n35027) );
  AND2X1 U35651 ( .A(n33681), .B(mem_d_data_rd_i[23]), .Y(n35026) );
  AND2X1 U35653 ( .A(mem_d_data_rd_i[31]), .B(n583), .Y(n35029) );
  AND2X1 U35654 ( .A(n33678), .B(mem_d_data_rd_i[7]), .Y(n35028) );
  NOR2X1 U35655 ( .A(n35030), .B(n35031), .Y(n34084) );
  AND2X1 U35792 ( .A(n584), .B(mem_d_data_rd_i[10]), .Y(n35166) );
  NOR2X1 U35793 ( .A(n581), .B(n73551), .Y(n35165) );
  NOR2X1 U35795 ( .A(n33543), .B(n395), .Y(n35168) );
  NOR2X1 U35796 ( .A(n577), .B(n437), .Y(n35167) );
  NOR2X1 U35932 ( .A(n431), .B(n32009), .Y(n35304) );
  NAND2X1 U35933 ( .A(n35305), .B(mem_d_resp_tag_i[5]), .Y(n32009) );
  NOR2X1 U35934 ( .A(mem_d_resp_tag_i[6]), .B(n585), .Y(n35305) );
  NOR2X1 U35935 ( .A(n581), .B(n73553), .Y(n35303) );
  NAND2X1 U35936 ( .A(n31923), .B(n35306), .Y(n33681) );
  NAND2X1 U35937 ( .A(n35307), .B(mem_d_resp_tag_i[6]), .Y(n35306) );
  NOR2X1 U35938 ( .A(mem_d_resp_tag_i[5]), .B(n585), .Y(n35307) );
  NOR2X1 U35940 ( .A(n577), .B(n73554), .Y(n35309) );
  NAND2X1 U35941 ( .A(n47178), .B(n35310), .Y(n33678) );
  NAND2X1 U35942 ( .A(n587), .B(n586), .Y(n35310) );
  NAND2X1 U35943 ( .A(n29623), .B(n35311), .Y(n31921) );
  NAND2X1 U35944 ( .A(n586), .B(n585), .Y(n35311) );
  AND2X1 U35945 ( .A(mem_d_data_rd_i[24]), .B(n583), .Y(n35308) );
  NAND2X1 U35946 ( .A(n35312), .B(mem_d_resp_tag_i[5]), .Y(n33543) );
  NOR2X1 U35947 ( .A(n585), .B(n586), .Y(n35312) );
  NAND2X1 U36534 ( .A(mem_d_resp_tag_i[10]), .B(n35892), .Y(n35891) );
  NAND2X1 U36535 ( .A(n34490), .B(n35893), .Y(n35892) );
  NAND2X1 U36536 ( .A(n35894), .B(n35895), .Y(n35893) );
  NOR2X1 U36537 ( .A(mem_d_resp_tag_i[7]), .B(mem_d_resp_tag_i[6]), .Y(n35895)
         );
  NOR2X1 U36538 ( .A(n582), .B(n429), .Y(n35894) );
  NAND2X1 U36539 ( .A(mem_d_data_rd_i[31]), .B(n73578), .Y(n34490) );
  NAND2X1 U36540 ( .A(n35896), .B(mem_d_resp_tag_i[6]), .Y(n31923) );
  NOR2X1 U36541 ( .A(mem_d_resp_tag_i[7]), .B(n582), .Y(n35896) );
  NAND2X1 U36542 ( .A(n35897), .B(n35898), .Y(n34489) );
  NOR2X1 U36543 ( .A(n35899), .B(n35900), .Y(n35898) );
  NOR2X1 U36544 ( .A(n35901), .B(n586), .Y(n35900) );
  NOR2X1 U36545 ( .A(n35902), .B(n35903), .Y(n35901) );
  NOR2X1 U36546 ( .A(mem_d_data_rd_i[31]), .B(n587), .Y(n35903) );
  NOR2X1 U36547 ( .A(mem_d_resp_tag_i[5]), .B(mem_d_data_rd_i[23]), .Y(n35902)
         );
  NOR2X1 U36548 ( .A(mem_d_resp_tag_i[6]), .B(n35904), .Y(n35899) );
  NOR2X1 U36549 ( .A(n35905), .B(n35906), .Y(n35904) );
  NOR2X1 U36550 ( .A(mem_d_resp_tag_i[5]), .B(mem_d_data_rd_i[7]), .Y(n35906)
         );
  NOR2X1 U36551 ( .A(mem_d_data_rd_i[15]), .B(n587), .Y(n35905) );
  AND2X1 U36552 ( .A(mem_d_resp_tag_i[7]), .B(mem_d_resp_tag_i[10]), .Y(n35897) );
  NAND2X1 U36596 ( .A(u_arb_src_mmu_q), .B(u_arb_read_hold_q), .Y(n35938) );
  NAND2X1 U36620 ( .A(n35952), .B(n8417), .Y(n35956) );
  NAND2X1 U36621 ( .A(n35957), .B(n35958), .Y(n35952) );
  NAND2X1 U36622 ( .A(n35959), .B(u_csr_N3161), .Y(n35958) );
  NAND2X1 U36623 ( .A(u_mmu_dtlb_entry_q_4), .B(n8835), .Y(n35959) );
  NAND2X1 U36624 ( .A(n73569), .B(u_mmu_dtlb_entry_q_4), .Y(n35957) );
  NAND2X1 U36646 ( .A(n35981), .B(n35982), .Y(n35970) );
  NAND2X1 U36647 ( .A(n35983), .B(u_decode_scoreboard_q[5]), .Y(n35982) );
  NAND2X1 U36653 ( .A(n35987), .B(n35988), .Y(n35981) );
  NAND2X1 U36654 ( .A(n35989), .B(n35990), .Y(n35988) );
  OR2X1 U36655 ( .A(n35991), .B(n569), .Y(n35990) );
  NAND2X1 U36656 ( .A(n73427), .B(n40841), .Y(n24134) );
  NAND2X1 U36661 ( .A(n553), .B(n35991), .Y(n35987) );
  NAND2X1 U36666 ( .A(n73427), .B(n35997), .Y(n24179) );
  NAND2X1 U36668 ( .A(n36000), .B(n36001), .Y(n35999) );
  NAND2X1 U36669 ( .A(n36002), .B(u_decode_scoreboard_q[18]), .Y(n36001) );
  NAND2X1 U36675 ( .A(n36006), .B(u_decode_scoreboard_q[28]), .Y(n36000) );
  AND2X1 U36727 ( .A(u_decode_scoreboard_q[24]), .B(n18296), .Y(n24239) );
  NAND2X1 U36728 ( .A(n36009), .B(n35922), .Y(n18296) );
  AND2X1 U36730 ( .A(u_decode_scoreboard_q[8]), .B(n21437), .Y(n24125) );
  AND2X1 U36735 ( .A(u_decode_scoreboard_q[17]), .B(n19670), .Y(n24298) );
  NAND2X1 U36736 ( .A(n40938), .B(n35922), .Y(n19670) );
  NAND2X1 U36856 ( .A(n73526), .B(n40938), .Y(n24263) );
  NOR2X1 U36858 ( .A(mem_d_resp_tag_i[3]), .B(n73557), .Y(n36163) );
  NAND2X1 U36876 ( .A(n36176), .B(n36177), .Y(n36175) );
  NAND2X1 U36877 ( .A(n36178), .B(u_decode_scoreboard_q[22]), .Y(n36177) );
  NAND2X1 U36883 ( .A(n36180), .B(u_decode_scoreboard_q[20]), .Y(n36176) );
  NAND2X1 U36914 ( .A(u_decode_scoreboard_q[25]), .B(n24101), .Y(n24229) );
  NAND2X1 U36915 ( .A(n35997), .B(n35922), .Y(n24101) );
  AND2X1 U36916 ( .A(n36197), .B(mem_d_resp_tag_i[0]), .Y(n35997) );
  NAND2X1 U36917 ( .A(n36198), .B(n36199), .Y(n36191) );
  NAND2X1 U36918 ( .A(n36200), .B(u_decode_scoreboard_q[10]), .Y(n36199) );
  NAND2X1 U36924 ( .A(n36202), .B(u_decode_scoreboard_q[6]), .Y(n36198) );
  NOR2X1 U36936 ( .A(n36208), .B(n36209), .Y(n36207) );
  NAND2X1 U36937 ( .A(n36210), .B(n36211), .Y(n36209) );
  NAND2X1 U36938 ( .A(n36212), .B(u_decode_scoreboard_q[11]), .Y(n36211) );
  NAND2X1 U36948 ( .A(n36217), .B(u_decode_scoreboard_q[26]), .Y(n36210) );
  AND2X1 U36956 ( .A(n36197), .B(n73557), .Y(n36009) );
  AND2X1 U36957 ( .A(mem_d_resp_tag_i[3]), .B(n73527), .Y(n36197) );
  NAND2X1 U36958 ( .A(n36219), .B(n36220), .Y(n36208) );
  NAND2X1 U36959 ( .A(n36221), .B(u_decode_scoreboard_q[4]), .Y(n36220) );
  AND2X1 U36973 ( .A(u_decode_scoreboard_q[16]), .B(n19867), .Y(n24306) );
  NAND2X1 U36974 ( .A(n73421), .B(n35922), .Y(n19867) );
  NOR2X1 U36977 ( .A(mem_d_resp_tag_i[3]), .B(mem_d_resp_tag_i[0]), .Y(n36227)
         );
  NAND2X1 U36996 ( .A(u_decode_scoreboard_q[1]), .B(n24109), .Y(n24275) );
  NAND2X1 U37000 ( .A(n36238), .B(n36239), .Y(n36228) );
  NAND2X1 U37001 ( .A(n36240), .B(u_decode_scoreboard_q[2]), .Y(n36239) );
  NAND2X1 U37014 ( .A(n36237), .B(n73557), .Y(n36244) );
  NOR2X1 U37015 ( .A(mem_d_resp_tag_i[4]), .B(mem_d_resp_tag_i[3]), .Y(n36237)
         );
  AND2X1 U37028 ( .A(u_decode_scoreboard_q[9]), .B(n21240), .Y(n24117) );
  NAND2X1 U37029 ( .A(n40937), .B(n35922), .Y(n21240) );
  NAND2X1 U37031 ( .A(n73556), .B(n73555), .Y(n36247) );
  NAND2X1 U37035 ( .A(n36250), .B(n36251), .Y(n36249) );
  OR2X1 U37036 ( .A(n576), .B(n30272), .Y(n36251) );
  NOR2X1 U37037 ( .A(n582), .B(n585), .Y(n30272) );
  NAND2X1 U37038 ( .A(n29623), .B(n576), .Y(n36250) );
  NAND2X1 U37039 ( .A(n582), .B(n585), .Y(n29623) );
  NOR2X1 U37040 ( .A(mem_d_resp_tag_i[4]), .B(n73557), .Y(n36248) );
  NOR2X1 \clk_gate_u_mmu_dtlb_entry_q_reg/U2  ( .A(
        \clk_gate_u_mmu_dtlb_entry_q_reg/n2 ), .B(n73546), .Y(net1782) );
  TLATX1 \clk_gate_u_mmu_dtlb_entry_q_reg/latch  ( .G(n73546), .D(n17208), 
        .QN(\clk_gate_u_mmu_dtlb_entry_q_reg/n2 ) );
  TLATX1 \clk_gate_u_mmu_dtlb_entry_q_reg_0/latch  ( .G(n73546), .D(n17209), 
        .QN(\clk_gate_u_mmu_dtlb_entry_q_reg_0/n2 ) );
  NOR2X1 \clk_gate_u_mmu_itlb_entry_q_reg/U2  ( .A(
        \clk_gate_u_mmu_itlb_entry_q_reg/n2 ), .B(n73546), .Y(net1792) );
  TLATX1 \clk_gate_u_mmu_itlb_entry_q_reg/latch  ( .G(n73546), .D(n17210), 
        .QN(\clk_gate_u_mmu_itlb_entry_q_reg/n2 ) );
  TLATX1 \clk_gate_u_mmu_itlb_entry_q_reg_0/latch  ( .G(n73546), .D(n17211), 
        .QN(\clk_gate_u_mmu_itlb_entry_q_reg_0/n2 ) );
  NOR2X1 \clk_gate_u_mmu_pte_entry_q_reg/U2  ( .A(
        \clk_gate_u_mmu_pte_entry_q_reg/n2 ), .B(n73546), .Y(net1802) );
  TLATX1 \clk_gate_u_mmu_pte_entry_q_reg/latch  ( .G(n73546), .D(n17212), .QN(
        \clk_gate_u_mmu_pte_entry_q_reg/n2 ) );
  TLATX1 \clk_gate_u_mmu_pte_addr_q_reg/latch  ( .G(n73546), .D(n17213), .QN(
        \clk_gate_u_mmu_pte_addr_q_reg/n2 ) );
  TLATX1 \clk_gate_u_mmu_pte_addr_q_reg_0/latch  ( .G(n73546), .D(n17214), 
        .QN(\clk_gate_u_mmu_pte_addr_q_reg_0/n2 ) );
  TLATX1 \clk_gate_u_mmu_virt_addr_q_reg/latch  ( .G(n73546), .D(n17215), .QN(
        \clk_gate_u_mmu_virt_addr_q_reg/n2 ) );
  TLATX1 \clk_gate_u_mmu_lsu_in_addr_q_reg/latch  ( .G(n73546), .D(n17216), 
        .QN(\clk_gate_u_mmu_lsu_in_addr_q_reg/n2 ) );
  TLATX1 \clk_gate_u_mmu_lsu_in_addr_q_reg_0/latch  ( .G(n73546), .D(n17217), 
        .QN(\clk_gate_u_mmu_lsu_in_addr_q_reg_0/n2 ) );
  TLATX1 \clk_gate_u_lsu_mem_cacheable_q_reg/latch  ( .G(n73546), .D(n17218), 
        .QN(\clk_gate_u_lsu_mem_cacheable_q_reg/n2 ) );
  TLATX1 \clk_gate_u_lsu_mem_addr_q_reg/latch  ( .G(n73546), .D(n17219), .QN(
        \clk_gate_u_lsu_mem_addr_q_reg/n2 ) );
  TLATX1 \clk_gate_u_lsu_mem_addr_q_reg_0/latch  ( .G(n73546), .D(n17220), 
        .QN(\clk_gate_u_lsu_mem_addr_q_reg_0/n2 ) );
  NOR2X1 \clk_gate_u_lsu_mem_data_wr_q_reg/U2  ( .A(
        \clk_gate_u_lsu_mem_data_wr_q_reg/n2 ), .B(n73546), .Y(net1847) );
  TLATX1 \clk_gate_u_lsu_mem_data_wr_q_reg/latch  ( .G(n73546), .D(n17221), 
        .QN(\clk_gate_u_lsu_mem_data_wr_q_reg/n2 ) );
  TLATX1 \clk_gate_u_lsu_mem_data_wr_q_reg_0/latch  ( .G(n73546), .D(n17222), 
        .QN(\clk_gate_u_lsu_mem_data_wr_q_reg_0/n2 ) );
  NOR2X1 \clk_gate_u_csr_writeback_value_q_reg/U2  ( .A(
        \clk_gate_u_csr_writeback_value_q_reg/n2 ), .B(n73546), .Y(net1857) );
  TLATX1 \clk_gate_u_csr_writeback_value_q_reg/latch  ( .G(n73546), .D(n17223), 
        .QN(\clk_gate_u_csr_writeback_value_q_reg/n2 ) );
  NOR2X1 \clk_gate_u_csr_writeback_value_q_reg_0/U2  ( .A(
        \clk_gate_u_csr_writeback_value_q_reg_0/n2 ), .B(n73546), .Y(net1862)
         );
  TLATX1 \clk_gate_u_csr_writeback_value_q_reg_0/latch  ( .G(n73546), .D(
        n17224), .QN(\clk_gate_u_csr_writeback_value_q_reg_0/n2 ) );
  NOR2X1 \clk_gate_u_csr_writeback_idx_q_reg/U2  ( .A(
        \clk_gate_u_csr_writeback_idx_q_reg/n2 ), .B(n73546), .Y(net1867) );
  TLATX1 \clk_gate_u_csr_writeback_idx_q_reg/latch  ( .G(n73546), .D(n17225), 
        .QN(\clk_gate_u_csr_writeback_idx_q_reg/n2 ) );
  NOR2X1 \clk_gate_u_csr_pc_m_q_reg/U2  ( .A(\clk_gate_u_csr_pc_m_q_reg/n2 ), 
        .B(n73546), .Y(net1872) );
  TLATX1 \clk_gate_u_csr_pc_m_q_reg/latch  ( .G(n73546), .D(n17226), .QN(
        \clk_gate_u_csr_pc_m_q_reg/n2 ) );
  NOR2X1 \clk_gate_u_csr_csr_sr_q_reg/U2  ( .A(
        \clk_gate_u_csr_csr_sr_q_reg/n2 ), .B(n73546), .Y(net1878) );
  TLATX1 \clk_gate_u_csr_csr_sr_q_reg/latch  ( .G(n73546), .D(n17227), .QN(
        \clk_gate_u_csr_csr_sr_q_reg/n2 ) );
  NOR2X1 \clk_gate_u_muldiv_divisor_q_reg/U2  ( .A(
        \clk_gate_u_muldiv_divisor_q_reg/n2 ), .B(n73546), .Y(net1883) );
  TLATX1 \clk_gate_u_muldiv_divisor_q_reg/latch  ( .G(n73546), .D(n17228), 
        .QN(\clk_gate_u_muldiv_divisor_q_reg/n2 ) );
  NOR2X1 \clk_gate_u_muldiv_divisor_q_reg_0/U2  ( .A(
        \clk_gate_u_muldiv_divisor_q_reg_0/n2 ), .B(n73546), .Y(net1888) );
  TLATX1 \clk_gate_u_muldiv_divisor_q_reg_0/latch  ( .G(n73546), .D(n17229), 
        .QN(\clk_gate_u_muldiv_divisor_q_reg_0/n2 ) );
  NOR2X1 \clk_gate_u_muldiv_divisor_q_reg_1/U2  ( .A(
        \clk_gate_u_muldiv_divisor_q_reg_1/n2 ), .B(n73546), .Y(net1893) );
  TLATX1 \clk_gate_u_muldiv_divisor_q_reg_1/latch  ( .G(n73546), .D(n17230), 
        .QN(\clk_gate_u_muldiv_divisor_q_reg_1/n2 ) );
  NOR2X1 \clk_gate_u_muldiv_divisor_q_reg_2/U2  ( .A(
        \clk_gate_u_muldiv_divisor_q_reg_2/n2 ), .B(n73546), .Y(net1898) );
  TLATX1 \clk_gate_u_muldiv_divisor_q_reg_2/latch  ( .G(n73546), .D(n17231), 
        .QN(\clk_gate_u_muldiv_divisor_q_reg_2/n2 ) );
  NOR2X1 \clk_gate_u_muldiv_q_mask_q_reg/U2  ( .A(
        \clk_gate_u_muldiv_q_mask_q_reg/n2 ), .B(n73546), .Y(net1903) );
  TLATX1 \clk_gate_u_muldiv_q_mask_q_reg/latch  ( .G(n73546), .D(n17232), .QN(
        \clk_gate_u_muldiv_q_mask_q_reg/n2 ) );
  NOR2X1 \clk_gate_u_muldiv_dividend_q_reg/U2  ( .A(
        \clk_gate_u_muldiv_dividend_q_reg/n2 ), .B(n73546), .Y(net1908) );
  TLATX1 \clk_gate_u_muldiv_dividend_q_reg/latch  ( .G(n73546), .D(n17233), 
        .QN(\clk_gate_u_muldiv_dividend_q_reg/n2 ) );
  NOR2X1 \clk_gate_u_muldiv_dividend_q_reg_0/U2  ( .A(
        \clk_gate_u_muldiv_dividend_q_reg_0/n2 ), .B(n73546), .Y(net1913) );
  TLATX1 \clk_gate_u_muldiv_dividend_q_reg_0/latch  ( .G(n73546), .D(n17234), 
        .QN(\clk_gate_u_muldiv_dividend_q_reg_0/n2 ) );
  NOR2X1 \clk_gate_u_muldiv_quotient_q_reg/U2  ( .A(
        \clk_gate_u_muldiv_quotient_q_reg/n2 ), .B(n73546), .Y(net1918) );
  TLATX1 \clk_gate_u_muldiv_quotient_q_reg/latch  ( .G(n73546), .D(n17235), 
        .QN(\clk_gate_u_muldiv_quotient_q_reg/n2 ) );
  NOR2X1 \clk_gate_u_muldiv_quotient_q_reg_0/U2  ( .A(
        \clk_gate_u_muldiv_quotient_q_reg_0/n2 ), .B(n73546), .Y(net1923) );
  TLATX1 \clk_gate_u_muldiv_quotient_q_reg_0/latch  ( .G(n73546), .D(n17236), 
        .QN(\clk_gate_u_muldiv_quotient_q_reg_0/n2 ) );
  TLATX1 \clk_gate_u_decode_opcode_instr_q_reg/latch  ( .G(n73546), .D(n17237), 
        .QN(\clk_gate_u_decode_opcode_instr_q_reg/n2 ) );
  TLATX1 \clk_gate_u_decode_opcode_instr_q_reg_0/latch  ( .G(n73546), .D(
        n17238), .QN(\clk_gate_u_decode_opcode_instr_q_reg_0/n2 ) );
  TLATX1 \clk_gate_u_decode_opcode_instr_q_reg_1/latch  ( .G(n73546), .D(
        n17239), .QN(\clk_gate_u_decode_opcode_instr_q_reg_1/n2 ) );
  TLATX1 \clk_gate_u_decode_opcode_instr_q_reg_2/latch  ( .G(n73546), .D(
        n17240), .QN(\clk_gate_u_decode_opcode_instr_q_reg_2/n2 ) );
  TLATX1 \clk_gate_u_decode_inst_q_reg/latch  ( .G(n73546), .D(n17241), .QN(
        \clk_gate_u_decode_inst_q_reg/n2 ) );
  TLATX1 \clk_gate_u_decode_pc_q_reg/latch  ( .G(n73546), .D(n17242), .QN(
        \clk_gate_u_decode_pc_q_reg/n2 ) );
  TLATX1 \clk_gate_u_decode_pc_q_reg_0/latch  ( .G(n73546), .D(n17243), .QN(
        \clk_gate_u_decode_pc_q_reg_0/n2 ) );
  TLATX1 \clk_gate_u_decode_u_regfile_reg_r21_q_reg/latch  ( .G(n73546), .D(
        n17244), .QN(\clk_gate_u_decode_u_regfile_reg_r21_q_reg/n2 ) );
  TLATX1 \clk_gate_u_decode_u_regfile_reg_r21_q_reg_0/latch  ( .G(n73546), .D(
        n17245), .QN(\clk_gate_u_decode_u_regfile_reg_r21_q_reg_0/n2 ) );
  TLATX1 \clk_gate_u_decode_u_regfile_reg_r20_q_reg/latch  ( .G(n73546), .D(
        n17246), .QN(\clk_gate_u_decode_u_regfile_reg_r20_q_reg/n2 ) );
  TLATX1 \clk_gate_u_decode_u_regfile_reg_r20_q_reg_0/latch  ( .G(n73546), .D(
        n17247), .QN(\clk_gate_u_decode_u_regfile_reg_r20_q_reg_0/n2 ) );
  TLATX1 \clk_gate_u_decode_u_regfile_reg_r19_q_reg/latch  ( .G(n73546), .D(
        n17248), .QN(\clk_gate_u_decode_u_regfile_reg_r19_q_reg/n2 ) );
  TLATX1 \clk_gate_u_decode_u_regfile_reg_r19_q_reg_0/latch  ( .G(n73546), .D(
        n17249), .QN(\clk_gate_u_decode_u_regfile_reg_r19_q_reg_0/n2 ) );
  TLATX1 \clk_gate_u_decode_u_regfile_reg_r18_q_reg/latch  ( .G(n73546), .D(
        n17250), .QN(\clk_gate_u_decode_u_regfile_reg_r18_q_reg/n2 ) );
  TLATX1 \clk_gate_u_decode_u_regfile_reg_r18_q_reg_0/latch  ( .G(n73546), .D(
        n17251), .QN(\clk_gate_u_decode_u_regfile_reg_r18_q_reg_0/n2 ) );
  TLATX1 \clk_gate_u_decode_u_regfile_reg_r17_q_reg/latch  ( .G(n73546), .D(
        n17252), .QN(\clk_gate_u_decode_u_regfile_reg_r17_q_reg/n2 ) );
  TLATX1 \clk_gate_u_decode_u_regfile_reg_r17_q_reg_0/latch  ( .G(n73546), .D(
        n17253), .QN(\clk_gate_u_decode_u_regfile_reg_r17_q_reg_0/n2 ) );
  TLATX1 \clk_gate_u_decode_u_regfile_reg_r16_q_reg/latch  ( .G(n73546), .D(
        n17254), .QN(\clk_gate_u_decode_u_regfile_reg_r16_q_reg/n2 ) );
  TLATX1 \clk_gate_u_decode_u_regfile_reg_r16_q_reg_0/latch  ( .G(n73546), .D(
        n17255), .QN(\clk_gate_u_decode_u_regfile_reg_r16_q_reg_0/n2 ) );
  TLATX1 \clk_gate_u_decode_u_regfile_reg_r15_q_reg/latch  ( .G(n73546), .D(
        n17256), .QN(\clk_gate_u_decode_u_regfile_reg_r15_q_reg/n2 ) );
  TLATX1 \clk_gate_u_decode_u_regfile_reg_r15_q_reg_0/latch  ( .G(n73546), .D(
        n17257), .QN(\clk_gate_u_decode_u_regfile_reg_r15_q_reg_0/n2 ) );
  TLATX1 \clk_gate_u_decode_u_regfile_reg_r14_q_reg/latch  ( .G(n73546), .D(
        n17258), .QN(\clk_gate_u_decode_u_regfile_reg_r14_q_reg/n2 ) );
  TLATX1 \clk_gate_u_decode_u_regfile_reg_r14_q_reg_0/latch  ( .G(n73546), .D(
        n17259), .QN(\clk_gate_u_decode_u_regfile_reg_r14_q_reg_0/n2 ) );
  TLATX1 \clk_gate_u_decode_u_regfile_reg_r13_q_reg/latch  ( .G(n73546), .D(
        n17260), .QN(\clk_gate_u_decode_u_regfile_reg_r13_q_reg/n2 ) );
  TLATX1 \clk_gate_u_decode_u_regfile_reg_r13_q_reg_0/latch  ( .G(n73546), .D(
        n17261), .QN(\clk_gate_u_decode_u_regfile_reg_r13_q_reg_0/n2 ) );
  TLATX1 \clk_gate_u_decode_u_regfile_reg_r12_q_reg/latch  ( .G(n73546), .D(
        n17262), .QN(\clk_gate_u_decode_u_regfile_reg_r12_q_reg/n2 ) );
  TLATX1 \clk_gate_u_decode_u_regfile_reg_r12_q_reg_0/latch  ( .G(n73546), .D(
        n17263), .QN(\clk_gate_u_decode_u_regfile_reg_r12_q_reg_0/n2 ) );
  TLATX1 \clk_gate_u_decode_u_regfile_reg_r11_q_reg/latch  ( .G(n73546), .D(
        n17264), .QN(\clk_gate_u_decode_u_regfile_reg_r11_q_reg/n2 ) );
  TLATX1 \clk_gate_u_decode_u_regfile_reg_r11_q_reg_0/latch  ( .G(n73546), .D(
        n17265), .QN(\clk_gate_u_decode_u_regfile_reg_r11_q_reg_0/n2 ) );
  TLATX1 \clk_gate_u_decode_u_regfile_reg_r10_q_reg/latch  ( .G(n73546), .D(
        n17266), .QN(\clk_gate_u_decode_u_regfile_reg_r10_q_reg/n2 ) );
  TLATX1 \clk_gate_u_decode_u_regfile_reg_r10_q_reg_0/latch  ( .G(n73546), .D(
        n17267), .QN(\clk_gate_u_decode_u_regfile_reg_r10_q_reg_0/n2 ) );
  TLATX1 \clk_gate_u_decode_u_regfile_reg_r9_q_reg/latch  ( .G(n73546), .D(
        n17268), .QN(\clk_gate_u_decode_u_regfile_reg_r9_q_reg/n2 ) );
  TLATX1 \clk_gate_u_decode_u_regfile_reg_r9_q_reg_0/latch  ( .G(n73546), .D(
        n17269), .QN(\clk_gate_u_decode_u_regfile_reg_r9_q_reg_0/n2 ) );
  TLATX1 \clk_gate_u_decode_u_regfile_reg_r8_q_reg/latch  ( .G(n73546), .D(
        n17270), .QN(\clk_gate_u_decode_u_regfile_reg_r8_q_reg/n2 ) );
  TLATX1 \clk_gate_u_decode_u_regfile_reg_r8_q_reg_0/latch  ( .G(n73546), .D(
        n17271), .QN(\clk_gate_u_decode_u_regfile_reg_r8_q_reg_0/n2 ) );
  TLATX1 \clk_gate_u_decode_u_regfile_reg_r7_q_reg/latch  ( .G(n73546), .D(
        n17272), .QN(\clk_gate_u_decode_u_regfile_reg_r7_q_reg/n2 ) );
  TLATX1 \clk_gate_u_decode_u_regfile_reg_r7_q_reg_0/latch  ( .G(n73546), .D(
        n17273), .QN(\clk_gate_u_decode_u_regfile_reg_r7_q_reg_0/n2 ) );
  TLATX1 \clk_gate_u_decode_u_regfile_reg_r6_q_reg/latch  ( .G(n73546), .D(
        n17274), .QN(\clk_gate_u_decode_u_regfile_reg_r6_q_reg/n2 ) );
  TLATX1 \clk_gate_u_decode_u_regfile_reg_r6_q_reg_0/latch  ( .G(n73546), .D(
        n17275), .QN(\clk_gate_u_decode_u_regfile_reg_r6_q_reg_0/n2 ) );
  TLATX1 \clk_gate_u_decode_u_regfile_reg_r5_q_reg/latch  ( .G(n73546), .D(
        n17276), .QN(\clk_gate_u_decode_u_regfile_reg_r5_q_reg/n2 ) );
  TLATX1 \clk_gate_u_decode_u_regfile_reg_r5_q_reg_0/latch  ( .G(n73546), .D(
        n17277), .QN(\clk_gate_u_decode_u_regfile_reg_r5_q_reg_0/n2 ) );
  TLATX1 \clk_gate_u_decode_u_regfile_reg_r4_q_reg/latch  ( .G(n73546), .D(
        n17278), .QN(\clk_gate_u_decode_u_regfile_reg_r4_q_reg/n2 ) );
  TLATX1 \clk_gate_u_decode_u_regfile_reg_r4_q_reg_0/latch  ( .G(n73546), .D(
        n17279), .QN(\clk_gate_u_decode_u_regfile_reg_r4_q_reg_0/n2 ) );
  TLATX1 \clk_gate_u_decode_u_regfile_reg_r3_q_reg/latch  ( .G(n73546), .D(
        n17280), .QN(\clk_gate_u_decode_u_regfile_reg_r3_q_reg/n2 ) );
  TLATX1 \clk_gate_u_decode_u_regfile_reg_r3_q_reg_0/latch  ( .G(n73546), .D(
        n17281), .QN(\clk_gate_u_decode_u_regfile_reg_r3_q_reg_0/n2 ) );
  TLATX1 \clk_gate_u_decode_u_regfile_reg_r2_q_reg/latch  ( .G(n73546), .D(
        n17282), .QN(\clk_gate_u_decode_u_regfile_reg_r2_q_reg/n2 ) );
  TLATX1 \clk_gate_u_decode_u_regfile_reg_r2_q_reg_0/latch  ( .G(n73546), .D(
        n17283), .QN(\clk_gate_u_decode_u_regfile_reg_r2_q_reg_0/n2 ) );
  TLATX1 \clk_gate_u_decode_u_regfile_reg_r1_q_reg/latch  ( .G(n73546), .D(
        n17284), .QN(\clk_gate_u_decode_u_regfile_reg_r1_q_reg/n2 ) );
  TLATX1 \clk_gate_u_decode_u_regfile_reg_r1_q_reg_0/latch  ( .G(n73546), .D(
        n17285), .QN(\clk_gate_u_decode_u_regfile_reg_r1_q_reg_0/n2 ) );
  TLATX1 \clk_gate_u_decode_u_regfile_reg_r31_q_reg/latch  ( .G(n73546), .D(
        n17286), .QN(\clk_gate_u_decode_u_regfile_reg_r31_q_reg/n2 ) );
  TLATX1 \clk_gate_u_decode_u_regfile_reg_r31_q_reg_0/latch  ( .G(n73546), .D(
        n17287), .QN(\clk_gate_u_decode_u_regfile_reg_r31_q_reg_0/n2 ) );
  TLATX1 \clk_gate_u_decode_u_regfile_reg_r26_q_reg/latch  ( .G(n73546), .D(
        n17288), .QN(\clk_gate_u_decode_u_regfile_reg_r26_q_reg/n2 ) );
  TLATX1 \clk_gate_u_decode_u_regfile_reg_r26_q_reg_0/latch  ( .G(n73546), .D(
        n17289), .QN(\clk_gate_u_decode_u_regfile_reg_r26_q_reg_0/n2 ) );
  TLATX1 \clk_gate_u_decode_u_regfile_reg_r27_q_reg/latch  ( .G(n73546), .D(
        n17290), .QN(\clk_gate_u_decode_u_regfile_reg_r27_q_reg/n2 ) );
  TLATX1 \clk_gate_u_decode_u_regfile_reg_r27_q_reg_0/latch  ( .G(n73546), .D(
        n17291), .QN(\clk_gate_u_decode_u_regfile_reg_r27_q_reg_0/n2 ) );
  TLATX1 \clk_gate_u_decode_u_regfile_reg_r25_q_reg/latch  ( .G(n73546), .D(
        n17292), .QN(\clk_gate_u_decode_u_regfile_reg_r25_q_reg/n2 ) );
  TLATX1 \clk_gate_u_decode_u_regfile_reg_r25_q_reg_0/latch  ( .G(n73546), .D(
        n17293), .QN(\clk_gate_u_decode_u_regfile_reg_r25_q_reg_0/n2 ) );
  TLATX1 \clk_gate_u_decode_u_regfile_reg_r28_q_reg/latch  ( .G(n73546), .D(
        n17294), .QN(\clk_gate_u_decode_u_regfile_reg_r28_q_reg/n2 ) );
  TLATX1 \clk_gate_u_decode_u_regfile_reg_r28_q_reg_0/latch  ( .G(n73546), .D(
        n17295), .QN(\clk_gate_u_decode_u_regfile_reg_r28_q_reg_0/n2 ) );
  TLATX1 \clk_gate_u_decode_u_regfile_reg_r24_q_reg/latch  ( .G(n73546), .D(
        n17296), .QN(\clk_gate_u_decode_u_regfile_reg_r24_q_reg/n2 ) );
  TLATX1 \clk_gate_u_decode_u_regfile_reg_r24_q_reg_0/latch  ( .G(n73546), .D(
        n17297), .QN(\clk_gate_u_decode_u_regfile_reg_r24_q_reg_0/n2 ) );
  TLATX1 \clk_gate_u_decode_u_regfile_reg_r29_q_reg/latch  ( .G(n73546), .D(
        n17298), .QN(\clk_gate_u_decode_u_regfile_reg_r29_q_reg/n2 ) );
  TLATX1 \clk_gate_u_decode_u_regfile_reg_r29_q_reg_0/latch  ( .G(n73546), .D(
        n17299), .QN(\clk_gate_u_decode_u_regfile_reg_r29_q_reg_0/n2 ) );
  TLATX1 \clk_gate_u_decode_u_regfile_reg_r23_q_reg/latch  ( .G(n73546), .D(
        n17300), .QN(\clk_gate_u_decode_u_regfile_reg_r23_q_reg/n2 ) );
  TLATX1 \clk_gate_u_decode_u_regfile_reg_r23_q_reg_0/latch  ( .G(n73546), .D(
        n17301), .QN(\clk_gate_u_decode_u_regfile_reg_r23_q_reg_0/n2 ) );
  TLATX1 \clk_gate_u_decode_u_regfile_reg_r30_q_reg/latch  ( .G(n73546), .D(
        n17302), .QN(\clk_gate_u_decode_u_regfile_reg_r30_q_reg/n2 ) );
  TLATX1 \clk_gate_u_decode_u_regfile_reg_r30_q_reg_0/latch  ( .G(n73546), .D(
        n17303), .QN(\clk_gate_u_decode_u_regfile_reg_r30_q_reg_0/n2 ) );
  TLATX1 \clk_gate_u_decode_u_regfile_reg_r22_q_reg/latch  ( .G(n73546), .D(
        n17304), .QN(\clk_gate_u_decode_u_regfile_reg_r22_q_reg/n2 ) );
  TLATX1 \clk_gate_u_decode_u_regfile_reg_r22_q_reg_0/latch  ( .G(n73546), .D(
        n17305), .QN(\clk_gate_u_decode_u_regfile_reg_r22_q_reg_0/n2 ) );
  TLATX1 \clk_gate_u_fetch_pc_d_q_reg/latch  ( .G(n73546), .D(n17306), .QN(
        \clk_gate_u_fetch_pc_d_q_reg/n2 ) );
  TLATX1 \clk_gate_u_fetch_pc_d_q_reg_0/latch  ( .G(n73546), .D(n17307), .QN(
        \clk_gate_u_fetch_pc_d_q_reg_0/n2 ) );
  TLATX1 \clk_gate_u_fetch_branch_pc_q_reg/latch  ( .G(n73546), .D(n17308), 
        .QN(\clk_gate_u_fetch_branch_pc_q_reg/n2 ) );
  TLATX1 \clk_gate_u_fetch_branch_pc_q_reg_0/latch  ( .G(n73546), .D(n17309), 
        .QN(\clk_gate_u_fetch_branch_pc_q_reg_0/n2 ) );
  TLATX1 \clk_gate_u_fetch_fetch_pc_q_reg/latch  ( .G(n73546), .D(n17310), 
        .QN(\clk_gate_u_fetch_fetch_pc_q_reg/n2 ) );
  TLATX1 \clk_gate_u_fetch_fetch_pc_q_reg_0/latch  ( .G(n73546), .D(n17311), 
        .QN(\clk_gate_u_fetch_fetch_pc_q_reg_0/n2 ) );
  TLATX1 \clk_gate_u_fetch_skid_buffer_q_reg/latch  ( .G(n73546), .D(n17312), 
        .QN(\clk_gate_u_fetch_skid_buffer_q_reg/n2 ) );
  TLATX1 \clk_gate_u_fetch_skid_buffer_q_reg_0/latch  ( .G(n73546), .D(n17313), 
        .QN(\clk_gate_u_fetch_skid_buffer_q_reg_0/n2 ) );
  TLATX1 \clk_gate_u_fetch_skid_buffer_q_reg_1/latch  ( .G(n73546), .D(n17314), 
        .QN(\clk_gate_u_fetch_skid_buffer_q_reg_1/n2 ) );
  TLATX1 \clk_gate_u_fetch_skid_buffer_q_reg_2/latch  ( .G(n73546), .D(n17315), 
        .QN(\clk_gate_u_fetch_skid_buffer_q_reg_2/n2 ) );
  DFFRHQX1 u_muldiv_mult_result_q_reg_24_ ( .D(u_muldiv_result_r[24]), .CK(
        clk_i), .RN(n38344), .Q(u_muldiv_mult_result_q[24]) );
  DFFRHQX1 u_muldiv_mult_result_q_reg_25_ ( .D(u_muldiv_result_r[25]), .CK(
        clk_i), .RN(n38346), .Q(u_muldiv_mult_result_q[25]) );
  DFFRHQX1 u_muldiv_mult_result_q_reg_26_ ( .D(u_muldiv_result_r[26]), .CK(
        clk_i), .RN(n38344), .Q(u_muldiv_mult_result_q[26]) );
  DFFRHQX1 u_muldiv_mult_result_q_reg_27_ ( .D(u_muldiv_result_r[27]), .CK(
        clk_i), .RN(n38345), .Q(u_muldiv_mult_result_q[27]) );
  DFFRHQX1 u_decode_u_regfile_reg_r16_q_reg_20_ ( .D(u_decode_u_regfile_N675), 
        .CK(n37815), .RN(n44247), .Q(n2408) );
  DFFRHQX1 u_decode_u_regfile_reg_r19_q_reg_20_ ( .D(u_decode_u_regfile_N786), 
        .CK(n37812), .RN(n44247), .Q(n2411) );
  DFFRHQX1 u_exec_result_q_reg_31_ ( .D(u_exec_alu_p_w[31]), .CK(clk_i), .RN(
        n38340), .Q(writeback_exec_value_w[31]) );
  DFFRHQX1 u_decode_opcode_instr_q_reg_48_ ( .D(u_decode_N784), .CK(n37885), 
        .RN(n44207), .Q(opcode_instr_w_48) );
  DFFRHQX1 u_decode_opcode_instr_q_reg_49_ ( .D(u_decode_N785), .CK(n37885), 
        .RN(n44207), .Q(n42614) );
  DFFRHQX1 u_exec_result_q_reg_30_ ( .D(u_exec_alu_p_w[30]), .CK(clk_i), .RN(
        n44180), .Q(n43235) );
  DFFRHQX1 u_exec_result_q_reg_27_ ( .D(u_exec_alu_p_w[27]), .CK(clk_i), .RN(
        n44189), .Q(n43216) );
  DFFRHQX1 u_decode_u_regfile_reg_r21_q_reg_0_ ( .D(u_decode_u_regfile_N840), 
        .CK(n37838), .RN(n38320), .Q(n1969) );
  DFFRHQX1 u_decode_u_regfile_reg_r21_q_reg_1_ ( .D(u_decode_u_regfile_N841), 
        .CK(n37838), .RN(n38336), .Q(n2001) );
  DFFRHQX1 u_decode_u_regfile_reg_r18_q_reg_1_ ( .D(u_decode_u_regfile_N730), 
        .CK(n37844), .RN(n38335), .Q(n1998) );
  DFFRHQX1 u_decode_u_regfile_reg_r8_q_reg_0_ ( .D(u_decode_u_regfile_N359), 
        .CK(n37839), .RN(n44119), .Q(n42613) );
  DFFRHQX1 u_decode_u_regfile_reg_r24_q_reg_0_ ( .D(u_decode_u_regfile_N951), 
        .CK(n37878), .RN(n44132), .Q(n42612) );
  DFFRHQX1 u_decode_u_regfile_reg_r5_q_reg_0_ ( .D(u_decode_u_regfile_N248), 
        .CK(n37840), .RN(n44130), .Q(n1953) );
  DFFRX1 u_decode_u_regfile_reg_r30_q_reg_21_ ( .D(u_decode_u_regfile_N1194), 
        .CK(n37832), .RN(n44247), .Q(n2556), .QN(n42820) );
  DFFRX1 u_decode_u_regfile_reg_r7_q_reg_21_ ( .D(u_decode_u_regfile_N343), 
        .CK(n37824), .RN(n44247), .QN(n46696) );
  DFFRX1 u_decode_u_regfile_reg_r7_q_reg_23_ ( .D(u_decode_u_regfile_N345), 
        .CK(n37824), .RN(n44248), .QN(n46626) );
  DFFRX1 u_decode_u_regfile_reg_r14_q_reg_1_ ( .D(u_decode_u_regfile_N582), 
        .CK(n37848), .RN(n73547), .Q(n1994), .QN(n48163) );
  DFFRX1 u_decode_u_regfile_reg_r3_q_reg_1_ ( .D(u_decode_u_regfile_N175), 
        .CK(n37857), .RN(n38336), .QN(n48211) );
  DFFRX1 u_decode_u_regfile_reg_r19_q_reg_1_ ( .D(u_decode_u_regfile_N767), 
        .CK(n37843), .RN(n38335), .QN(n48180) );
  DFFRX1 u_exec_rd_x_q_reg_1_ ( .D(u_exec_N239), .CK(clk_i), .RN(n38321), .Q(
        writeback_exec_idx_w[1]), .QN(n50720) );
  DFFRX1 u_exec_rd_x_q_reg_0_ ( .D(u_exec_N238), .CK(clk_i), .RN(n38322), .Q(
        writeback_exec_idx_w[0]), .QN(n50824) );
  DFFRHQX1 u_muldiv_mult_result_q_reg_28_ ( .D(u_muldiv_result_r[28]), .CK(
        clk_i), .RN(n38347), .Q(u_muldiv_mult_result_q[28]) );
  DFFRHQX1 u_muldiv_mult_result_q_reg_29_ ( .D(u_muldiv_result_r[29]), .CK(
        clk_i), .RN(n38345), .Q(u_muldiv_mult_result_q[29]) );
  DFFRX1 u_decode_inst_q_reg_18_ ( .D(u_decode_N340), .CK(n37870), .RN(n73547), 
        .Q(opcode_opcode_w[18]), .QN(n42666) );
  DFFRX1 u_decode_inst_q_reg_15_ ( .D(u_decode_N337), .CK(n37870), .RN(n44252), 
        .Q(opcode_opcode_w[15]), .QN(n42732) );
  DFFRX1 u_decode_inst_q_reg_22_ ( .D(n8511), .CK(clk_i), .RN(n38350), .Q(
        opcode_opcode_w[22]), .QN(n42814) );
  DFFRX1 u_decode_inst_q_reg_21_ ( .D(n73540), .CK(n37870), .RN(n38349), .Q(
        opcode_opcode_w[21]), .QN(n42763) );
  DFFRX1 u_decode_inst_q_reg_23_ ( .D(n8512), .CK(clk_i), .RN(n38351), .Q(
        opcode_opcode_w[23]), .QN(n42761) );
  DFFRX1 u_decode_inst_q_reg_20_ ( .D(u_decode_N342), .CK(n37870), .RN(n38351), 
        .Q(opcode_opcode_w[20]), .QN(n42740) );
  DFFRX1 u_decode_inst_q_reg_24_ ( .D(n8513), .CK(clk_i), .RN(n73547), .Q(
        opcode_opcode_w[24]), .QN(n42750) );
  DFFRHQX1 u_csr_csr_stval_q_reg_12_ ( .D(u_csr_csr_stval_r[12]), .CK(clk_i), 
        .RN(n38332), .Q(u_csr_csr_stval_q[12]) );
  DFFRHQX1 u_csr_csr_stval_q_reg_11_ ( .D(u_csr_csr_stval_r[11]), .CK(clk_i), 
        .RN(n38331), .Q(u_csr_csr_stval_q[11]) );
  DFFRHQX1 u_csr_csr_stval_q_reg_10_ ( .D(u_csr_csr_stval_r[10]), .CK(clk_i), 
        .RN(n38330), .Q(u_csr_csr_stval_q[10]) );
  DFFRHQX1 u_csr_csr_sscratch_q_reg_3_ ( .D(u_csr_csr_sscratch_r[3]), .CK(
        clk_i), .RN(n38355), .Q(u_csr_csr_sscratch_q[3]) );
  DFFRHQX1 u_csr_csr_sscratch_q_reg_1_ ( .D(u_csr_csr_sscratch_r[1]), .CK(
        clk_i), .RN(n38354), .Q(u_csr_csr_sscratch_q[1]) );
  DFFRHQX1 u_csr_csr_sscratch_q_reg_4_ ( .D(u_csr_csr_sscratch_r[4]), .CK(
        clk_i), .RN(n38357), .Q(u_csr_csr_sscratch_q[4]) );
  DFFRHQX1 u_csr_csr_sscratch_q_reg_0_ ( .D(u_csr_csr_sscratch_r[0]), .CK(
        clk_i), .RN(n38356), .Q(u_csr_csr_sscratch_q[0]) );
  DFFRHQX1 u_csr_csr_sscratch_q_reg_2_ ( .D(u_csr_csr_sscratch_r[2]), .CK(
        clk_i), .RN(n38355), .Q(u_csr_csr_sscratch_q[2]) );
  DFFRHQX1 u_muldiv_divisor_q_reg_59_ ( .D(u_muldiv_N324), .CK(net1898), .RN(
        n38333), .Q(u_muldiv_divisor_q[59]) );
  DFFRHQX1 u_csr_csr_mscratch_q_reg_11_ ( .D(u_csr_csr_mscratch_r[11]), .CK(
        clk_i), .RN(n38328), .Q(u_csr_csr_mscratch_q[11]) );
  DFFRHQX1 u_csr_csr_mscratch_q_reg_8_ ( .D(u_csr_csr_mscratch_r[8]), .CK(
        clk_i), .RN(n38327), .Q(u_csr_csr_mscratch_q[8]) );
  DFFRHQX1 u_csr_csr_mscratch_q_reg_7_ ( .D(u_csr_csr_mscratch_r[7]), .CK(
        clk_i), .RN(n38326), .Q(u_csr_csr_mscratch_q[7]) );
  DFFRHQX1 u_csr_csr_mscratch_q_reg_5_ ( .D(u_csr_csr_mscratch_r[5]), .CK(
        clk_i), .RN(n38325), .Q(u_csr_csr_mscratch_q[5]) );
  DFFRHQX1 u_csr_csr_mscratch_q_reg_31_ ( .D(u_csr_csr_mscratch_r[31]), .CK(
        clk_i), .RN(n38328), .Q(u_csr_csr_mscratch_q[31]) );
  DFFRHQX1 u_csr_csr_mscratch_q_reg_30_ ( .D(u_csr_csr_mscratch_r[30]), .CK(
        clk_i), .RN(n38327), .Q(u_csr_csr_mscratch_q[30]) );
  DFFRHQX1 u_csr_csr_mscratch_q_reg_29_ ( .D(u_csr_csr_mscratch_r[29]), .CK(
        clk_i), .RN(n38326), .Q(u_csr_csr_mscratch_q[29]) );
  DFFRHQX1 u_csr_csr_mscratch_q_reg_28_ ( .D(u_csr_csr_mscratch_r[28]), .CK(
        clk_i), .RN(n38325), .Q(u_csr_csr_mscratch_q[28]) );
  DFFRHQX1 u_csr_csr_mscratch_q_reg_27_ ( .D(u_csr_csr_mscratch_r[27]), .CK(
        clk_i), .RN(n38328), .Q(u_csr_csr_mscratch_q[27]) );
  DFFRHQX1 u_csr_csr_mscratch_q_reg_26_ ( .D(u_csr_csr_mscratch_r[26]), .CK(
        clk_i), .RN(n38327), .Q(u_csr_csr_mscratch_q[26]) );
  DFFRHQX1 u_csr_csr_mscratch_q_reg_25_ ( .D(u_csr_csr_mscratch_r[25]), .CK(
        clk_i), .RN(n38326), .Q(u_csr_csr_mscratch_q[25]) );
  DFFRHQX1 u_csr_csr_mscratch_q_reg_24_ ( .D(u_csr_csr_mscratch_r[24]), .CK(
        clk_i), .RN(n38325), .Q(u_csr_csr_mscratch_q[24]) );
  DFFRHQX1 u_csr_csr_mscratch_q_reg_23_ ( .D(u_csr_csr_mscratch_r[23]), .CK(
        clk_i), .RN(n38328), .Q(u_csr_csr_mscratch_q[23]) );
  DFFRHQX1 u_csr_csr_mscratch_q_reg_22_ ( .D(u_csr_csr_mscratch_r[22]), .CK(
        clk_i), .RN(n38327), .Q(u_csr_csr_mscratch_q[22]) );
  DFFRHQX1 u_csr_csr_mscratch_q_reg_21_ ( .D(u_csr_csr_mscratch_r[21]), .CK(
        clk_i), .RN(n38326), .Q(u_csr_csr_mscratch_q[21]) );
  DFFRHQX1 u_csr_csr_mscratch_q_reg_20_ ( .D(u_csr_csr_mscratch_r[20]), .CK(
        clk_i), .RN(n38325), .Q(u_csr_csr_mscratch_q[20]) );
  DFFRHQX1 u_csr_csr_mscratch_q_reg_19_ ( .D(u_csr_csr_mscratch_r[19]), .CK(
        clk_i), .RN(n38328), .Q(u_csr_csr_mscratch_q[19]) );
  DFFRHQX1 u_csr_csr_mscratch_q_reg_18_ ( .D(u_csr_csr_mscratch_r[18]), .CK(
        clk_i), .RN(n38327), .Q(u_csr_csr_mscratch_q[18]) );
  DFFRHQX1 u_csr_csr_mscratch_q_reg_17_ ( .D(u_csr_csr_mscratch_r[17]), .CK(
        clk_i), .RN(n38326), .Q(u_csr_csr_mscratch_q[17]) );
  DFFRHQX1 u_csr_csr_mscratch_q_reg_16_ ( .D(u_csr_csr_mscratch_r[16]), .CK(
        clk_i), .RN(n38325), .Q(u_csr_csr_mscratch_q[16]) );
  DFFRHQX1 u_csr_csr_mscratch_q_reg_13_ ( .D(u_csr_csr_mscratch_r[13]), .CK(
        clk_i), .RN(n38328), .Q(u_csr_csr_mscratch_q[13]) );
  DFFRHQX1 u_csr_csr_mscratch_q_reg_12_ ( .D(u_csr_csr_mscratch_r[12]), .CK(
        clk_i), .RN(n38327), .Q(u_csr_csr_mscratch_q[12]) );
  DFFRHQX1 u_csr_csr_mscratch_q_reg_15_ ( .D(u_csr_csr_mscratch_r[15]), .CK(
        clk_i), .RN(n38326), .Q(u_csr_csr_mscratch_q[15]) );
  DFFRHQX1 u_csr_csr_mscratch_q_reg_14_ ( .D(u_csr_csr_mscratch_r[14]), .CK(
        clk_i), .RN(n38325), .Q(u_csr_csr_mscratch_q[14]) );
  DFFRHQX1 u_csr_csr_stvec_q_reg_11_ ( .D(u_csr_csr_stvec_r[11]), .CK(clk_i), 
        .RN(n44249), .Q(u_csr_csr_stvec_q[11]) );
  DFFRHQX1 u_csr_csr_stvec_q_reg_10_ ( .D(u_csr_csr_stvec_r[10]), .CK(clk_i), 
        .RN(n38354), .Q(u_csr_csr_stvec_q[10]) );
  DFFRHQX1 u_csr_csr_stvec_q_reg_12_ ( .D(u_csr_csr_stvec_r[12]), .CK(clk_i), 
        .RN(n38357), .Q(u_csr_csr_stvec_q[12]) );
  DFFRHQX1 u_csr_csr_sscratch_q_reg_11_ ( .D(u_csr_csr_sscratch_r[11]), .CK(
        clk_i), .RN(n44249), .Q(u_csr_csr_sscratch_q[11]) );
  DFFRHQX1 u_csr_csr_sscratch_q_reg_5_ ( .D(u_csr_csr_sscratch_r[5]), .CK(
        clk_i), .RN(n38356), .Q(u_csr_csr_sscratch_q[5]) );
  DFFRHQX1 u_csr_csr_sscratch_q_reg_31_ ( .D(u_csr_csr_sscratch_r[31]), .CK(
        clk_i), .RN(n38355), .Q(u_csr_csr_sscratch_q[31]) );
  DFFRHQX1 u_csr_csr_sscratch_q_reg_30_ ( .D(u_csr_csr_sscratch_r[30]), .CK(
        clk_i), .RN(n38354), .Q(u_csr_csr_sscratch_q[30]) );
  DFFRHQX1 u_csr_csr_sscratch_q_reg_29_ ( .D(u_csr_csr_sscratch_r[29]), .CK(
        clk_i), .RN(n38357), .Q(u_csr_csr_sscratch_q[29]) );
  DFFRHQX1 u_csr_csr_sscratch_q_reg_28_ ( .D(u_csr_csr_sscratch_r[28]), .CK(
        clk_i), .RN(n38356), .Q(u_csr_csr_sscratch_q[28]) );
  DFFRHQX1 u_csr_csr_sscratch_q_reg_27_ ( .D(u_csr_csr_sscratch_r[27]), .CK(
        clk_i), .RN(n38355), .Q(u_csr_csr_sscratch_q[27]) );
  DFFRHQX1 u_csr_csr_sscratch_q_reg_26_ ( .D(u_csr_csr_sscratch_r[26]), .CK(
        clk_i), .RN(n38354), .Q(u_csr_csr_sscratch_q[26]) );
  DFFRHQX1 u_csr_csr_sscratch_q_reg_25_ ( .D(u_csr_csr_sscratch_r[25]), .CK(
        clk_i), .RN(n38357), .Q(u_csr_csr_sscratch_q[25]) );
  DFFRHQX1 u_csr_csr_sscratch_q_reg_24_ ( .D(u_csr_csr_sscratch_r[24]), .CK(
        clk_i), .RN(n38356), .Q(u_csr_csr_sscratch_q[24]) );
  DFFRHQX1 u_csr_csr_sscratch_q_reg_23_ ( .D(u_csr_csr_sscratch_r[23]), .CK(
        clk_i), .RN(n38355), .Q(u_csr_csr_sscratch_q[23]) );
  DFFRHQX1 u_csr_csr_sscratch_q_reg_22_ ( .D(u_csr_csr_sscratch_r[22]), .CK(
        clk_i), .RN(n38354), .Q(u_csr_csr_sscratch_q[22]) );
  DFFRHQX1 u_csr_csr_sscratch_q_reg_10_ ( .D(u_csr_csr_sscratch_r[10]), .CK(
        clk_i), .RN(n38357), .Q(u_csr_csr_sscratch_q[10]) );
  DFFRHQX1 u_csr_csr_sscratch_q_reg_6_ ( .D(u_csr_csr_sscratch_r[6]), .CK(
        clk_i), .RN(n38356), .Q(u_csr_csr_sscratch_q[6]) );
  DFFRHQX1 u_csr_csr_sscratch_q_reg_21_ ( .D(u_csr_csr_sscratch_r[21]), .CK(
        clk_i), .RN(n38355), .Q(u_csr_csr_sscratch_q[21]) );
  DFFRHQX1 u_csr_csr_sscratch_q_reg_20_ ( .D(u_csr_csr_sscratch_r[20]), .CK(
        clk_i), .RN(n38354), .Q(u_csr_csr_sscratch_q[20]) );
  DFFRHQX1 u_csr_csr_sscratch_q_reg_19_ ( .D(u_csr_csr_sscratch_r[19]), .CK(
        clk_i), .RN(n38357), .Q(u_csr_csr_sscratch_q[19]) );
  DFFRHQX1 u_csr_csr_sscratch_q_reg_18_ ( .D(u_csr_csr_sscratch_r[18]), .CK(
        clk_i), .RN(n38356), .Q(u_csr_csr_sscratch_q[18]) );
  DFFRHQX1 u_csr_csr_sscratch_q_reg_17_ ( .D(u_csr_csr_sscratch_r[17]), .CK(
        clk_i), .RN(n38355), .Q(u_csr_csr_sscratch_q[17]) );
  DFFRHQX1 u_csr_csr_sscratch_q_reg_16_ ( .D(u_csr_csr_sscratch_r[16]), .CK(
        clk_i), .RN(n38354), .Q(u_csr_csr_sscratch_q[16]) );
  DFFRHQX1 u_csr_csr_sscratch_q_reg_13_ ( .D(u_csr_csr_sscratch_r[13]), .CK(
        clk_i), .RN(n38357), .Q(u_csr_csr_sscratch_q[13]) );
  DFFRHQX1 u_csr_csr_sscratch_q_reg_12_ ( .D(u_csr_csr_sscratch_r[12]), .CK(
        clk_i), .RN(n38356), .Q(u_csr_csr_sscratch_q[12]) );
  DFFRHQX1 u_csr_csr_sscratch_q_reg_15_ ( .D(u_csr_csr_sscratch_r[15]), .CK(
        clk_i), .RN(n38355), .Q(u_csr_csr_sscratch_q[15]) );
  DFFRHQX1 u_csr_csr_sscratch_q_reg_14_ ( .D(u_csr_csr_sscratch_r[14]), .CK(
        clk_i), .RN(n38354), .Q(u_csr_csr_sscratch_q[14]) );
  DFFRHQX1 u_csr_csr_stval_q_reg_9_ ( .D(u_csr_csr_stval_r[9]), .CK(clk_i), 
        .RN(n38332), .Q(u_csr_csr_stval_q[9]) );
  DFFRHQX1 u_csr_csr_stval_q_reg_8_ ( .D(u_csr_csr_stval_r[8]), .CK(clk_i), 
        .RN(n38331), .Q(u_csr_csr_stval_q[8]) );
  DFFRHQX1 u_csr_csr_stval_q_reg_7_ ( .D(u_csr_csr_stval_r[7]), .CK(clk_i), 
        .RN(n38330), .Q(u_csr_csr_stval_q[7]) );
  DFFRHQX1 u_csr_csr_stval_q_reg_31_ ( .D(u_csr_csr_stval_r[31]), .CK(clk_i), 
        .RN(n44249), .Q(u_csr_csr_stval_q[31]) );
  DFFRHQX1 u_csr_csr_stval_q_reg_6_ ( .D(u_csr_csr_stval_r[6]), .CK(clk_i), 
        .RN(n38333), .Q(u_csr_csr_stval_q[6]) );
  DFFRHQX1 u_csr_csr_stval_q_reg_5_ ( .D(u_csr_csr_stval_r[5]), .CK(clk_i), 
        .RN(n38332), .Q(u_csr_csr_stval_q[5]) );
  DFFRHQX1 u_csr_csr_stval_q_reg_30_ ( .D(u_csr_csr_stval_r[30]), .CK(clk_i), 
        .RN(n44249), .Q(u_csr_csr_stval_q[30]) );
  DFFRHQX1 u_csr_csr_stval_q_reg_29_ ( .D(u_csr_csr_stval_r[29]), .CK(clk_i), 
        .RN(n44249), .Q(u_csr_csr_stval_q[29]) );
  DFFRHQX1 u_csr_csr_stval_q_reg_28_ ( .D(u_csr_csr_stval_r[28]), .CK(clk_i), 
        .RN(n38331), .Q(u_csr_csr_stval_q[28]) );
  DFFRHQX1 u_csr_csr_stval_q_reg_27_ ( .D(u_csr_csr_stval_r[27]), .CK(clk_i), 
        .RN(n38330), .Q(u_csr_csr_stval_q[27]) );
  DFFRHQX1 u_csr_csr_stval_q_reg_26_ ( .D(u_csr_csr_stval_r[26]), .CK(clk_i), 
        .RN(n38333), .Q(u_csr_csr_stval_q[26]) );
  DFFRHQX1 u_csr_csr_stval_q_reg_25_ ( .D(u_csr_csr_stval_r[25]), .CK(clk_i), 
        .RN(n38332), .Q(u_csr_csr_stval_q[25]) );
  DFFRHQX1 u_csr_csr_stval_q_reg_24_ ( .D(u_csr_csr_stval_r[24]), .CK(clk_i), 
        .RN(n38331), .Q(u_csr_csr_stval_q[24]) );
  DFFRHQX1 u_csr_csr_stval_q_reg_23_ ( .D(u_csr_csr_stval_r[23]), .CK(clk_i), 
        .RN(n38330), .Q(u_csr_csr_stval_q[23]) );
  DFFRHQX1 u_csr_csr_stval_q_reg_22_ ( .D(u_csr_csr_stval_r[22]), .CK(clk_i), 
        .RN(n38333), .Q(u_csr_csr_stval_q[22]) );
  DFFRHQX1 u_csr_csr_stval_q_reg_21_ ( .D(u_csr_csr_stval_r[21]), .CK(clk_i), 
        .RN(n38332), .Q(u_csr_csr_stval_q[21]) );
  DFFRHQX1 u_csr_csr_stval_q_reg_20_ ( .D(u_csr_csr_stval_r[20]), .CK(clk_i), 
        .RN(n38331), .Q(u_csr_csr_stval_q[20]) );
  DFFRHQX1 u_csr_csr_stval_q_reg_19_ ( .D(u_csr_csr_stval_r[19]), .CK(clk_i), 
        .RN(n38330), .Q(u_csr_csr_stval_q[19]) );
  DFFRHQX1 u_csr_csr_stval_q_reg_18_ ( .D(u_csr_csr_stval_r[18]), .CK(clk_i), 
        .RN(n38333), .Q(u_csr_csr_stval_q[18]) );
  DFFRHQX1 u_csr_csr_stval_q_reg_17_ ( .D(u_csr_csr_stval_r[17]), .CK(clk_i), 
        .RN(n38332), .Q(u_csr_csr_stval_q[17]) );
  DFFRHQX1 u_csr_csr_stval_q_reg_16_ ( .D(u_csr_csr_stval_r[16]), .CK(clk_i), 
        .RN(n38331), .Q(u_csr_csr_stval_q[16]) );
  DFFRHQX1 u_csr_csr_stval_q_reg_15_ ( .D(u_csr_csr_stval_r[15]), .CK(clk_i), 
        .RN(n44249), .Q(u_csr_csr_stval_q[15]) );
  DFFRHQX1 u_csr_csr_stval_q_reg_14_ ( .D(u_csr_csr_stval_r[14]), .CK(clk_i), 
        .RN(n44249), .Q(u_csr_csr_stval_q[14]) );
  DFFRHQX1 u_csr_csr_stval_q_reg_13_ ( .D(u_csr_csr_stval_r[13]), .CK(clk_i), 
        .RN(n38330), .Q(u_csr_csr_stval_q[13]) );
  DFFRHQX1 u_csr_csr_stvec_q_reg_8_ ( .D(u_csr_csr_stvec_r[8]), .CK(clk_i), 
        .RN(n38357), .Q(u_csr_csr_stvec_q[8]) );
  DFFRHQX1 u_csr_csr_stvec_q_reg_7_ ( .D(u_csr_csr_stvec_r[7]), .CK(clk_i), 
        .RN(n38356), .Q(u_csr_csr_stvec_q[7]) );
  DFFRHQX1 u_csr_csr_stvec_q_reg_5_ ( .D(u_csr_csr_stvec_r[5]), .CK(clk_i), 
        .RN(n38355), .Q(u_csr_csr_stvec_q[5]) );
  DFFRHQX1 u_csr_csr_stvec_q_reg_31_ ( .D(u_csr_csr_stvec_r[31]), .CK(clk_i), 
        .RN(n38354), .Q(u_csr_csr_stvec_q[31]) );
  DFFRHQX1 u_csr_csr_stvec_q_reg_30_ ( .D(u_csr_csr_stvec_r[30]), .CK(clk_i), 
        .RN(n38357), .Q(u_csr_csr_stvec_q[30]) );
  DFFRHQX1 u_csr_csr_stvec_q_reg_29_ ( .D(u_csr_csr_stvec_r[29]), .CK(clk_i), 
        .RN(n38356), .Q(u_csr_csr_stvec_q[29]) );
  DFFRHQX1 u_csr_csr_stvec_q_reg_28_ ( .D(u_csr_csr_stvec_r[28]), .CK(clk_i), 
        .RN(n38355), .Q(u_csr_csr_stvec_q[28]) );
  DFFRHQX1 u_csr_csr_stvec_q_reg_27_ ( .D(u_csr_csr_stvec_r[27]), .CK(clk_i), 
        .RN(n38354), .Q(u_csr_csr_stvec_q[27]) );
  DFFRHQX1 u_csr_csr_stvec_q_reg_26_ ( .D(u_csr_csr_stvec_r[26]), .CK(clk_i), 
        .RN(n38357), .Q(u_csr_csr_stvec_q[26]) );
  DFFRHQX1 u_csr_csr_stvec_q_reg_25_ ( .D(u_csr_csr_stvec_r[25]), .CK(clk_i), 
        .RN(n38356), .Q(u_csr_csr_stvec_q[25]) );
  DFFRHQX1 u_csr_csr_stvec_q_reg_24_ ( .D(u_csr_csr_stvec_r[24]), .CK(clk_i), 
        .RN(n38355), .Q(u_csr_csr_stvec_q[24]) );
  DFFRHQX1 u_csr_csr_stvec_q_reg_23_ ( .D(u_csr_csr_stvec_r[23]), .CK(clk_i), 
        .RN(n38354), .Q(u_csr_csr_stvec_q[23]) );
  DFFRHQX1 u_csr_csr_stvec_q_reg_22_ ( .D(u_csr_csr_stvec_r[22]), .CK(clk_i), 
        .RN(n38357), .Q(u_csr_csr_stvec_q[22]) );
  DFFRHQX1 u_csr_csr_stvec_q_reg_9_ ( .D(u_csr_csr_stvec_r[9]), .CK(clk_i), 
        .RN(n38356), .Q(u_csr_csr_stvec_q[9]) );
  DFFRHQX1 u_csr_csr_stvec_q_reg_6_ ( .D(u_csr_csr_stvec_r[6]), .CK(clk_i), 
        .RN(n38355), .Q(u_csr_csr_stvec_q[6]) );
  DFFRHQX1 u_csr_csr_stvec_q_reg_21_ ( .D(u_csr_csr_stvec_r[21]), .CK(clk_i), 
        .RN(n38354), .Q(u_csr_csr_stvec_q[21]) );
  DFFRHQX1 u_csr_csr_stvec_q_reg_20_ ( .D(u_csr_csr_stvec_r[20]), .CK(clk_i), 
        .RN(n38357), .Q(u_csr_csr_stvec_q[20]) );
  DFFRHQX1 u_csr_csr_stvec_q_reg_19_ ( .D(u_csr_csr_stvec_r[19]), .CK(clk_i), 
        .RN(n38356), .Q(u_csr_csr_stvec_q[19]) );
  DFFRHQX1 u_csr_csr_stvec_q_reg_18_ ( .D(u_csr_csr_stvec_r[18]), .CK(clk_i), 
        .RN(n38355), .Q(u_csr_csr_stvec_q[18]) );
  DFFRHQX1 u_csr_csr_stvec_q_reg_17_ ( .D(u_csr_csr_stvec_r[17]), .CK(clk_i), 
        .RN(n38354), .Q(u_csr_csr_stvec_q[17]) );
  DFFRHQX1 u_csr_csr_stvec_q_reg_16_ ( .D(u_csr_csr_stvec_r[16]), .CK(clk_i), 
        .RN(n38357), .Q(u_csr_csr_stvec_q[16]) );
  DFFRHQX1 u_csr_csr_stvec_q_reg_13_ ( .D(u_csr_csr_stvec_r[13]), .CK(clk_i), 
        .RN(n38356), .Q(u_csr_csr_stvec_q[13]) );
  DFFRHQX1 u_csr_csr_stvec_q_reg_15_ ( .D(u_csr_csr_stvec_r[15]), .CK(clk_i), 
        .RN(n38355), .Q(u_csr_csr_stvec_q[15]) );
  DFFRHQX1 u_csr_csr_stvec_q_reg_14_ ( .D(u_csr_csr_stvec_r[14]), .CK(clk_i), 
        .RN(n38354), .Q(u_csr_csr_stvec_q[14]) );
  DFFRHQX1 u_muldiv_divisor_q_reg_60_ ( .D(u_muldiv_N325), .CK(net1898), .RN(
        n38333), .Q(u_muldiv_divisor_q[60]) );
  DFFRHQX1 u_muldiv_dividend_q_reg_19_ ( .D(u_muldiv_N251), .CK(net1913), .RN(
        n38332), .Q(u_muldiv_dividend_q[19]) );
  DFFRHQX1 u_muldiv_divisor_q_reg_61_ ( .D(u_muldiv_N326), .CK(net1898), .RN(
        n38331), .Q(u_muldiv_divisor_q[61]) );
  DFFRHQX1 u_muldiv_divisor_q_reg_62_ ( .D(u_muldiv_N327), .CK(net1898), .RN(
        n38346), .Q(u_muldiv_divisor_q[62]) );
  DFFRHQX1 u_muldiv_dividend_q_reg_20_ ( .D(u_muldiv_N252), .CK(net1913), .RN(
        n38330), .Q(u_muldiv_dividend_q[20]) );
  DFFRHQX1 u_muldiv_invert_res_q_reg ( .D(n8520), .CK(clk_i), .RN(n44249), .Q(
        u_muldiv_invert_res_q) );
  DFFRHQX1 u_muldiv_dividend_q_reg_21_ ( .D(u_muldiv_N253), .CK(net1913), .RN(
        n38333), .Q(u_muldiv_dividend_q[21]) );
  DFFRHQX1 u_muldiv_dividend_q_reg_22_ ( .D(u_muldiv_N254), .CK(net1913), .RN(
        n38332), .Q(u_muldiv_dividend_q[22]) );
  DFFRHQX1 u_muldiv_dividend_q_reg_23_ ( .D(u_muldiv_N255), .CK(net1913), .RN(
        n38331), .Q(u_muldiv_dividend_q[23]) );
  DFFRHQX1 u_muldiv_dividend_q_reg_24_ ( .D(u_muldiv_N256), .CK(net1913), .RN(
        n38330), .Q(u_muldiv_dividend_q[24]) );
  DFFRHQX1 u_muldiv_dividend_q_reg_25_ ( .D(u_muldiv_N257), .CK(net1913), .RN(
        n38333), .Q(u_muldiv_dividend_q[25]) );
  DFFRHQX1 u_muldiv_dividend_q_reg_26_ ( .D(u_muldiv_N258), .CK(net1913), .RN(
        n38332), .Q(u_muldiv_dividend_q[26]) );
  DFFRHQX1 u_muldiv_dividend_q_reg_27_ ( .D(u_muldiv_N259), .CK(net1913), .RN(
        n38331), .Q(u_muldiv_dividend_q[27]) );
  DFFRHQX1 u_muldiv_dividend_q_reg_28_ ( .D(u_muldiv_N260), .CK(net1913), .RN(
        n44249), .Q(u_muldiv_dividend_q[28]) );
  DFFRHQX1 u_muldiv_dividend_q_reg_29_ ( .D(u_muldiv_N261), .CK(net1913), .RN(
        n38330), .Q(u_muldiv_dividend_q[29]) );
  DFFRHQX1 u_muldiv_dividend_q_reg_30_ ( .D(u_muldiv_N262), .CK(net1913), .RN(
        n44249), .Q(u_muldiv_dividend_q[30]) );
  DFFRHQX1 u_muldiv_dividend_q_reg_31_ ( .D(u_muldiv_N263), .CK(net1913), .RN(
        n44249), .Q(u_muldiv_dividend_q[31]) );
  DFFRX1 u_csr_branch_q_reg ( .D(u_csr_N3697), .CK(clk_i), .RN(n73547), .Q(
        n42596), .QN(n8696) );
  DFFRX1 u_muldiv_mult_result_q_reg_0_ ( .D(u_muldiv_result_r[0]), .CK(clk_i), 
        .RN(n38326), .Q(u_muldiv_mult_result_q[0]) );
  DFFRX1 u_muldiv_mult_result_q_reg_1_ ( .D(u_muldiv_result_r[1]), .CK(clk_i), 
        .RN(n38344), .Q(u_muldiv_mult_result_q[1]) );
  DFFRX1 u_muldiv_mult_result_q_reg_3_ ( .D(u_muldiv_result_r[3]), .CK(clk_i), 
        .RN(n38347), .Q(u_muldiv_mult_result_q[3]) );
  DFFRX1 u_muldiv_mult_result_q_reg_4_ ( .D(u_muldiv_result_r[4]), .CK(clk_i), 
        .RN(n38346), .Q(u_muldiv_mult_result_q[4]) );
  DFFRX1 u_fetch_active_q_reg ( .D(n8443), .CK(clk_i), .RN(n38356), .Q(
        u_fetch_active_q), .QN(n50044) );
  DFFRX1 u_decode_opcode_instr_q_reg_39_ ( .D(u_decode_N775), .CK(n37807), 
        .RN(n38350), .Q(opcode_instr_w_39), .QN(n58249) );
  DFFRX1 u_decode_opcode_instr_q_reg_38_ ( .D(u_decode_N774), .CK(n37807), 
        .RN(n38349), .Q(opcode_instr_w_38), .QN(n51407) );
  DFFRX1 u_muldiv_mult_result_q_reg_5_ ( .D(u_muldiv_result_r[5]), .CK(clk_i), 
        .RN(n38345), .Q(u_muldiv_mult_result_q[5]) );
  DFFRX1 u_decode_opcode_instr_q_reg_12_ ( .D(u_decode_N748), .CK(n37806), 
        .RN(n38321), .Q(opcode_instr_w[12]) );
  DFFRX1 u_decode_inst_q_reg_12_ ( .D(u_decode_N334), .CK(n37870), .RN(n38360), 
        .Q(opcode_opcode_w[12]), .QN(n56860) );
  DFFRX1 u_decode_inst_q_reg_10_ ( .D(u_decode_N332), .CK(n37870), .RN(n38352), 
        .Q(opcode_opcode_w[10]), .QN(n54447) );
  DFFRX1 u_decode_inst_q_reg_9_ ( .D(u_decode_N331), .CK(n37870), .RN(n38351), 
        .Q(opcode_opcode_w[9]), .QN(n57436) );
  DFFRX1 u_decode_inst_q_reg_7_ ( .D(u_decode_N329), .CK(n37870), .RN(n38350), 
        .Q(opcode_opcode_w[7]), .QN(n50700) );
  DFFRX1 u_decode_inst_q_reg_11_ ( .D(u_decode_N333), .CK(n37870), .RN(n38349), 
        .Q(opcode_opcode_w[11]), .QN(n54586) );
  DFFRX1 u_decode_inst_q_reg_8_ ( .D(u_decode_N330), .CK(n37870), .RN(n38352), 
        .Q(opcode_opcode_w[8]), .QN(n57429) );
  DFFRX1 u_decode_opcode_instr_q_reg_56_ ( .D(u_decode_N792), .CK(n37885), 
        .RN(n38338), .Q(opcode_instr_w_56) );
  DFFRX1 u_decode_valid_q_reg ( .D(n36342), .CK(n37870), .RN(n44252), .Q(
        u_decode_valid_q), .QN(n54383) );
  DFFRX1 u_muldiv_mult_result_q_reg_6_ ( .D(u_muldiv_result_r[6]), .CK(clk_i), 
        .RN(n38344), .Q(u_muldiv_mult_result_q[6]) );
  DFFRX1 u_decode_ifence_q_reg ( .D(u_decode_N180), .CK(clk_i), .RN(n38325), 
        .Q(mem_i_flush_o) );
  DFFRX1 u_fetch_pc_d_q_reg_31_ ( .D(\mmu_ifetch_pc_w[31] ), .CK(n37805), .RN(
        n38340), .QN(n56570) );
  DFFRX1 u_fetch_pc_d_q_reg_12_ ( .D(n21), .CK(n37804), .RN(n38359), .QN(
        n55090) );
  DFFRX1 u_fetch_pc_d_q_reg_30_ ( .D(n16), .CK(n37805), .RN(n38343), .QN(
        n56374) );
  DFFRX1 u_fetch_pc_d_q_reg_26_ ( .D(n13), .CK(n37805), .RN(n38337), .QN(
        n54376) );
  DFFRX1 u_fetch_pc_d_q_reg_22_ ( .D(n17), .CK(n37805), .RN(n38362), .QN(
        n55628) );
  DFFRX1 u_fetch_pc_d_q_reg_14_ ( .D(n24), .CK(n37804), .RN(n38361), .QN(
        n55195) );
  DFFRX1 u_fetch_pc_d_q_reg_29_ ( .D(n14), .CK(n37805), .RN(n38317), .QN(
        n56183) );
  DFFRX1 u_fetch_pc_d_q_reg_20_ ( .D(n7), .CK(n37805), .RN(n38360), .QN(n55526) );
  DFFRX1 u_fetch_pc_d_q_reg_16_ ( .D(n8), .CK(n37805), .RN(n38359), .QN(n55316) );
  DFFRX1 u_fetch_pc_d_q_reg_27_ ( .D(n19), .CK(n37805), .RN(n38316), .QN(
        n55997) );
  DFFRX1 u_fetch_pc_d_q_reg_15_ ( .D(n22), .CK(n37804), .RN(n38362), .QN(
        n55256) );
  DFFRX1 u_decode_inst_q_reg_13_ ( .D(n42425), .CK(n37870), .RN(n38361), .Q(
        opcode_opcode_w[13]), .QN(n56868) );
  DFFRX1 u_fetch_pc_d_q_reg_25_ ( .D(n23), .CK(n37805), .RN(n38342), .QN(
        n55772) );
  DFFRX1 u_fetch_pc_d_q_reg_1_ ( .D(mem_i_pc_o[1]), .CK(n37804), .RN(n38341), 
        .QN(n56781) );
  DFFRX1 u_fetch_pc_d_q_reg_0_ ( .D(mem_i_pc_o[0]), .CK(n37804), .RN(n38347), 
        .QN(n57283) );
  DFFRX1 u_fetch_pc_d_q_reg_10_ ( .D(mem_i_pc_o[10]), .CK(n37804), .RN(n38360), 
        .QN(n54963) );
  DFFRX1 u_fetch_pc_d_q_reg_6_ ( .D(mem_i_pc_o[6]), .CK(n37804), .RN(n38336), 
        .QN(n54715) );
  DFFRX1 u_fetch_pc_d_q_reg_11_ ( .D(mem_i_pc_o[11]), .CK(n37804), .RN(n38359), 
        .QN(n55028) );
  DFFRX1 u_fetch_pc_d_q_reg_7_ ( .D(mem_i_pc_o[7]), .CK(n37804), .RN(n38335), 
        .QN(n54775) );
  DFFRX1 u_fetch_pc_d_q_reg_8_ ( .D(mem_i_pc_o[8]), .CK(n37804), .RN(n38340), 
        .QN(n56811) );
  DFFRX1 u_fetch_pc_d_q_reg_4_ ( .D(mem_i_pc_o[4]), .CK(n37804), .RN(n38338), 
        .QN(n54581) );
  DFFRX1 u_fetch_pc_d_q_reg_5_ ( .D(mem_i_pc_o[5]), .CK(n37804), .RN(n38337), 
        .QN(n54652) );
  DFFRX1 u_fetch_pc_d_q_reg_3_ ( .D(mem_i_pc_o[3]), .CK(n37804), .RN(n38343), 
        .QN(n56789) );
  DFFRX1 u_fetch_pc_d_q_reg_9_ ( .D(mem_i_pc_o[9]), .CK(n37804), .RN(n38362), 
        .QN(n54892) );
  DFFRX1 u_decode_inst_q_reg_14_ ( .D(n42424), .CK(n37870), .RN(n38361), .Q(
        opcode_opcode_w[14]), .QN(n56876) );
  DFFRX1 u_fetch_pc_d_q_reg_2_ ( .D(mem_i_pc_o[2]), .CK(n37804), .RN(n38336), 
        .QN(n54440) );
  DFFRX1 u_fetch_pc_d_q_reg_18_ ( .D(n10), .CK(n37805), .RN(n38360), .QN(
        n55421) );
  DFFRX1 u_fetch_pc_d_q_reg_28_ ( .D(n18), .CK(n37805), .RN(n38315), .QN(
        n56173) );
  DFFRX1 u_fetch_pc_d_q_reg_23_ ( .D(n15), .CK(n37805), .RN(n38359), .QN(
        n55676) );
  DFFRX1 u_fetch_pc_d_q_reg_19_ ( .D(n20), .CK(n37805), .RN(n38362), .QN(
        n55473) );
  DFFRX1 u_fetch_pc_d_q_reg_17_ ( .D(n6), .CK(n37805), .RN(n38361), .QN(n55367) );
  DFFRX1 u_fetch_pc_d_q_reg_24_ ( .D(n11), .CK(n37805), .RN(n38342), .QN(
        n55724) );
  DFFRX1 u_fetch_pc_d_q_reg_21_ ( .D(n12), .CK(n37805), .RN(n38360), .QN(
        n55578) );
  DFFRX1 u_fetch_pc_d_q_reg_13_ ( .D(n9), .CK(n37804), .RN(n38359), .QN(n55139) );
  DFFRX1 u_muldiv_mult_result_q_reg_7_ ( .D(u_muldiv_result_r[7]), .CK(clk_i), 
        .RN(n38346), .Q(u_muldiv_mult_result_q[7]) );
  DFFRX1 u_decode_inst_q_reg_25_ ( .D(n8514), .CK(clk_i), .RN(n38351), .Q(
        opcode_opcode_w[25]), .QN(n58817) );
  DFFRX1 u_decode_inst_q_reg_30_ ( .D(n8519), .CK(clk_i), .RN(n38350), .Q(
        opcode_opcode_w[30]), .QN(n57889) );
  DFFRX1 u_decode_inst_q_reg_26_ ( .D(n8515), .CK(clk_i), .RN(n38349), .Q(
        opcode_opcode_w[26]), .QN(n73364) );
  DFFRX1 u_decode_inst_q_reg_27_ ( .D(n8516), .CK(clk_i), .RN(n38352), .Q(
        opcode_opcode_w[27]), .QN(n58818) );
  DFFRX1 u_decode_inst_q_reg_31_ ( .D(n8538), .CK(clk_i), .RN(n38351), .Q(
        opcode_opcode_w[31]), .QN(n44832) );
  DFFRX1 u_decode_opcode_instr_q_reg_55_ ( .D(u_decode_N791), .CK(n37885), 
        .RN(n44252), .Q(opcode_instr_w_55), .QN(n58212) );
  DFFRX1 u_decode_opcode_instr_q_reg_9_ ( .D(u_decode_N745), .CK(n37806), .RN(
        n38320), .QN(n50694) );
  DFFRX1 u_mmu_virt_addr_q_reg_14_ ( .D(u_mmu_request_addr_w[14]), .CK(n37803), 
        .RN(n38341), .Q(u_mmu_virt_addr_q[14]) );
  DFFRX1 u_mmu_virt_addr_q_reg_12_ ( .D(u_mmu_request_addr_w[12]), .CK(n37803), 
        .RN(n38340), .Q(u_mmu_virt_addr_q[12]) );
  DFFRX1 u_mmu_virt_addr_q_reg_20_ ( .D(u_mmu_request_addr_w[20]), .CK(n37803), 
        .RN(n38343), .Q(u_mmu_virt_addr_q[20]) );
  DFFRX1 u_mmu_virt_addr_q_reg_16_ ( .D(u_mmu_request_addr_w[16]), .CK(n37803), 
        .RN(n38342), .Q(u_mmu_virt_addr_q[16]) );
  DFFRX1 u_mmu_virt_addr_q_reg_15_ ( .D(u_mmu_request_addr_w[15]), .CK(n37803), 
        .RN(n38341), .Q(u_mmu_virt_addr_q[15]) );
  DFFRX1 u_decode_opcode_instr_q_reg_2_ ( .D(u_decode_N738), .CK(n37806), .RN(
        n38323), .Q(n1854), .QN(n50657) );
  DFFRX1 u_mmu_virt_addr_q_reg_18_ ( .D(u_mmu_request_addr_w[18]), .CK(n37803), 
        .RN(n38340), .Q(u_mmu_virt_addr_q[18]) );
  DFFRX1 u_mmu_virt_addr_q_reg_19_ ( .D(u_mmu_request_addr_w[19]), .CK(n37803), 
        .RN(n38343), .Q(u_mmu_virt_addr_q[19]) );
  DFFRX1 u_decode_opcode_instr_q_reg_42_ ( .D(u_decode_N778), .CK(n37807), 
        .RN(n38362), .Q(n1852) );
  DFFRX1 u_decode_opcode_instr_q_reg_31_ ( .D(u_decode_N767), .CK(n37802), 
        .RN(n38350), .Q(n1853), .QN(n58811) );
  DFFRX1 u_decode_opcode_instr_q_reg_13_ ( .D(u_decode_N749), .CK(n37806), 
        .RN(n38322), .QN(n50678) );
  DFFRX1 u_mmu_virt_addr_q_reg_17_ ( .D(u_mmu_request_addr_w[17]), .CK(n37803), 
        .RN(n38342), .Q(u_mmu_virt_addr_q[17]) );
  DFFRX1 u_decode_opcode_instr_q_reg_37_ ( .D(u_decode_N773), .CK(n37807), 
        .RN(n38335), .Q(opcode_instr_w_37), .QN(n58812) );
  DFFRX1 u_mmu_virt_addr_q_reg_21_ ( .D(u_mmu_request_addr_w[21]), .CK(n37803), 
        .RN(n38341), .Q(u_mmu_virt_addr_q[21]) );
  DFFRX1 u_mmu_virt_addr_q_reg_13_ ( .D(u_mmu_request_addr_w[13]), .CK(n37803), 
        .RN(n38340), .Q(u_mmu_virt_addr_q[13]) );
  DFFRX1 u_csr_csr_sepc_q_reg_2_ ( .D(u_csr_csr_sepc_r[2]), .CK(clk_i), .RN(
        n38338), .Q(u_csr_csr_sepc_q[2]), .QN(n58487) );
  DFFRX1 u_fetch_skid_buffer_q_reg_6_ ( .D(net2343), .CK(n37801), .RN(n38349), 
        .Q(u_fetch_skid_buffer_q[6]) );
  DFFRX1 u_fetch_skid_buffer_q_reg_4_ ( .D(net2341), .CK(n37801), .RN(n38352), 
        .Q(u_fetch_skid_buffer_q[4]) );
  DFFRX1 u_fetch_skid_buffer_q_reg_1_ ( .D(net2337), .CK(n37801), .RN(n38345), 
        .Q(u_fetch_skid_buffer_q[1]) );
  DFFRX1 u_fetch_skid_buffer_q_reg_0_ ( .D(net2336), .CK(n37801), .RN(n38344), 
        .Q(u_fetch_skid_buffer_q[0]) );
  DFFRX1 u_csr_csr_mepc_q_reg_0_ ( .D(u_csr_csr_mepc_r[0]), .CK(clk_i), .RN(
        n38347), .Q(u_csr_csr_mepc_q[0]), .QN(n58456) );
  DFFRX1 u_csr_csr_mepc_q_reg_1_ ( .D(u_csr_csr_mepc_r[1]), .CK(clk_i), .RN(
        n38355), .Q(u_csr_csr_mepc_q[1]), .QN(n58476) );
  DFFRX1 u_csr_csr_sepc_q_reg_0_ ( .D(u_csr_csr_sepc_r[0]), .CK(clk_i), .RN(
        n38346), .Q(u_csr_csr_sepc_q[0]), .QN(n58455) );
  DFFRX1 u_csr_csr_sepc_q_reg_1_ ( .D(u_csr_csr_sepc_r[1]), .CK(clk_i), .RN(
        n38354), .Q(u_csr_csr_sepc_q[1]), .QN(n58475) );
  DFFRX1 u_decode_opcode_instr_q_reg_47_ ( .D(u_decode_N783), .CK(n37807), 
        .RN(n44252), .Q(n1837) );
  DFFRX1 u_decode_opcode_instr_q_reg_29_ ( .D(u_decode_N765), .CK(n37802), 
        .RN(n38351), .QN(n73363) );
  DFFRX1 u_decode_opcode_instr_q_reg_23_ ( .D(u_decode_N759), .CK(n37802), 
        .RN(n38350), .Q(n1888), .QN(n50039) );
  DFFRX1 u_decode_opcode_instr_q_reg_11_ ( .D(u_decode_N747), .CK(n37806), 
        .RN(n38321), .Q(opcode_instr_w[11]), .QN(n50856) );
  DFFRX1 u_decode_opcode_instr_q_reg_1_ ( .D(u_decode_N737), .CK(n37806), .RN(
        n38320), .Q(opcode_instr_w_1), .QN(n58541) );
  DFFRX1 u_decode_opcode_instr_q_reg_35_ ( .D(u_decode_N771), .CK(n37807), 
        .RN(n38349), .Q(opcode_instr_w_35), .QN(n57360) );
  DFFRX1 u_csr_csr_mepc_q_reg_2_ ( .D(u_csr_csr_mepc_r[2]), .CK(clk_i), .RN(
        n38337), .Q(u_csr_csr_mepc_q[2]), .QN(n58488) );
  DFFRX1 u_decode_opcode_instr_q_reg_54_ ( .D(u_decode_N790), .CK(n37885), 
        .RN(n44252), .Q(n1891) );
  DFFRX1 u_decode_opcode_instr_q_reg_46_ ( .D(u_decode_N782), .CK(n37807), 
        .RN(n38336), .Q(opcode_instr_w_46) );
  DFFRX1 u_decode_opcode_instr_q_reg_28_ ( .D(u_decode_N764), .CK(n37802), 
        .RN(n38352), .Q(opcode_instr_w_28) );
  DFFRX1 u_decode_opcode_instr_q_reg_17_ ( .D(u_decode_N753), .CK(n37802), 
        .RN(n38323), .Q(opcode_instr_w_17), .QN(n50850) );
  DFFRX1 u_decode_opcode_instr_q_reg_0_ ( .D(u_decode_N736), .CK(n37806), .RN(
        n38322), .QN(n50658) );
  DFFRX1 u_decode_opcode_instr_q_reg_41_ ( .D(u_decode_N777), .CK(n37807), 
        .RN(n38321), .Q(opcode_instr_w_41), .QN(n55034) );
  DFFRX1 u_decode_opcode_instr_q_reg_30_ ( .D(u_decode_N766), .CK(n37802), 
        .RN(n38351), .Q(n1855) );
  DFFRX1 u_decode_opcode_instr_q_reg_24_ ( .D(u_decode_N760), .CK(n37802), 
        .RN(n38345), .Q(opcode_instr_w_24) );
  DFFRX1 u_decode_opcode_instr_q_reg_6_ ( .D(u_decode_N742), .CK(n37806), .RN(
        n38320), .Q(opcode_instr_w[6]), .QN(n57096) );
  DFFRX1 u_decode_opcode_instr_q_reg_36_ ( .D(u_decode_N772), .CK(n37807), 
        .RN(n38335), .Q(opcode_instr_w_36) );
  DFFRX1 u_decode_opcode_instr_q_reg_51_ ( .D(u_decode_N787), .CK(n37885), 
        .RN(n44252), .Q(opcode_instr_w_51), .QN(n58164) );
  DFFRX1 u_decode_opcode_instr_q_reg_25_ ( .D(u_decode_N761), .CK(n37802), 
        .RN(n38344), .Q(opcode_instr_w_25), .QN(n50028) );
  DFFRX1 u_decode_opcode_instr_q_reg_15_ ( .D(u_decode_N751), .CK(n37806), 
        .RN(n38323), .Q(n1926), .QN(n50682) );
  DFFRX1 u_decode_opcode_instr_q_reg_5_ ( .D(u_decode_N741), .CK(n37806), .RN(
        n38322), .Q(opcode_instr_w[5]) );
  DFFRX1 u_muldiv_mult_result_q_reg_8_ ( .D(u_muldiv_result_r[8]), .CK(clk_i), 
        .RN(n38347), .Q(u_muldiv_mult_result_q[8]) );
  DFFRX1 u_decode_opcode_instr_q_reg_53_ ( .D(u_decode_N789), .CK(n37885), 
        .RN(n44252), .Q(n8887), .QN(n44954) );
  DFFRX1 u_decode_opcode_instr_q_reg_45_ ( .D(u_decode_N781), .CK(n37807), 
        .RN(n38338), .Q(opcode_instr_w_45) );
  DFFRX1 u_decode_opcode_instr_q_reg_34_ ( .D(u_decode_N770), .CK(n37807), 
        .RN(n38350), .Q(n1850), .QN(n58815) );
  DFFRX1 u_decode_opcode_instr_q_reg_27_ ( .D(u_decode_N763), .CK(n37802), 
        .RN(n38349), .Q(n36761), .QN(n44810) );
  DFFRX1 u_decode_opcode_instr_q_reg_16_ ( .D(u_decode_N752), .CK(n37802), 
        .RN(n38321), .Q(opcode_instr_w_16), .QN(n50859) );
  DFFRX1 u_decode_opcode_instr_q_reg_52_ ( .D(u_decode_N788), .CK(n37885), 
        .RN(n44252), .Q(n1848), .QN(n58165) );
  DFFRX1 u_decode_opcode_instr_q_reg_44_ ( .D(u_decode_N780), .CK(n37807), 
        .RN(n38337), .QN(n55033) );
  DFFRX1 u_decode_opcode_instr_q_reg_33_ ( .D(u_decode_N769), .CK(n37807), 
        .RN(n38352), .Q(n1849) );
  DFFRX1 u_csr_csr_sepc_q_reg_14_ ( .D(u_csr_csr_sepc_r[14]), .CK(clk_i), .RN(
        n38361), .Q(u_csr_csr_sepc_q[14]), .QN(n55182) );
  DFFRX1 u_csr_csr_sepc_q_reg_12_ ( .D(u_csr_csr_sepc_r[12]), .CK(clk_i), .RN(
        n38360), .Q(u_csr_csr_sepc_q[12]), .QN(n55078) );
  DFFRX1 u_csr_csr_sepc_q_reg_15_ ( .D(u_csr_csr_sepc_r[15]), .CK(clk_i), .RN(
        n38359), .Q(u_csr_csr_sepc_q[15]), .QN(n55242) );
  DFFRX1 u_csr_csr_sepc_q_reg_10_ ( .D(u_csr_csr_sepc_r[10]), .CK(clk_i), .RN(
        n38362), .Q(u_csr_csr_sepc_q[10]), .QN(n58463) );
  DFFRX1 u_csr_csr_sepc_q_reg_8_ ( .D(u_csr_csr_sepc_r[8]), .CK(clk_i), .RN(
        n44248), .Q(u_csr_csr_sepc_q[8]), .QN(n58502) );
  DFFRX1 u_decode_opcode_instr_q_reg_57_ ( .D(u_decode_N793), .CK(n37885), 
        .RN(n44252), .Q(opcode_instr_w_57) );
  DFFRX1 u_mmu_pte_entry_q_reg_12_ ( .D(u_mmu_N239), .CK(net1802), .RN(n44252), 
        .Q(u_mmu_pte_entry_q[12]) );
  DFFRX1 u_mmu_pte_entry_q_reg_14_ ( .D(u_mmu_N241), .CK(net1802), .RN(n44252), 
        .Q(u_mmu_pte_entry_q[14]) );
  DFFRX1 u_mmu_pte_entry_q_reg_16_ ( .D(u_mmu_N243), .CK(net1802), .RN(n38346), 
        .Q(u_mmu_pte_entry_q[16]) );
  DFFRX1 u_mmu_pte_entry_q_reg_20_ ( .D(u_mmu_N247), .CK(net1802), .RN(n38318), 
        .Q(u_mmu_pte_entry_q[20]) );
  DFFRX1 u_mmu_pte_entry_q_reg_15_ ( .D(u_mmu_N242), .CK(net1802), .RN(n44252), 
        .Q(u_mmu_pte_entry_q[15]) );
  DFFRX1 u_decode_opcode_instr_q_reg_40_ ( .D(u_decode_N776), .CK(n37807), 
        .RN(n38357), .Q(opcode_instr_w_40), .QN(n58211) );
  DFFRX1 u_mmu_pte_entry_q_reg_18_ ( .D(u_mmu_N245), .CK(net1802), .RN(n38317), 
        .Q(u_mmu_pte_entry_q[18]) );
  DFFRX1 u_mmu_pte_entry_q_reg_19_ ( .D(u_mmu_N246), .CK(net1802), .RN(n38316), 
        .Q(u_mmu_pte_entry_q[19]) );
  DFFRX1 u_mmu_pte_entry_q_reg_17_ ( .D(u_mmu_N244), .CK(net1802), .RN(n38315), 
        .Q(u_mmu_pte_entry_q[17]) );
  DFFRX1 u_muldiv_mult_result_q_reg_9_ ( .D(u_muldiv_result_r[9]), .CK(clk_i), 
        .RN(n38345), .Q(u_muldiv_mult_result_q[9]) );
  DFFRX1 u_decode_pc_q_reg_31_ ( .D(u_decode_N321), .CK(n37800), .RN(n38343), 
        .Q(opcode_pc_w[31]), .QN(n58416) );
  DFFRX1 u_decode_pc_q_reg_30_ ( .D(u_decode_N320), .CK(n37800), .RN(n38342), 
        .Q(opcode_pc_w[30]), .QN(n58409) );
  DFFRX1 u_decode_pc_q_reg_8_ ( .D(u_decode_N298), .CK(n37799), .RN(n38341), 
        .Q(opcode_pc_w[8]), .QN(n58441) );
  DFFRX1 u_decode_pc_q_reg_29_ ( .D(u_decode_N319), .CK(n37800), .RN(n38318), 
        .Q(opcode_pc_w[29]), .QN(n58403) );
  DFFRX1 u_decode_pc_q_reg_28_ ( .D(u_decode_N318), .CK(n37800), .RN(n38317), 
        .Q(opcode_pc_w[28]), .QN(n58396) );
  DFFRX1 u_decode_pc_q_reg_3_ ( .D(u_decode_N293), .CK(n37799), .RN(n38340), 
        .Q(opcode_pc_w[3]), .QN(n54529) );
  DFFRX1 u_decode_pc_q_reg_1_ ( .D(u_decode_N291), .CK(n37799), .RN(n38343), 
        .Q(opcode_pc_w[1]), .QN(n56782) );
  DFFRX1 u_decode_pc_q_reg_0_ ( .D(u_decode_N290), .CK(n37799), .RN(n38344), 
        .Q(u_csr_N184), .QN(n57284) );
  DFFRX1 u_mmu_pte_entry_q_reg_21_ ( .D(u_mmu_N248), .CK(net1802), .RN(n38316), 
        .Q(u_mmu_pte_entry_q[21]) );
  DFFRX1 u_mmu_pte_entry_q_reg_13_ ( .D(u_mmu_N240), .CK(net1802), .RN(n44252), 
        .Q(u_mmu_pte_entry_q[13]) );
  DFFRX1 u_csr_csr_mepc_q_reg_18_ ( .D(u_csr_csr_mepc_r[18]), .CK(clk_i), .RN(
        n38361), .Q(u_csr_csr_mepc_q[18]), .QN(n55406) );
  DFFRX1 u_csr_csr_mepc_q_reg_5_ ( .D(u_csr_csr_mepc_r[5]), .CK(clk_i), .RN(
        n38336), .Q(u_csr_csr_mepc_q[5]), .QN(n58496) );
  DFFRX1 u_csr_csr_mepc_q_reg_7_ ( .D(u_csr_csr_mepc_r[7]), .CK(clk_i), .RN(
        n38335), .Q(u_csr_csr_mepc_q[7]), .QN(n58500) );
  DFFRX1 u_csr_csr_mepc_q_reg_3_ ( .D(u_csr_csr_mepc_r[3]), .CK(clk_i), .RN(
        n38338), .Q(u_csr_csr_mepc_q[3]), .QN(n58492) );
  DFFRX1 u_csr_csr_mepc_q_reg_4_ ( .D(u_csr_csr_mepc_r[4]), .CK(clk_i), .RN(
        n38337), .Q(u_csr_csr_mepc_q[4]), .QN(n58494) );
  DFFRX1 u_csr_csr_mepc_q_reg_6_ ( .D(u_csr_csr_mepc_r[6]), .CK(clk_i), .RN(
        n38336), .Q(u_csr_csr_mepc_q[6]), .QN(n58498) );
  DFFRX1 u_csr_csr_sepc_q_reg_18_ ( .D(u_csr_csr_sepc_r[18]), .CK(clk_i), .RN(
        n38360), .Q(u_csr_csr_sepc_q[18]), .QN(n55407) );
  DFFRX1 u_csr_csr_mepc_q_reg_21_ ( .D(u_csr_csr_mepc_r[21]), .CK(clk_i), .RN(
        n38359), .Q(u_csr_csr_mepc_q[21]), .QN(n55565) );
  DFFRX1 u_csr_csr_mepc_q_reg_20_ ( .D(u_csr_csr_mepc_r[20]), .CK(clk_i), .RN(
        n38362), .Q(u_csr_csr_mepc_q[20]), .QN(n55512) );
  DFFRX1 u_csr_csr_mepc_q_reg_17_ ( .D(u_csr_csr_mepc_r[17]), .CK(clk_i), .RN(
        n38361), .Q(u_csr_csr_mepc_q[17]), .QN(n55354) );
  DFFRX1 u_csr_csr_mepc_q_reg_16_ ( .D(u_csr_csr_mepc_r[16]), .CK(clk_i), .RN(
        n38360), .Q(u_csr_csr_mepc_q[16]), .QN(n55294) );
  DFFRX1 u_csr_csr_mepc_q_reg_14_ ( .D(u_csr_csr_mepc_r[14]), .CK(clk_i), .RN(
        n38359), .Q(u_csr_csr_mepc_q[14]), .QN(n55181) );
  DFFRX1 u_csr_csr_mepc_q_reg_13_ ( .D(u_csr_csr_mepc_r[13]), .CK(clk_i), .RN(
        n38362), .Q(u_csr_csr_mepc_q[13]), .QN(n55126) );
  DFFRX1 u_csr_csr_mepc_q_reg_12_ ( .D(u_csr_csr_mepc_r[12]), .CK(clk_i), .RN(
        n38361), .Q(u_csr_csr_mepc_q[12]), .QN(n55077) );
  DFFRX1 u_csr_csr_mepc_q_reg_19_ ( .D(u_csr_csr_mepc_r[19]), .CK(clk_i), .RN(
        n38360), .Q(u_csr_csr_mepc_q[19]), .QN(n55457) );
  DFFRX1 u_csr_csr_mepc_q_reg_15_ ( .D(u_csr_csr_mepc_r[15]), .CK(clk_i), .RN(
        n38359), .Q(u_csr_csr_mepc_q[15]), .QN(n55241) );
  DFFRX1 u_csr_csr_mepc_q_reg_26_ ( .D(u_csr_csr_mepc_r[26]), .CK(clk_i), .RN(
        n38342), .Q(u_csr_csr_mepc_q[26]), .QN(n55806) );
  DFFRX1 u_csr_csr_mepc_q_reg_25_ ( .D(u_csr_csr_mepc_r[25]), .CK(clk_i), .RN(
        n38341), .Q(u_csr_csr_mepc_q[25]), .QN(n55760) );
  DFFRX1 u_csr_csr_mepc_q_reg_24_ ( .D(u_csr_csr_mepc_r[24]), .CK(clk_i), .RN(
        n38335), .Q(u_csr_csr_mepc_q[24]), .QN(n55712) );
  DFFRX1 u_csr_csr_mepc_q_reg_23_ ( .D(u_csr_csr_mepc_r[23]), .CK(clk_i), .RN(
        n38362), .Q(u_csr_csr_mepc_q[23]), .QN(n55661) );
  DFFRX1 u_csr_csr_mepc_q_reg_22_ ( .D(u_csr_csr_mepc_r[22]), .CK(clk_i), .RN(
        n38361), .Q(u_csr_csr_mepc_q[22]), .QN(n55614) );
  DFFRX1 u_csr_csr_mepc_q_reg_31_ ( .D(u_csr_csr_mepc_r[31]), .CK(clk_i), .RN(
        n38340), .Q(u_csr_csr_mepc_q[31]), .QN(n58490) );
  DFFRX1 u_csr_csr_mepc_q_reg_30_ ( .D(u_csr_csr_mepc_r[30]), .CK(clk_i), .RN(
        n38343), .Q(u_csr_csr_mepc_q[30]), .QN(n58489) );
  DFFRX1 u_csr_csr_mepc_q_reg_29_ ( .D(u_csr_csr_mepc_r[29]), .CK(clk_i), .RN(
        n38315), .Q(u_csr_csr_mepc_q[29]), .QN(n56343) );
  DFFRX1 u_csr_csr_mepc_q_reg_28_ ( .D(u_csr_csr_mepc_r[28]), .CK(clk_i), .RN(
        n38318), .Q(u_csr_csr_mepc_q[28]), .QN(n56160) );
  DFFRX1 u_csr_csr_mepc_q_reg_27_ ( .D(u_csr_csr_mepc_r[27]), .CK(clk_i), .RN(
        n38317), .Q(u_csr_csr_mepc_q[27]), .QN(n55983) );
  DFFRX1 u_csr_csr_mepc_q_reg_9_ ( .D(u_csr_csr_mepc_r[9]), .CK(clk_i), .RN(
        n44248), .Q(u_csr_csr_mepc_q[9]), .QN(n58505) );
  DFFRX1 u_csr_csr_mepc_q_reg_10_ ( .D(u_csr_csr_mepc_r[10]), .CK(clk_i), .RN(
        n38360), .Q(u_csr_csr_mepc_q[10]), .QN(n58464) );
  DFFRX1 u_csr_csr_mepc_q_reg_8_ ( .D(u_csr_csr_mepc_r[8]), .CK(clk_i), .RN(
        n44248), .Q(u_csr_csr_mepc_q[8]), .QN(n58503) );
  DFFRX1 u_csr_csr_mepc_q_reg_11_ ( .D(u_csr_csr_mepc_r[11]), .CK(clk_i), .RN(
        n38359), .Q(u_csr_csr_mepc_q[11]), .QN(n58466) );
  DFFRX1 u_csr_csr_sepc_q_reg_30_ ( .D(u_csr_csr_sepc_r[30]), .CK(clk_i), .RN(
        n38342), .Q(u_csr_csr_sepc_q[30]), .QN(n56536) );
  DFFRX1 u_csr_csr_sepc_q_reg_29_ ( .D(u_csr_csr_sepc_r[29]), .CK(clk_i), .RN(
        n38316), .Q(u_csr_csr_sepc_q[29]), .QN(n58486) );
  DFFRX1 u_csr_csr_sepc_q_reg_28_ ( .D(u_csr_csr_sepc_r[28]), .CK(clk_i), .RN(
        n38315), .Q(u_csr_csr_sepc_q[28]), .QN(n58485) );
  DFFRX1 u_csr_csr_sepc_q_reg_27_ ( .D(u_csr_csr_sepc_r[27]), .CK(clk_i), .RN(
        n38318), .Q(u_csr_csr_sepc_q[27]), .QN(n58484) );
  DFFRX1 u_csr_csr_sepc_q_reg_26_ ( .D(u_csr_csr_sepc_r[26]), .CK(clk_i), .RN(
        n38317), .Q(u_csr_csr_sepc_q[26]), .QN(n58483) );
  DFFRX1 u_csr_csr_sepc_q_reg_25_ ( .D(u_csr_csr_sepc_r[25]), .CK(clk_i), .RN(
        n38341), .Q(u_csr_csr_sepc_q[25]), .QN(n58482) );
  DFFRX1 u_csr_csr_sepc_q_reg_24_ ( .D(u_csr_csr_sepc_r[24]), .CK(clk_i), .RN(
        n38316), .Q(u_csr_csr_sepc_q[24]), .QN(n58481) );
  DFFRX1 u_csr_csr_sepc_q_reg_23_ ( .D(u_csr_csr_sepc_r[23]), .CK(clk_i), .RN(
        n38362), .Q(u_csr_csr_sepc_q[23]), .QN(n58480) );
  DFFRX1 u_csr_csr_sepc_q_reg_22_ ( .D(u_csr_csr_sepc_r[22]), .CK(clk_i), .RN(
        n38361), .Q(u_csr_csr_sepc_q[22]), .QN(n58479) );
  DFFRX1 u_csr_csr_sepc_q_reg_21_ ( .D(u_csr_csr_sepc_r[21]), .CK(clk_i), .RN(
        n38360), .Q(u_csr_csr_sepc_q[21]), .QN(n55566) );
  DFFRX1 u_csr_csr_sepc_q_reg_20_ ( .D(u_csr_csr_sepc_r[20]), .CK(clk_i), .RN(
        n38359), .Q(u_csr_csr_sepc_q[20]), .QN(n55513) );
  DFFRX1 u_csr_csr_sepc_q_reg_19_ ( .D(u_csr_csr_sepc_r[19]), .CK(clk_i), .RN(
        n38362), .Q(u_csr_csr_sepc_q[19]), .QN(n55458) );
  DFFRX1 u_csr_csr_sepc_q_reg_17_ ( .D(u_csr_csr_sepc_r[17]), .CK(clk_i), .RN(
        n38361), .Q(u_csr_csr_sepc_q[17]), .QN(n55355) );
  DFFRX1 u_csr_csr_sepc_q_reg_16_ ( .D(u_csr_csr_sepc_r[16]), .CK(clk_i), .RN(
        n38360), .Q(u_csr_csr_sepc_q[16]), .QN(n55295) );
  DFFRX1 u_csr_csr_sepc_q_reg_13_ ( .D(u_csr_csr_sepc_r[13]), .CK(clk_i), .RN(
        n38359), .Q(u_csr_csr_sepc_q[13]), .QN(n55127) );
  DFFRX1 u_csr_csr_sepc_q_reg_6_ ( .D(u_csr_csr_sepc_r[6]), .CK(clk_i), .RN(
        n38338), .Q(u_csr_csr_sepc_q[6]), .QN(n58497) );
  DFFRX1 u_csr_csr_sepc_q_reg_5_ ( .D(u_csr_csr_sepc_r[5]), .CK(clk_i), .RN(
        n38337), .Q(u_csr_csr_sepc_q[5]), .QN(n58495) );
  DFFRX1 u_csr_csr_sepc_q_reg_7_ ( .D(u_csr_csr_sepc_r[7]), .CK(clk_i), .RN(
        n38336), .Q(u_csr_csr_sepc_q[7]), .QN(n58499) );
  DFFRX1 u_csr_csr_sepc_q_reg_4_ ( .D(u_csr_csr_sepc_r[4]), .CK(clk_i), .RN(
        n38335), .Q(u_csr_csr_sepc_q[4]), .QN(n58493) );
  DFFRX1 u_csr_csr_sepc_q_reg_3_ ( .D(u_csr_csr_sepc_r[3]), .CK(clk_i), .RN(
        n38338), .Q(u_csr_csr_sepc_q[3]), .QN(n58491) );
  DFFRX1 u_csr_csr_sepc_q_reg_9_ ( .D(u_csr_csr_sepc_r[9]), .CK(clk_i), .RN(
        n44248), .Q(u_csr_csr_sepc_q[9]), .QN(n58504) );
  DFFRX1 u_decode_opcode_instr_q_reg_43_ ( .D(u_decode_N779), .CK(n37807), 
        .RN(n38347), .Q(n40925) );
  DFFRX1 u_decode_opcode_instr_q_reg_3_ ( .D(u_decode_N739), .CK(n37806), .RN(
        n38320), .Q(n1890) );
  DFFRX1 u_decode_opcode_instr_q_reg_50_ ( .D(u_decode_N786), .CK(n37885), 
        .RN(n44252), .Q(n42546) );
  DFFRX1 u_decode_opcode_instr_q_reg_14_ ( .D(u_decode_N750), .CK(n37806), 
        .RN(n38323), .QN(n58540) );
  DFFRX1 u_csr_csr_sepc_q_reg_31_ ( .D(u_csr_csr_sepc_r[31]), .CK(clk_i), .RN(
        n38340), .Q(u_csr_csr_sepc_q[31]), .QN(n56607) );
  DFFRX1 u_csr_csr_sepc_q_reg_11_ ( .D(u_csr_csr_sepc_r[11]), .CK(clk_i), .RN(
        n38362), .Q(u_csr_csr_sepc_q[11]), .QN(n58465) );
  DFFRX1 u_fetch_skid_buffer_q_reg_19_ ( .D(net2361), .CK(n37798), .RN(n38322), 
        .Q(u_fetch_skid_buffer_q[19]) );
  DFFRX1 u_fetch_skid_buffer_q_reg_18_ ( .D(net2360), .CK(n37798), .RN(n44252), 
        .QN(n57599) );
  DFFRX1 u_fetch_skid_buffer_q_reg_31_ ( .D(net2374), .CK(n37798), .RN(n38351), 
        .Q(u_fetch_skid_buffer_q[31]) );
  DFFRX1 u_fetch_skid_buffer_q_reg_30_ ( .D(net2373), .CK(n37798), .RN(n38350), 
        .Q(u_fetch_skid_buffer_q[30]) );
  DFFRX1 u_fetch_skid_buffer_q_reg_29_ ( .D(net2372), .CK(n37798), .RN(n38349), 
        .Q(u_fetch_skid_buffer_q[29]) );
  DFFRX1 u_fetch_skid_buffer_q_reg_26_ ( .D(net2368), .CK(n37798), .RN(n38352), 
        .Q(u_fetch_skid_buffer_q[26]) );
  DFFRX1 u_fetch_skid_buffer_q_reg_24_ ( .D(net2366), .CK(n37798), .RN(n38351), 
        .Q(u_fetch_skid_buffer_q[24]) );
  DFFRX1 u_fetch_skid_buffer_q_reg_23_ ( .D(net2365), .CK(n37798), .RN(n38350), 
        .Q(u_fetch_skid_buffer_q[23]) );
  DFFRX1 u_fetch_skid_buffer_q_reg_17_ ( .D(net2359), .CK(n37798), .RN(n38349), 
        .Q(u_fetch_skid_buffer_q[17]) );
  DFFRX1 u_fetch_skid_buffer_q_reg_10_ ( .D(net2347), .CK(n37801), .RN(n38352), 
        .Q(u_fetch_skid_buffer_q[10]) );
  DFFRX1 u_fetch_skid_buffer_q_reg_9_ ( .D(net2346), .CK(n37801), .RN(n38351), 
        .Q(u_fetch_skid_buffer_q[9]) );
  DFFRX1 u_fetch_skid_buffer_q_reg_8_ ( .D(net2345), .CK(n37801), .RN(n38350), 
        .Q(u_fetch_skid_buffer_q[8]) );
  DFFRX1 u_fetch_skid_buffer_q_reg_2_ ( .D(net2339), .CK(n37801), .RN(n38346), 
        .Q(u_fetch_skid_buffer_q[2]) );
  DFFRX1 u_decode_pc_q_reg_9_ ( .D(u_decode_N299), .CK(n37799), .RN(n38361), 
        .Q(opcode_pc_w[9]), .QN(n58446) );
  DFFRX1 u_decode_pc_q_reg_7_ ( .D(u_decode_N297), .CK(n37799), .RN(n38360), 
        .Q(opcode_pc_w[7]), .QN(n58436) );
  DFFRX1 u_decode_pc_q_reg_4_ ( .D(u_decode_N294), .CK(n37799), .RN(n38337), 
        .Q(opcode_pc_w[4]), .QN(n54591) );
  DFFRX1 u_decode_pc_q_reg_23_ ( .D(u_decode_N313), .CK(n37800), .RN(n38359), 
        .Q(opcode_pc_w[23]), .QN(n58363) );
  DFFRX1 u_decode_pc_q_reg_15_ ( .D(u_decode_N305), .CK(n37799), .RN(n38362), 
        .Q(opcode_pc_w[15]), .QN(n58312) );
  DFFRX1 u_decode_pc_q_reg_14_ ( .D(u_decode_N304), .CK(n37799), .RN(n38361), 
        .Q(opcode_pc_w[14]), .QN(n58305) );
  DFFRX1 u_decode_pc_q_reg_13_ ( .D(u_decode_N303), .CK(n37799), .RN(n38360), 
        .Q(opcode_pc_w[13]), .QN(n58298) );
  DFFRX1 u_decode_pc_q_reg_12_ ( .D(u_decode_N302), .CK(n37799), .RN(n38359), 
        .Q(opcode_pc_w[12]), .QN(n58291) );
  DFFRX1 u_decode_pc_q_reg_11_ ( .D(u_decode_N301), .CK(n37799), .RN(n38362), 
        .Q(opcode_pc_w[11]), .QN(n58286) );
  DFFRX1 u_decode_pc_q_reg_10_ ( .D(u_decode_N300), .CK(n37799), .RN(n38361), 
        .Q(opcode_pc_w[10]), .QN(n58280) );
  DFFRX1 u_decode_pc_q_reg_22_ ( .D(u_decode_N312), .CK(n37800), .RN(n38360), 
        .Q(opcode_pc_w[22]), .QN(n58356) );
  DFFRX1 u_decode_pc_q_reg_24_ ( .D(u_decode_N314), .CK(n37800), .RN(n38343), 
        .Q(opcode_pc_w[24]), .QN(n58370) );
  DFFRX1 u_decode_pc_q_reg_20_ ( .D(u_decode_N310), .CK(n37800), .RN(n38359), 
        .Q(opcode_pc_w[20]), .QN(n58344) );
  DFFRX1 u_decode_pc_q_reg_18_ ( .D(u_decode_N308), .CK(n37800), .RN(n38362), 
        .Q(opcode_pc_w[18]), .QN(n58331) );
  DFFRX1 u_decode_pc_q_reg_27_ ( .D(u_decode_N317), .CK(n37800), .RN(n38315), 
        .Q(opcode_pc_w[27]), .QN(n58389) );
  DFFRX1 u_decode_pc_q_reg_26_ ( .D(u_decode_N316), .CK(n37800), .RN(n38336), 
        .Q(opcode_pc_w[26]), .QN(n58382) );
  DFFRX1 u_decode_pc_q_reg_25_ ( .D(u_decode_N315), .CK(n37800), .RN(n38342), 
        .Q(opcode_pc_w[25]), .QN(n58377) );
  DFFRX1 u_decode_pc_q_reg_21_ ( .D(u_decode_N311), .CK(n37800), .RN(n38361), 
        .Q(opcode_pc_w[21]), .QN(n58349) );
  DFFRX1 u_decode_pc_q_reg_17_ ( .D(u_decode_N307), .CK(n37800), .RN(n38360), 
        .Q(opcode_pc_w[17]), .QN(n58324) );
  DFFRX1 u_decode_pc_q_reg_16_ ( .D(u_decode_N306), .CK(n37800), .RN(n38359), 
        .Q(opcode_pc_w[16]), .QN(n58319) );
  DFFRX1 u_fetch_skid_buffer_q_reg_28_ ( .D(net2371), .CK(n37798), .RN(n38349), 
        .Q(u_fetch_skid_buffer_q[28]) );
  DFFRX1 u_fetch_skid_buffer_q_reg_25_ ( .D(net2367), .CK(n37798), .RN(n38352), 
        .Q(u_fetch_skid_buffer_q[25]) );
  DFFRX1 u_fetch_skid_buffer_q_reg_22_ ( .D(net2364), .CK(n37798), .RN(n38351), 
        .Q(u_fetch_skid_buffer_q[22]) );
  DFFRX1 u_fetch_skid_buffer_q_reg_21_ ( .D(net2363), .CK(n37798), .RN(n38350), 
        .Q(u_fetch_skid_buffer_q[21]) );
  DFFRX1 u_fetch_skid_buffer_q_reg_20_ ( .D(net2362), .CK(n37798), .RN(n38349), 
        .Q(u_fetch_skid_buffer_q[20]), .QN(n58513) );
  DFFRX1 u_fetch_skid_buffer_q_reg_16_ ( .D(net2358), .CK(n37798), .RN(n38352), 
        .QN(n50503) );
  DFFRX1 u_fetch_skid_buffer_q_reg_15_ ( .D(net2352), .CK(n37801), .RN(n44252), 
        .QN(n57549) );
  DFFRX1 u_fetch_skid_buffer_q_reg_14_ ( .D(net2351), .CK(n37801), .RN(n38351), 
        .Q(u_fetch_skid_buffer_q[14]) );
  DFFRX1 u_fetch_skid_buffer_q_reg_13_ ( .D(net2350), .CK(n37801), .RN(n38350), 
        .Q(u_fetch_skid_buffer_q[13]) );
  DFFRX1 u_fetch_skid_buffer_q_reg_12_ ( .D(net2349), .CK(n37801), .RN(n38349), 
        .Q(u_fetch_skid_buffer_q[12]) );
  DFFRX1 u_fetch_skid_buffer_q_reg_11_ ( .D(net2348), .CK(n37801), .RN(n38352), 
        .Q(u_fetch_skid_buffer_q[11]) );
  DFFRX1 u_fetch_skid_buffer_q_reg_7_ ( .D(net2344), .CK(n37801), .RN(n38351), 
        .QN(n50512) );
  DFFRX1 u_fetch_skid_buffer_q_reg_5_ ( .D(net2342), .CK(n37801), .RN(n38350), 
        .Q(u_fetch_skid_buffer_q[5]) );
  DFFRX1 u_fetch_skid_buffer_q_reg_3_ ( .D(net2340), .CK(n37801), .RN(n38321), 
        .Q(u_fetch_skid_buffer_q[3]) );
  DFFRX1 u_decode_pc_q_reg_2_ ( .D(u_decode_N292), .CK(n37799), .RN(n38335), 
        .Q(opcode_pc_w[2]), .QN(n54528) );
  DFFRX1 u_decode_opcode_instr_q_reg_8_ ( .D(u_decode_N744), .CK(n37806), .RN(
        n38320), .Q(opcode_instr_w[8]), .QN(n50665) );
  DFFRX1 u_decode_opcode_instr_q_reg_7_ ( .D(u_decode_N743), .CK(n37806), .RN(
        n38323), .QN(n57095) );
  DFFRX1 u_decode_opcode_instr_q_reg_20_ ( .D(u_decode_N756), .CK(n37802), 
        .RN(n38322), .QN(n50858) );
  DFFRX1 u_muldiv_mult_result_q_reg_10_ ( .D(u_muldiv_result_r[10]), .CK(clk_i), .RN(n38345), .Q(u_muldiv_mult_result_q[10]) );
  DFFRX1 u_muldiv_mult_result_q_reg_11_ ( .D(u_muldiv_result_r[11]), .CK(clk_i), .RN(n38344), .Q(u_muldiv_mult_result_q[11]) );
  DFFRX1 u_muldiv_mult_result_q_reg_12_ ( .D(u_muldiv_result_r[12]), .CK(clk_i), .RN(n38347), .Q(u_muldiv_mult_result_q[12]) );
  DFFRX1 u_fetch_fetch_page_fault_q_reg ( .D(u_fetch_N157), .CK(clk_i), .RN(
        n38349), .Q(u_fetch_fetch_page_fault_q), .QN(n50534) );
  DFFRX1 u_fetch_branch_valid_q_reg ( .D(u_fetch_N15), .CK(clk_i), .RN(n44252), 
        .Q(u_fetch_branch_valid_q), .QN(n50043) );
  DFFRX1 u_muldiv_mult_result_q_reg_13_ ( .D(u_muldiv_result_r[13]), .CK(clk_i), .RN(n38346), .Q(u_muldiv_mult_result_q[13]) );
  DFFRX1 u_fetch_icache_fetch_q_reg ( .D(n8561), .CK(clk_i), .RN(n44252), .Q(
        u_fetch_icache_fetch_q) );
  DFFRX1 u_muldiv_mult_result_q_reg_15_ ( .D(u_muldiv_result_r[15]), .CK(clk_i), .RN(n38345), .Q(u_muldiv_mult_result_q[15]) );
  DFFRX1 u_muldiv_mult_result_q_reg_14_ ( .D(u_muldiv_result_r[14]), .CK(clk_i), .RN(n38344), .Q(u_muldiv_mult_result_q[14]) );
  DFFRX1 u_mmu_state_q_reg_0_ ( .D(n8555), .CK(clk_i), .RN(n38347), .Q(
        u_mmu_state_q[0]), .QN(n57380) );
  DFFRX1 u_mmu_dtlb_req_q_reg ( .D(n8554), .CK(clk_i), .RN(n38356), .Q(
        u_mmu_dtlb_req_q), .QN(n55819) );
  DFFRX1 u_mmu_pte_addr_q_reg_7_ ( .D(U1_U7_Z_7), .CK(n37884), .RN(n38346), 
        .Q(arb_mmu_addr_w[7]) );
  DFFRX1 u_mmu_pte_addr_q_reg_6_ ( .D(U1_U7_Z_6), .CK(n37884), .RN(n38345), 
        .Q(arb_mmu_addr_w[6]) );
  DFFRX1 u_mmu_pte_addr_q_reg_5_ ( .D(U1_U7_Z_5), .CK(n37884), .RN(n38344), 
        .Q(arb_mmu_addr_w[5]) );
  DFFRX1 u_mmu_pte_addr_q_reg_4_ ( .D(U1_U7_Z_4), .CK(n37884), .RN(n38347), 
        .Q(arb_mmu_addr_w[4]) );
  DFFRX1 u_mmu_pte_addr_q_reg_3_ ( .D(U1_U7_Z_3), .CK(n37884), .RN(n38346), 
        .Q(arb_mmu_addr_w[3]) );
  DFFRX1 u_mmu_pte_addr_q_reg_2_ ( .D(U1_U7_Z_2), .CK(n37884), .RN(n38345), 
        .Q(arb_mmu_addr_w[2]) );
  DFFRX1 u_muldiv_mult_result_q_reg_16_ ( .D(u_muldiv_result_r[16]), .CK(clk_i), .RN(n38344), .Q(u_muldiv_mult_result_q[16]) );
  DFFRX1 u_muldiv_mult_result_q_reg_17_ ( .D(u_muldiv_result_r[17]), .CK(clk_i), .RN(n38347), .Q(u_muldiv_mult_result_q[17]) );
  DFFRX1 u_muldiv_mult_result_q_reg_18_ ( .D(u_muldiv_result_r[18]), .CK(clk_i), .RN(n38346), .Q(u_muldiv_mult_result_q[18]) );
  DFFRX1 u_mmu_virt_addr_q_reg_31_ ( .D(n8560), .CK(clk_i), .RN(n38341), .Q(
        u_mmu_virt_addr_q_31) );
  DFFRX1 u_mmu_virt_addr_q_reg_30_ ( .D(n8553), .CK(clk_i), .RN(n38340), .Q(
        u_mmu_virt_addr_q_30) );
  DFFRX1 u_mmu_virt_addr_q_reg_29_ ( .D(n8552), .CK(clk_i), .RN(n38343), .Q(
        u_mmu_virt_addr_q_29) );
  DFFRX1 u_mmu_virt_addr_q_reg_28_ ( .D(n8551), .CK(clk_i), .RN(n38342), .Q(
        u_mmu_virt_addr_q_28) );
  DFFRX1 u_mmu_pte_addr_q_reg_11_ ( .D(U1_U7_Z_11), .CK(n37884), .RN(n44252), 
        .Q(arb_mmu_addr_w[11]) );
  DFFRX1 u_mmu_pte_addr_q_reg_10_ ( .D(U1_U7_Z_10), .CK(n37884), .RN(n44252), 
        .Q(arb_mmu_addr_w[10]) );
  DFFRX1 u_mmu_pte_addr_q_reg_9_ ( .D(U1_U7_Z_9), .CK(n37884), .RN(n38345), 
        .Q(arb_mmu_addr_w[9]) );
  DFFRX1 u_mmu_pte_addr_q_reg_8_ ( .D(U1_U7_Z_8), .CK(n37884), .RN(n38344), 
        .Q(arb_mmu_addr_w[8]) );
  DFFRX1 u_muldiv_mult_result_q_reg_19_ ( .D(u_muldiv_result_r[19]), .CK(clk_i), .RN(n38347), .Q(u_muldiv_mult_result_q[19]) );
  DFFRX1 u_muldiv_mult_result_q_reg_21_ ( .D(u_muldiv_result_r[21]), .CK(clk_i), .RN(n38346), .Q(u_muldiv_mult_result_q[21]) );
  DFFRX1 u_muldiv_mult_result_q_reg_20_ ( .D(u_muldiv_result_r[20]), .CK(clk_i), .RN(n38345), .Q(u_muldiv_mult_result_q[20]) );
  DFFRX1 u_muldiv_mult_result_q_reg_22_ ( .D(u_muldiv_result_r[22]), .CK(clk_i), .RN(n38344), .Q(u_muldiv_mult_result_q[22]) );
  DFFRX1 u_muldiv_mult_result_q_reg_23_ ( .D(u_muldiv_result_r[23]), .CK(clk_i), .RN(n38347), .Q(u_muldiv_mult_result_q[23]) );
  DFFRX1 u_exec_result_q_reg_26_ ( .D(u_exec_alu_p_w[26]), .CK(clk_i), .RN(
        n38338), .Q(n37406) );
  DFFRX1 u_decode_u_regfile_reg_r21_q_reg_30_ ( .D(u_decode_u_regfile_N870), 
        .CK(n37810), .RN(n38341), .Q(n2981) );
  DFFRX1 u_decode_u_regfile_reg_r21_q_reg_26_ ( .D(u_decode_u_regfile_N866), 
        .CK(n37810), .RN(n38337), .Q(n2646), .QN(n46032) );
  DFFRX1 u_decode_u_regfile_reg_r21_q_reg_29_ ( .D(u_decode_u_regfile_N869), 
        .CK(n37810), .RN(n38318), .Q(n3010), .QN(n45466) );
  DFFRX1 u_decode_u_regfile_reg_r20_q_reg_29_ ( .D(u_decode_u_regfile_N832), 
        .CK(n37811), .RN(n38317), .Q(n3009), .QN(n45483) );
  DFFRX1 u_decode_u_regfile_reg_r18_q_reg_30_ ( .D(u_decode_u_regfile_N759), 
        .CK(n37813), .RN(n38340), .Q(n2978), .QN(n45631) );
  DFFRX1 u_decode_u_regfile_reg_r27_q_reg_1_ ( .D(u_decode_u_regfile_N1063), 
        .CK(n37863), .RN(n38336), .Q(n1977), .QN(n48213) );
  DFFRX1 u_decode_u_regfile_reg_r11_q_reg_1_ ( .D(u_decode_u_regfile_N471), 
        .CK(n37851), .RN(n38335), .QN(n48161) );
  DFFRX1 u_muldiv_mult_result_q_reg_2_ ( .D(u_muldiv_result_r[2]), .CK(clk_i), 
        .RN(n38346), .QN(n1889) );
  DFFRX1 u_fetch_fetch_pc_q_reg_1_ ( .D(mem_i_pc_o[1]), .CK(n37882), .RN(
        n38343), .QN(n1759) );
  DFFRX1 u_fetch_fetch_pc_q_reg_0_ ( .D(mem_i_pc_o[0]), .CK(n37882), .RN(
        n38345), .QN(n1758) );
  DFFRX1 u_fetch_skid_valid_q_reg ( .D(n43319), .CK(clk_i), .RN(n38321), .Q(
        n58511), .QN(n8801) );
  DFFRX1 u_fetch_fetch_pc_q_reg_2_ ( .D(n36343), .CK(n37882), .RN(n38338), 
        .QN(n1760) );
  DFFRX1 u_decode_opcode_instr_q_reg_21_ ( .D(u_decode_N757), .CK(n37802), 
        .RN(n38320), .Q(n43012), .QN(n37342) );
  DFFRX1 u_fetch_fetch_pc_q_reg_3_ ( .D(u_fetch_N52), .CK(n37882), .RN(n38337), 
        .QN(n1761) );
  DFFRX1 u_mmu_virt_addr_q_reg_26_ ( .D(u_mmu_request_addr_w[26]), .CK(n37803), 
        .RN(n38316), .Q(n57389) );
  DFFRX1 u_mmu_virt_addr_q_reg_22_ ( .D(u_mmu_request_addr_w[22]), .CK(n37803), 
        .RN(n38342), .Q(n57388) );
  DFFRX1 u_mmu_virt_addr_q_reg_27_ ( .D(u_mmu_request_addr_w[27]), .CK(n37803), 
        .RN(n38341), .Q(n57390) );
  DFFRX1 u_mmu_virt_addr_q_reg_25_ ( .D(u_mmu_request_addr_w[25]), .CK(n37803), 
        .RN(n38340), .Q(n57391) );
  DFFRX1 u_mmu_virt_addr_q_reg_23_ ( .D(u_mmu_request_addr_w[23]), .CK(n37803), 
        .RN(n38343), .Q(n57387) );
  DFFRX1 u_mmu_virt_addr_q_reg_24_ ( .D(u_mmu_request_addr_w[24]), .CK(n37803), 
        .RN(n38342), .Q(n57386) );
  DFFRX1 u_fetch_fetch_pc_q_reg_4_ ( .D(u_fetch_N53), .CK(n37882), .RN(n38336), 
        .QN(n1762) );
  DFFRX1 u_fetch_skid_buffer_q_reg_27_ ( .D(net2370), .CK(n37798), .RN(n38352), 
        .QN(n1836) );
  DFFRX1 u_fetch_skid_buffer_q_reg_58_ ( .D(net2411), .CK(n37797), .RN(n38335), 
        .QN(n2190) );
  DFFRX1 u_fetch_skid_buffer_q_reg_42_ ( .D(net2390), .CK(n37796), .RN(n38362), 
        .QN(n2143) );
  DFFRX1 u_fetch_skid_buffer_q_reg_41_ ( .D(net2389), .CK(n37796), .RN(n38361), 
        .QN(n2140) );
  DFFRX1 u_fetch_skid_buffer_q_reg_39_ ( .D(net2387), .CK(n37796), .RN(n38338), 
        .QN(n2134) );
  DFFRX1 u_fetch_skid_buffer_q_reg_38_ ( .D(net2386), .CK(n37796), .RN(n38337), 
        .QN(n2131) );
  DFFRX1 u_fetch_skid_buffer_q_reg_37_ ( .D(net2385), .CK(n37796), .RN(n38336), 
        .QN(n2099) );
  DFFRX1 u_fetch_skid_buffer_q_reg_36_ ( .D(net2384), .CK(n37796), .RN(n38335), 
        .QN(n2067) );
  DFFRX1 u_fetch_skid_buffer_q_reg_34_ ( .D(net2382), .CK(n37796), .RN(n38338), 
        .QN(n2005) );
  DFFRX1 u_decode_opcode_instr_q_reg_32_ ( .D(u_decode_N768), .CK(n37807), 
        .RN(n38351), .Q(n50611), .QN(n17098) );
  DFFRX1 u_fetch_skid_buffer_q_reg_63_ ( .D(net2416), .CK(n37797), .RN(n38341), 
        .QN(n1930) );
  DFFRX1 u_fetch_skid_buffer_q_reg_62_ ( .D(net2415), .CK(n37797), .RN(n38340), 
        .QN(n1929) );
  DFFRX1 u_fetch_skid_buffer_q_reg_61_ ( .D(net2414), .CK(n37797), .RN(n38315), 
        .QN(n1935) );
  DFFRX1 u_fetch_skid_buffer_q_reg_60_ ( .D(net2413), .CK(n37797), .RN(n38318), 
        .QN(n1937) );
  DFFRX1 u_fetch_skid_buffer_q_reg_59_ ( .D(net2412), .CK(n37797), .RN(n38317), 
        .QN(n1939) );
  DFFRX1 u_fetch_skid_buffer_q_reg_57_ ( .D(net2410), .CK(n37797), .RN(n38343), 
        .QN(n2187) );
  DFFRX1 u_fetch_skid_buffer_q_reg_56_ ( .D(net2409), .CK(n37797), .RN(n38342), 
        .QN(n2184) );
  DFFRX1 u_fetch_skid_buffer_q_reg_55_ ( .D(net2408), .CK(n37797), .RN(n38360), 
        .QN(n2181) );
  DFFRX1 u_fetch_skid_buffer_q_reg_54_ ( .D(net2407), .CK(n37797), .RN(n38359), 
        .QN(n2178) );
  DFFRX1 u_fetch_skid_buffer_q_reg_53_ ( .D(net2406), .CK(n37797), .RN(n38362), 
        .QN(n2175) );
  DFFRX1 u_fetch_skid_buffer_q_reg_52_ ( .D(net2405), .CK(n37797), .RN(n38361), 
        .QN(n2172) );
  DFFRX1 u_fetch_skid_buffer_q_reg_51_ ( .D(net2404), .CK(n37797), .RN(n38360), 
        .QN(n2169) );
  DFFRX1 u_fetch_skid_buffer_q_reg_50_ ( .D(net2403), .CK(n37797), .RN(n38359), 
        .QN(n2166) );
  DFFRX1 u_fetch_skid_buffer_q_reg_49_ ( .D(net2402), .CK(n37797), .RN(n38362), 
        .QN(n2163) );
  DFFRX1 u_fetch_skid_buffer_q_reg_48_ ( .D(net2401), .CK(n37797), .RN(n38361), 
        .QN(n2160) );
  DFFRX1 u_fetch_skid_buffer_q_reg_47_ ( .D(net2395), .CK(n37796), .RN(n38360), 
        .QN(n2156) );
  DFFRX1 u_fetch_skid_buffer_q_reg_46_ ( .D(net2394), .CK(n37796), .RN(n38359), 
        .QN(n2152) );
  DFFRX1 u_fetch_skid_buffer_q_reg_45_ ( .D(net2393), .CK(n37796), .RN(n38362), 
        .QN(n2149) );
  DFFRX1 u_fetch_skid_buffer_q_reg_44_ ( .D(net2392), .CK(n37796), .RN(n38361), 
        .QN(n2146) );
  DFFRX1 u_fetch_skid_buffer_q_reg_43_ ( .D(net2391), .CK(n37796), .RN(n38360), 
        .QN(n1932) );
  DFFRX1 u_fetch_skid_buffer_q_reg_40_ ( .D(net2388), .CK(n37796), .RN(n38341), 
        .QN(n2137) );
  DFFRX1 u_fetch_skid_buffer_q_reg_35_ ( .D(net2383), .CK(n37796), .RN(n38340), 
        .QN(n2036) );
  DFFRX1 u_fetch_skid_buffer_q_reg_33_ ( .D(net2381), .CK(n37796), .RN(n38343), 
        .QN(n1973) );
  DFFRX1 u_fetch_skid_buffer_q_reg_32_ ( .D(net2380), .CK(n37796), .RN(n38344), 
        .QN(n1941) );
  DFFRX1 u_fetch_fetch_pc_q_reg_5_ ( .D(u_fetch_N54), .CK(n37882), .RN(n38337), 
        .QN(n1763) );
  DFFRX1 u_fetch_fetch_pc_q_reg_6_ ( .D(u_fetch_N55), .CK(n37882), .RN(n38336), 
        .QN(n1764) );
  DFFRX1 u_fetch_fetch_pc_q_reg_7_ ( .D(u_fetch_N56), .CK(n37882), .RN(n38335), 
        .QN(n1765) );
  DFFRX1 u_fetch_fetch_pc_q_reg_8_ ( .D(u_fetch_N57), .CK(n37882), .RN(n38359), 
        .QN(n1766) );
  DFFRX1 u_fetch_fetch_pc_q_reg_9_ ( .D(u_fetch_N58), .CK(n37882), .RN(n38362), 
        .QN(n1767) );
  DFFRX1 u_fetch_fetch_pc_q_reg_10_ ( .D(u_fetch_N59), .CK(n37882), .RN(n38361), .QN(n1768) );
  DFFRX1 u_fetch_fetch_pc_q_reg_11_ ( .D(u_fetch_N60), .CK(n37882), .RN(n38360), .QN(n1769) );
  DFFRX1 u_mmu_mem_req_q_reg ( .D(n8559), .CK(clk_i), .RN(n44252), .Q(n58183)
         );
  DFFRX1 u_fetch_fetch_pc_q_reg_12_ ( .D(u_fetch_N61), .CK(n37882), .RN(n38359), .QN(n1770) );
  DFFRX1 u_fetch_fetch_pc_q_reg_13_ ( .D(u_fetch_N62), .CK(n37882), .RN(n38362), .QN(n1771) );
  DFFRX1 u_fetch_fetch_pc_q_reg_14_ ( .D(u_fetch_N63), .CK(n37882), .RN(n38361), .QN(n1772) );
  DFFRX1 u_fetch_branch_pc_q_reg_26_ ( .D(net2312), .CK(n37866), .RN(n38316), 
        .QN(n2189) );
  DFFRX1 u_fetch_branch_pc_q_reg_25_ ( .D(net2311), .CK(n37866), .RN(n38342), 
        .QN(n2186) );
  DFFRX1 u_fetch_branch_pc_q_reg_0_ ( .D(net2281), .CK(n37867), .RN(n38347), 
        .QN(n1940) );
  DFFRX1 u_fetch_branch_pc_q_reg_30_ ( .D(net2316), .CK(n37866), .RN(n38341), 
        .QN(n2221) );
  DFFRX1 u_fetch_branch_pc_q_reg_29_ ( .D(net2315), .CK(n37866), .RN(n38315), 
        .QN(n1934) );
  DFFRX1 u_decode_inst_q_reg_28_ ( .D(n8517), .CK(clk_i), .RN(n38350), .Q(
        opcode_opcode_w[28]), .QN(n58457) );
  DFFRX1 u_decode_inst_q_reg_29_ ( .D(n8518), .CK(clk_i), .RN(n38349), .Q(
        opcode_opcode_w[29]), .QN(n73367) );
  DFFRX1 u_decode_opcode_instr_q_reg_10_ ( .D(u_decode_N746), .CK(n37806), 
        .RN(n38323), .Q(opcode_instr_w[10]), .QN(n40919) );
  DFFRX1 u_decode_opcode_instr_q_reg_18_ ( .D(u_decode_N754), .CK(n37802), 
        .RN(n38322), .Q(opcode_instr_w_18), .QN(n40931) );
  DFFRX1 u_decode_opcode_instr_q_reg_4_ ( .D(u_decode_N740), .CK(n37806), .RN(
        n38321), .Q(n1851), .QN(n40934) );
  DFFRX1 u_decode_opcode_instr_q_reg_26_ ( .D(u_decode_N762), .CK(n37802), 
        .RN(n38352), .Q(opcode_instr_w_26), .QN(n45704) );
  DFFRX1 u_decode_opcode_instr_q_reg_19_ ( .D(u_decode_N755), .CK(n37802), 
        .RN(n38320), .Q(n40917), .QN(n8955) );
  DFFRX1 u_decode_pc_q_reg_19_ ( .D(u_decode_N309), .CK(n37800), .RN(n38360), 
        .Q(opcode_pc_w[19]), .QN(n58338) );
  DFFRX1 u_decode_pc_q_reg_6_ ( .D(u_decode_N296), .CK(n37799), .RN(n38338), 
        .Q(opcode_pc_w[6]), .QN(n58431) );
  DFFRX1 u_decode_pc_q_reg_5_ ( .D(u_decode_N295), .CK(n37799), .RN(n38337), 
        .Q(opcode_pc_w[5]), .QN(n58426) );
  DFFRX1 u_decode_opcode_instr_q_reg_22_ ( .D(u_decode_N758), .CK(n37802), 
        .RN(n38323), .Q(n40930) );
  DFFRX1 u_exec_rd_x_q_reg_4_ ( .D(u_exec_N242), .CK(clk_i), .RN(n73547), .Q(
        writeback_exec_idx_w[4]), .QN(n50838) );
  DFFRHQX1 u_muldiv_mult_result_q_reg_30_ ( .D(u_muldiv_result_r[30]), .CK(
        clk_i), .RN(n73547), .Q(u_muldiv_mult_result_q[30]) );
  DFFRX1 u_exec_rd_x_q_reg_2_ ( .D(u_exec_N240), .CK(clk_i), .RN(n73547), .Q(
        writeback_exec_idx_w[2]), .QN(n50802) );
  DFFRX1 u_muldiv_mult_result_q_reg_31_ ( .D(u_muldiv_result_r[31]), .CK(clk_i), .RN(n73547), .Q(n38972) );
  AND2X1 U37134 ( .A(n61404), .B(n61403), .Y(n36346) );
  NOR2X1 U37135 ( .A(n36348), .B(n36349), .Y(n36347) );
  INVX1 U37136 ( .A(n36347), .Y(n61736) );
  AND2X1 U37137 ( .A(n61762), .B(n61734), .Y(n36348) );
  AND2X1 U37138 ( .A(n42042), .B(n61735), .Y(n36349) );
  NOR2X1 U37139 ( .A(n36351), .B(n36352), .Y(n36350) );
  INVX1 U37140 ( .A(n36350), .Y(n62777) );
  AND2X1 U37141 ( .A(n62775), .B(n70799), .Y(n36351) );
  AND2X1 U37142 ( .A(n42109), .B(n62776), .Y(n36352) );
  NOR2X1 U37143 ( .A(n36354), .B(n36355), .Y(n36353) );
  INVX1 U37144 ( .A(n36353), .Y(n62780) );
  AND2X1 U37145 ( .A(n62778), .B(n62777), .Y(n36354) );
  AND2X1 U37146 ( .A(n42115), .B(n62779), .Y(n36355) );
  AND2X1 U37147 ( .A(n63071), .B(n63070), .Y(n36356) );
  AND2X1 U37148 ( .A(n63955), .B(n63954), .Y(n36357) );
  NOR2X1 U37149 ( .A(n36359), .B(n36360), .Y(n36358) );
  INVX1 U37150 ( .A(n36358), .Y(n65941) );
  AND2X1 U37151 ( .A(n62701), .B(n62700), .Y(n36359) );
  AND2X1 U37152 ( .A(n41950), .B(n62702), .Y(n36360) );
  NOR2X1 U37153 ( .A(n40292), .B(n40293), .Y(n36361) );
  XNOR2X1 U37154 ( .A(n66904), .B(n66903), .Y(n36362) );
  XOR2X1 U37155 ( .A(n40087), .B(n36363), .Y(n68536) );
  XOR2X1 U37156 ( .A(n43708), .B(n37955), .Y(n36363) );
  OR2X1 U37157 ( .A(n62090), .B(n62158), .Y(n62091) );
  NOR2X1 U37158 ( .A(n36365), .B(n36366), .Y(n36364) );
  INVX1 U37159 ( .A(n36364), .Y(n62298) );
  AND2X1 U37160 ( .A(n62600), .B(n62295), .Y(n36365) );
  AND2X1 U37161 ( .A(n42055), .B(n62297), .Y(n36366) );
  NOR2X1 U37162 ( .A(n36368), .B(n36369), .Y(n36367) );
  INVX1 U37163 ( .A(n36367), .Y(n62301) );
  AND2X1 U37164 ( .A(n62598), .B(n62298), .Y(n36368) );
  AND2X1 U37165 ( .A(n42066), .B(n62300), .Y(n36369) );
  NOR2X1 U37166 ( .A(n36371), .B(n36372), .Y(n36370) );
  INVX1 U37167 ( .A(n36370), .Y(n61849) );
  AND2X1 U37168 ( .A(n61997), .B(n61845), .Y(n36371) );
  AND2X1 U37169 ( .A(n41875), .B(n61847), .Y(n36372) );
  OR2X1 U37170 ( .A(n36373), .B(n36374), .Y(n62324) );
  INVX1 U37171 ( .A(n42118), .Y(n36373) );
  AND2X1 U37172 ( .A(n38419), .B(n62323), .Y(n36374) );
  OR2X1 U37173 ( .A(n36375), .B(n36376), .Y(n40174) );
  INVX1 U37174 ( .A(n67919), .Y(n36375) );
  NAND2X1 U37175 ( .A(n67920), .B(n68544), .Y(n36376) );
  OR2X1 U37176 ( .A(n38430), .B(n38431), .Y(n36377) );
  NOR2X1 U37177 ( .A(n36379), .B(n36380), .Y(n36378) );
  INVX1 U37178 ( .A(n36378), .Y(n62295) );
  AND2X1 U37179 ( .A(n62292), .B(n62293), .Y(n36379) );
  AND2X1 U37180 ( .A(n42041), .B(n62294), .Y(n36380) );
  XNOR2X1 U37181 ( .A(n66928), .B(n66894), .Y(n36381) );
  AND2X1 U37182 ( .A(n61905), .B(n61904), .Y(n36382) );
  OR2X1 U37183 ( .A(n36383), .B(n36384), .Y(n65568) );
  AND2X1 U37184 ( .A(n64903), .B(n43711), .Y(n36383) );
  NOR2X1 U37185 ( .A(n39143), .B(n39144), .Y(n36384) );
  NOR2X1 U37186 ( .A(n36386), .B(n36387), .Y(n36385) );
  INVX1 U37187 ( .A(n36385), .Y(n62220) );
  AND2X1 U37188 ( .A(n62647), .B(n62216), .Y(n36386) );
  AND2X1 U37189 ( .A(n41872), .B(n62218), .Y(n36387) );
  AND2X1 U37190 ( .A(n62013), .B(n62012), .Y(n36388) );
  NOR2X1 U37191 ( .A(n36390), .B(n36391), .Y(n36389) );
  INVX1 U37192 ( .A(n36389), .Y(n62216) );
  AND2X1 U37193 ( .A(n62213), .B(n62214), .Y(n36390) );
  AND2X1 U37194 ( .A(n41860), .B(n62215), .Y(n36391) );
  XOR2X1 U37195 ( .A(n36402), .B(n67903), .Y(n36392) );
  AND2X1 U37196 ( .A(n38024), .B(n38025), .Y(n36393) );
  AND2X1 U37197 ( .A(n61411), .B(n61410), .Y(n36394) );
  AND2X1 U37198 ( .A(n61562), .B(n61561), .Y(n36395) );
  AND2X1 U37199 ( .A(n61925), .B(n61924), .Y(n36396) );
  AND2X1 U37200 ( .A(n61503), .B(n61502), .Y(n36397) );
  NOR2X1 U37201 ( .A(n36399), .B(n36400), .Y(n36398) );
  INVX1 U37202 ( .A(n36398), .Y(n62054) );
  AND2X1 U37203 ( .A(n62182), .B(n62051), .Y(n36399) );
  NOR2X1 U37204 ( .A(n38589), .B(n38590), .Y(n36400) );
  XNOR2X1 U37205 ( .A(n38491), .B(n36401), .Y(n65511) );
  XOR2X1 U37206 ( .A(n65480), .B(n65153), .Y(n36401) );
  OR2X1 U37207 ( .A(n67614), .B(n67615), .Y(n36402) );
  NOR2X1 U37208 ( .A(n65985), .B(n36403), .Y(n39840) );
  NAND2X1 U37209 ( .A(n65984), .B(n65986), .Y(n36403) );
  XNOR2X1 U37210 ( .A(n36404), .B(n66501), .Y(n41366) );
  INVX1 U37211 ( .A(n66622), .Y(n36404) );
  OR2X1 U37212 ( .A(n36411), .B(n38606), .Y(n36405) );
  NAND2X1 U37213 ( .A(n36406), .B(n61449), .Y(n61423) );
  NOR2X1 U37214 ( .A(n40231), .B(n40232), .Y(n36406) );
  OR2X1 U37215 ( .A(n63054), .B(n36407), .Y(n63056) );
  INVX1 U37216 ( .A(n63055), .Y(n36407) );
  AND2X1 U37217 ( .A(n36409), .B(n36408), .Y(n67254) );
  INVX1 U37218 ( .A(n41110), .Y(n36408) );
  NAND2X1 U37219 ( .A(n67248), .B(n40090), .Y(n36409) );
  NOR2X1 U37220 ( .A(n43698), .B(n66918), .Y(n36410) );
  OR2X1 U37221 ( .A(n36411), .B(n38606), .Y(n67563) );
  AND2X1 U37222 ( .A(n66620), .B(n43540), .Y(n36411) );
  OR2X1 U37223 ( .A(n70187), .B(n36412), .Y(n69229) );
  INVX1 U37224 ( .A(n43697), .Y(n36412) );
  NOR2X1 U37225 ( .A(n36414), .B(n36415), .Y(n36413) );
  INVX1 U37226 ( .A(n36413), .Y(n61712) );
  AND2X1 U37227 ( .A(n61709), .B(n61710), .Y(n36414) );
  AND2X1 U37228 ( .A(n41963), .B(n61711), .Y(n36415) );
  AND2X1 U37229 ( .A(n61715), .B(n61714), .Y(n36416) );
  XNOR2X1 U37230 ( .A(n60720), .B(n60721), .Y(n38290) );
  XOR2X1 U37231 ( .A(n69215), .B(n36752), .Y(n69216) );
  OR2X1 U37232 ( .A(n39099), .B(n39100), .Y(n36417) );
  AND2X1 U37233 ( .A(n61720), .B(n61719), .Y(n36418) );
  OR2X1 U37234 ( .A(n40667), .B(n40668), .Y(n36419) );
  OR2X1 U37235 ( .A(n36420), .B(n61296), .Y(n61293) );
  INVX1 U37236 ( .A(n61292), .Y(n36420) );
  AND2X1 U37237 ( .A(n63732), .B(n63733), .Y(n40752) );
  OR2X1 U37238 ( .A(n66616), .B(n36421), .Y(n66618) );
  INVX1 U37239 ( .A(n43559), .Y(n36421) );
  XNOR2X1 U37240 ( .A(n36422), .B(n65619), .Y(n65531) );
  INVX1 U37241 ( .A(n65625), .Y(n36422) );
  XOR2X1 U37242 ( .A(n36423), .B(n69565), .Y(n69570) );
  OR2X1 U37243 ( .A(n40400), .B(n38062), .Y(n36423) );
  AND2X1 U37244 ( .A(n66294), .B(n67179), .Y(n36424) );
  XNOR2X1 U37245 ( .A(n67217), .B(n67218), .Y(n36425) );
  NOR2X1 U37246 ( .A(n43636), .B(n67219), .Y(n36426) );
  OR2X1 U37247 ( .A(n40348), .B(n40349), .Y(n36427) );
  OR2X1 U37248 ( .A(n40348), .B(n40349), .Y(n36428) );
  XNOR2X1 U37249 ( .A(n36430), .B(n36429), .Y(n61084) );
  INVX1 U37250 ( .A(n39042), .Y(n36429) );
  XOR2X1 U37251 ( .A(n60888), .B(n60886), .Y(n36430) );
  OR2X1 U37252 ( .A(n36431), .B(n36432), .Y(n68886) );
  INVX1 U37253 ( .A(n43653), .Y(n36431) );
  AND2X1 U37254 ( .A(n67945), .B(n67946), .Y(n36432) );
  AND2X1 U37255 ( .A(n38061), .B(n39226), .Y(n36433) );
  INVX1 U37256 ( .A(n36433), .Y(n69553) );
  XNOR2X1 U37257 ( .A(n69224), .B(n69223), .Y(n36434) );
  XOR2X1 U37258 ( .A(n40020), .B(n36435), .Y(n69910) );
  XOR2X1 U37259 ( .A(n69914), .B(n43707), .Y(n36435) );
  XOR2X1 U37260 ( .A(n69904), .B(n69905), .Y(n36436) );
  NOR2X1 U37261 ( .A(n36438), .B(n36439), .Y(n36437) );
  INVX1 U37262 ( .A(n36437), .Y(n59667) );
  AND2X1 U37263 ( .A(n59381), .B(n59451), .Y(n36438) );
  AND2X1 U37264 ( .A(n41495), .B(n59384), .Y(n36439) );
  AND2X1 U37265 ( .A(n61892), .B(n61891), .Y(n36440) );
  OR2X1 U37266 ( .A(n64577), .B(n36441), .Y(n65590) );
  INVX1 U37267 ( .A(n43508), .Y(n36441) );
  XOR2X1 U37268 ( .A(n41750), .B(n59265), .Y(n36442) );
  XOR2X1 U37269 ( .A(n38396), .B(n38472), .Y(n36443) );
  INVX1 U37270 ( .A(n68831), .Y(n36444) );
  XNOR2X1 U37271 ( .A(n41139), .B(n68520), .Y(n36445) );
  AND2X1 U37272 ( .A(n60166), .B(n36446), .Y(n39494) );
  NOR2X1 U37273 ( .A(n40547), .B(n40548), .Y(n36446) );
  OR2X1 U37274 ( .A(n36447), .B(n36448), .Y(n47700) );
  OR2X1 U37275 ( .A(n47663), .B(n47662), .Y(n36447) );
  OR2X1 U37276 ( .A(n47684), .B(n47683), .Y(n36448) );
  OR2X1 U37277 ( .A(n36449), .B(n36450), .Y(n42352) );
  OR2X1 U37278 ( .A(n36481), .B(n46586), .Y(n36449) );
  OR2X1 U37279 ( .A(n36470), .B(n46587), .Y(n36450) );
  NAND2X1 U37280 ( .A(n46396), .B(n36451), .Y(n40290) );
  NOR2X1 U37281 ( .A(n36452), .B(n46397), .Y(n36451) );
  AND2X1 U37282 ( .A(n46395), .B(n1825), .Y(n36452) );
  OR2X1 U37283 ( .A(n36453), .B(n69226), .Y(n68544) );
  INVX1 U37284 ( .A(n43691), .Y(n36453) );
  AND2X1 U37285 ( .A(n62835), .B(n62834), .Y(n36454) );
  XOR2X1 U37286 ( .A(n61059), .B(n61123), .Y(n36455) );
  OR2X1 U37287 ( .A(n60863), .B(n61313), .Y(n60864) );
  OR2X1 U37288 ( .A(n37948), .B(n37949), .Y(n36456) );
  OR2X1 U37289 ( .A(n62824), .B(n62823), .Y(n62826) );
  INVX1 U37290 ( .A(n63722), .Y(n36457) );
  OR2X1 U37291 ( .A(n36458), .B(n36459), .Y(n63987) );
  INVX1 U37292 ( .A(n63719), .Y(n36458) );
  NAND2X1 U37293 ( .A(n36457), .B(n63718), .Y(n36459) );
  AND2X1 U37294 ( .A(n60521), .B(n60520), .Y(n36460) );
  NOR2X1 U37295 ( .A(n36462), .B(n36463), .Y(n36461) );
  INVX1 U37296 ( .A(n36461), .Y(n60858) );
  AND2X1 U37297 ( .A(n61318), .B(n60855), .Y(n36462) );
  AND2X1 U37298 ( .A(n41943), .B(n60857), .Y(n36463) );
  NOR2X1 U37299 ( .A(n70187), .B(n69231), .Y(n36464) );
  AND2X1 U37300 ( .A(n36465), .B(n67590), .Y(n67593) );
  INVX1 U37301 ( .A(n43507), .Y(n36465) );
  OR2X1 U37302 ( .A(n36466), .B(n38285), .Y(n64599) );
  INVX1 U37303 ( .A(n64596), .Y(n36466) );
  OR2X1 U37304 ( .A(n36467), .B(n36468), .Y(n64303) );
  AND2X1 U37305 ( .A(n64302), .B(n64301), .Y(n36467) );
  AND2X1 U37306 ( .A(n64298), .B(n64297), .Y(n36468) );
  OR2X1 U37307 ( .A(n36469), .B(n62340), .Y(n62341) );
  OR2X1 U37308 ( .A(n39088), .B(n39089), .Y(n36469) );
  INVX1 U37309 ( .A(n38690), .Y(n36470) );
  OR2X1 U37310 ( .A(n36471), .B(n66588), .Y(n66593) );
  INVX1 U37311 ( .A(n40142), .Y(n36471) );
  XNOR2X1 U37312 ( .A(n41058), .B(n67228), .Y(n36472) );
  XNOR2X1 U37313 ( .A(n41578), .B(n64869), .Y(n36473) );
  XOR2X1 U37314 ( .A(n39018), .B(n36474), .Y(n65965) );
  XOR2X1 U37315 ( .A(n66534), .B(n43643), .Y(n36474) );
  INVX1 U37316 ( .A(n61747), .Y(n36475) );
  AND2X1 U37317 ( .A(n36476), .B(n61746), .Y(n39086) );
  NOR2X1 U37318 ( .A(n36475), .B(n61751), .Y(n36476) );
  OR2X1 U37319 ( .A(n39398), .B(n39399), .Y(n36477) );
  NOR2X1 U37320 ( .A(n36479), .B(n36480), .Y(n36478) );
  INVX1 U37321 ( .A(n36478), .Y(n60069) );
  AND2X1 U37322 ( .A(n60060), .B(n60059), .Y(n36479) );
  AND2X1 U37323 ( .A(n60079), .B(n60081), .Y(n36480) );
  AND2X1 U37324 ( .A(n2508), .B(n40521), .Y(n36481) );
  INVX1 U37325 ( .A(n42370), .Y(n36482) );
  AND2X1 U37326 ( .A(n60411), .B(n60410), .Y(n36483) );
  OR2X1 U37327 ( .A(n59856), .B(n36484), .Y(n59858) );
  INVX1 U37328 ( .A(n59857), .Y(n36484) );
  OR2X1 U37329 ( .A(n36485), .B(n36486), .Y(n63898) );
  INVX1 U37330 ( .A(n41992), .Y(n36485) );
  NOR2X1 U37331 ( .A(n38099), .B(n39158), .Y(n36486) );
  AND2X1 U37332 ( .A(n63897), .B(n63898), .Y(n36487) );
  OR2X1 U37333 ( .A(n40369), .B(n40370), .Y(n36488) );
  NAND2X1 U37334 ( .A(n59954), .B(n59953), .Y(n36489) );
  NOR2X1 U37335 ( .A(n36491), .B(n36492), .Y(n36490) );
  INVX1 U37336 ( .A(n36490), .Y(n60154) );
  AND2X1 U37337 ( .A(n36749), .B(n60149), .Y(n36491) );
  AND2X1 U37338 ( .A(n60151), .B(n60150), .Y(n36492) );
  AND2X1 U37339 ( .A(n60156), .B(n60155), .Y(n36493) );
  OR2X1 U37340 ( .A(n36494), .B(n36495), .Y(n61110) );
  OR2X1 U37341 ( .A(n60572), .B(n41337), .Y(n36494) );
  AND2X1 U37342 ( .A(n60895), .B(n60573), .Y(n36495) );
  OR2X1 U37343 ( .A(n39539), .B(n36496), .Y(n62529) );
  NAND2X1 U37344 ( .A(n39416), .B(n62528), .Y(n36496) );
  NOR2X1 U37345 ( .A(n38646), .B(n36497), .Y(n41613) );
  OR2X1 U37346 ( .A(n38647), .B(n36498), .Y(n36497) );
  INVX1 U37347 ( .A(n61102), .Y(n36498) );
  OR2X1 U37348 ( .A(n42353), .B(n42354), .Y(n36499) );
  OR2X1 U37349 ( .A(n59853), .B(n59665), .Y(n59666) );
  NAND2X1 U37350 ( .A(n67259), .B(n36503), .Y(n36500) );
  NAND2X1 U37351 ( .A(n36500), .B(n36501), .Y(n41096) );
  OR2X1 U37352 ( .A(n36502), .B(n67258), .Y(n36501) );
  INVX1 U37353 ( .A(n67261), .Y(n36502) );
  AND2X1 U37354 ( .A(n67260), .B(n67261), .Y(n36503) );
  OR2X1 U37355 ( .A(n60727), .B(n36504), .Y(n60732) );
  INVX1 U37356 ( .A(n60730), .Y(n36504) );
  AND2X1 U37357 ( .A(n36505), .B(n36506), .Y(n67234) );
  OR2X1 U37358 ( .A(n41110), .B(n67248), .Y(n36505) );
  AND2X1 U37359 ( .A(n67233), .B(n67249), .Y(n36506) );
  NOR2X1 U37360 ( .A(n66922), .B(n36508), .Y(n36507) );
  INVX1 U37361 ( .A(n36507), .Y(n67591) );
  INVX1 U37362 ( .A(n43513), .Y(n36508) );
  OR2X1 U37363 ( .A(n67247), .B(n36509), .Y(n67233) );
  INVX1 U37364 ( .A(n43684), .Y(n36509) );
  INVX1 U37365 ( .A(n39091), .Y(n36510) );
  OR2X1 U37366 ( .A(n36511), .B(n69219), .Y(n69222) );
  NAND2X1 U37367 ( .A(n36510), .B(n69221), .Y(n36511) );
  AND2X1 U37368 ( .A(n60555), .B(n60554), .Y(n36512) );
  OR2X1 U37369 ( .A(n39667), .B(n39668), .Y(n36513) );
  OR2X1 U37370 ( .A(n36514), .B(n36515), .Y(n65237) );
  OR2X1 U37371 ( .A(n65231), .B(n65230), .Y(n36514) );
  OR2X1 U37372 ( .A(n65236), .B(n65235), .Y(n36515) );
  NAND2X1 U37373 ( .A(n67920), .B(n69225), .Y(n36516) );
  OR2X1 U37374 ( .A(n38874), .B(n38875), .Y(n36517) );
  XOR2X1 U37375 ( .A(n69564), .B(n36518), .Y(n69572) );
  NAND2X1 U37376 ( .A(n70185), .B(n38006), .Y(n36518) );
  OR2X1 U37377 ( .A(n36519), .B(n36520), .Y(n64651) );
  INVX1 U37378 ( .A(n64650), .Y(n36519) );
  AND2X1 U37379 ( .A(n64311), .B(n40198), .Y(n36520) );
  OR2X1 U37380 ( .A(n36521), .B(n36522), .Y(n69571) );
  OR2X1 U37381 ( .A(n69239), .B(n41180), .Y(n36521) );
  NOR2X1 U37382 ( .A(n40087), .B(n41410), .Y(n36522) );
  XOR2X1 U37383 ( .A(n39973), .B(n68522), .Y(n36523) );
  OR2X1 U37384 ( .A(n38530), .B(n38531), .Y(n36524) );
  INVX1 U37385 ( .A(n36524), .Y(n38529) );
  AND2X1 U37386 ( .A(n65266), .B(n65265), .Y(n36525) );
  OR2X1 U37387 ( .A(n36526), .B(n61098), .Y(n62354) );
  AND2X1 U37388 ( .A(n61090), .B(n61089), .Y(n36526) );
  OR2X1 U37389 ( .A(n39593), .B(n39594), .Y(n36527) );
  OR2X1 U37390 ( .A(n36528), .B(n36529), .Y(n63453) );
  AND2X1 U37391 ( .A(n63381), .B(n63380), .Y(n36528) );
  OR2X1 U37392 ( .A(n63379), .B(n39536), .Y(n36529) );
  OR2X1 U37393 ( .A(n39569), .B(n36530), .Y(n60710) );
  INVX1 U37394 ( .A(n60711), .Y(n36530) );
  AND2X1 U37395 ( .A(n64328), .B(n64327), .Y(n36531) );
  INVX1 U37396 ( .A(n36531), .Y(n64330) );
  OR2X1 U37397 ( .A(n36532), .B(n36533), .Y(n62535) );
  AND2X1 U37398 ( .A(n61294), .B(n61293), .Y(n36532) );
  AND2X1 U37399 ( .A(n61296), .B(n61295), .Y(n36533) );
  AND2X1 U37400 ( .A(n38782), .B(n36534), .Y(n65873) );
  NOR2X1 U37401 ( .A(n65978), .B(n65977), .Y(n36534) );
  AND2X1 U37402 ( .A(n36536), .B(n36535), .Y(n69913) );
  INVX1 U37403 ( .A(n40456), .Y(n36535) );
  OR2X1 U37404 ( .A(n41197), .B(n69911), .Y(n36536) );
  OR2X1 U37405 ( .A(n69912), .B(n69913), .Y(n36537) );
  AND2X1 U37406 ( .A(n36538), .B(n36539), .Y(n70201) );
  NAND2X1 U37407 ( .A(n38007), .B(n38074), .Y(n36538) );
  OR2X1 U37408 ( .A(n38053), .B(n69915), .Y(n36539) );
  XOR2X1 U37409 ( .A(n64510), .B(n64245), .Y(n36540) );
  NOR2X1 U37410 ( .A(n39418), .B(n39419), .Y(n36541) );
  XNOR2X1 U37411 ( .A(n69885), .B(n36542), .Y(n69574) );
  XOR2X1 U37412 ( .A(n69540), .B(n43523), .Y(n36542) );
  XOR2X1 U37413 ( .A(n69559), .B(n69558), .Y(n36543) );
  XOR2X1 U37414 ( .A(n41033), .B(n69574), .Y(n36544) );
  AND2X1 U37415 ( .A(n70783), .B(n36545), .Y(n70784) );
  INVX1 U37416 ( .A(n43514), .Y(n36545) );
  OR2X1 U37417 ( .A(n36546), .B(n70190), .Y(n71129) );
  INVX1 U37418 ( .A(n43691), .Y(n36546) );
  OR2X1 U37419 ( .A(n36547), .B(n70200), .Y(n70806) );
  INVX1 U37420 ( .A(n36436), .Y(n36547) );
  OR2X1 U37421 ( .A(n70479), .B(n38047), .Y(n36548) );
  INVX1 U37422 ( .A(n36548), .Y(n38046) );
  NAND2X1 U37423 ( .A(n70481), .B(n70480), .Y(n36549) );
  AND2X1 U37424 ( .A(n36549), .B(n36550), .Y(n70483) );
  AND2X1 U37425 ( .A(n38047), .B(n36548), .Y(n36550) );
  NOR2X1 U37426 ( .A(n41029), .B(n40395), .Y(n36551) );
  OR2X1 U37427 ( .A(n36552), .B(n69583), .Y(n69555) );
  INVX1 U37428 ( .A(n43505), .Y(n36552) );
  NOR2X1 U37429 ( .A(n36554), .B(n36555), .Y(n36553) );
  INVX1 U37430 ( .A(n36553), .Y(n61575) );
  AND2X1 U37431 ( .A(n61572), .B(n40156), .Y(n36554) );
  AND2X1 U37432 ( .A(n42024), .B(n61573), .Y(n36555) );
  NOR2X1 U37433 ( .A(n36557), .B(n36558), .Y(n36556) );
  INVX1 U37434 ( .A(n36556), .Y(n61582) );
  AND2X1 U37435 ( .A(n61594), .B(n61579), .Y(n36557) );
  AND2X1 U37436 ( .A(n42051), .B(n61581), .Y(n36558) );
  XNOR2X1 U37437 ( .A(n70171), .B(n38049), .Y(n36559) );
  XNOR2X1 U37438 ( .A(n70171), .B(n38049), .Y(n36560) );
  XOR2X1 U37439 ( .A(n71109), .B(n41281), .Y(n36561) );
  OR2X1 U37440 ( .A(n36563), .B(n36562), .Y(n70791) );
  INVX1 U37441 ( .A(n70790), .Y(n36562) );
  OR2X1 U37442 ( .A(n43508), .B(n36561), .Y(n36563) );
  XOR2X1 U37443 ( .A(n41020), .B(n41028), .Y(n36564) );
  OR2X1 U37444 ( .A(n40395), .B(n41029), .Y(n36565) );
  XOR2X1 U37445 ( .A(n64638), .B(n41292), .Y(n36566) );
  OR2X1 U37446 ( .A(n39314), .B(n39315), .Y(n36567) );
  OR2X1 U37447 ( .A(n39696), .B(n39697), .Y(n36568) );
  AND2X1 U37448 ( .A(n70803), .B(n40456), .Y(n36569) );
  INVX1 U37449 ( .A(n36569), .Y(n71125) );
  NAND2X1 U37450 ( .A(n71704), .B(n71703), .Y(n36570) );
  NAND2X1 U37451 ( .A(n40457), .B(n36571), .Y(n38969) );
  NOR2X1 U37452 ( .A(n36572), .B(n72657), .Y(n36571) );
  INVX1 U37453 ( .A(n72732), .Y(n36572) );
  AND2X1 U37454 ( .A(n70821), .B(n70820), .Y(n36573) );
  AND2X1 U37455 ( .A(n38818), .B(n36574), .Y(n72111) );
  INVX1 U37456 ( .A(n37357), .Y(n36574) );
  NAND2X1 U37457 ( .A(n72126), .B(n36575), .Y(u_muldiv_result_r[30]) );
  NOR2X1 U37458 ( .A(n72121), .B(n72120), .Y(n36575) );
  NAND2X1 U37459 ( .A(n71704), .B(n71703), .Y(n36576) );
  OR2X1 U37460 ( .A(n36577), .B(n36578), .Y(n69171) );
  OR2X1 U37461 ( .A(n69166), .B(n38144), .Y(n36577) );
  OR2X1 U37462 ( .A(n69297), .B(n43588), .Y(n36578) );
  NOR2X1 U37463 ( .A(n36580), .B(n36581), .Y(n36579) );
  INVX1 U37464 ( .A(n36579), .Y(n61429) );
  AND2X1 U37465 ( .A(n61445), .B(n61426), .Y(n36580) );
  NOR2X1 U37466 ( .A(n39322), .B(n39323), .Y(n36581) );
  OR2X1 U37467 ( .A(n39088), .B(n39089), .Y(n36582) );
  INVX1 U37468 ( .A(n36582), .Y(n38925) );
  OR2X1 U37469 ( .A(n39112), .B(n62377), .Y(n36583) );
  NOR2X1 U37470 ( .A(n36583), .B(n36584), .Y(n38721) );
  OR2X1 U37471 ( .A(n36585), .B(n39110), .Y(n36584) );
  INVX1 U37472 ( .A(n63140), .Y(n36585) );
  OR2X1 U37473 ( .A(n65288), .B(n38457), .Y(n36586) );
  OR2X1 U37474 ( .A(n65288), .B(n38457), .Y(n36587) );
  NAND2X1 U37475 ( .A(n69197), .B(n36591), .Y(n36588) );
  NAND2X1 U37476 ( .A(n36588), .B(n36589), .Y(n38826) );
  OR2X1 U37477 ( .A(n36590), .B(n69283), .Y(n36589) );
  INVX1 U37478 ( .A(n69284), .Y(n36590) );
  AND2X1 U37479 ( .A(n69196), .B(n69284), .Y(n36591) );
  OR2X1 U37480 ( .A(n36593), .B(n36592), .Y(n65667) );
  INVX1 U37481 ( .A(n65293), .Y(n36592) );
  OR2X1 U37482 ( .A(n41557), .B(n41608), .Y(n36593) );
  OR2X1 U37483 ( .A(n65918), .B(n36594), .Y(n65919) );
  INVX1 U37484 ( .A(n43672), .Y(n36594) );
  OR2X1 U37485 ( .A(n36595), .B(n36596), .Y(n66931) );
  AND2X1 U37486 ( .A(n66588), .B(n43649), .Y(n36595) );
  AND2X1 U37487 ( .A(n66593), .B(n66592), .Y(n36596) );
  OR2X1 U37488 ( .A(n36597), .B(n39769), .Y(n63142) );
  NOR2X1 U37489 ( .A(n38720), .B(n38721), .Y(n36597) );
  INVX1 U37490 ( .A(opcode_opcode_w[22]), .Y(n36598) );
  INVX1 U37491 ( .A(n36598), .Y(n36599) );
  OR2X1 U37492 ( .A(n42469), .B(n42763), .Y(n36600) );
  OR2X1 U37493 ( .A(n40604), .B(n42740), .Y(n36601) );
  OR2X1 U37494 ( .A(n40623), .B(n40624), .Y(n36602) );
  AND2X1 U37495 ( .A(n40753), .B(n40754), .Y(n36603) );
  AND2X1 U37496 ( .A(n70239), .B(n70238), .Y(n36604) );
  OR2X1 U37497 ( .A(n36605), .B(n36606), .Y(n70900) );
  AND2X1 U37498 ( .A(n70565), .B(n43573), .Y(n36605) );
  AND2X1 U37499 ( .A(n70566), .B(n38889), .Y(n36606) );
  OR2X1 U37500 ( .A(n38646), .B(n38647), .Y(n36607) );
  OR2X1 U37501 ( .A(n42469), .B(n42763), .Y(n36608) );
  OR2X1 U37502 ( .A(n42702), .B(n46326), .Y(n36609) );
  INVX1 U37503 ( .A(n42892), .Y(n36610) );
  OR2X1 U37504 ( .A(n36611), .B(n66926), .Y(n67261) );
  INVX1 U37505 ( .A(n43522), .Y(n36611) );
  OR2X1 U37506 ( .A(n36612), .B(n36613), .Y(n64949) );
  OR2X1 U37507 ( .A(n41562), .B(n42005), .Y(n36612) );
  OR2X1 U37508 ( .A(n41535), .B(n40052), .Y(n36613) );
  OR2X1 U37509 ( .A(n36614), .B(n36615), .Y(n66494) );
  OR2X1 U37510 ( .A(n41302), .B(n40225), .Y(n36614) );
  AND2X1 U37511 ( .A(n66008), .B(n66007), .Y(n36615) );
  OR2X1 U37512 ( .A(n36616), .B(n65478), .Y(n65658) );
  INVX1 U37513 ( .A(n65656), .Y(n36616) );
  AND2X1 U37514 ( .A(n59231), .B(n59123), .Y(n36617) );
  AND2X1 U37515 ( .A(n59715), .B(n59718), .Y(n36618) );
  OR2X1 U37516 ( .A(n39471), .B(n36785), .Y(n36619) );
  AND2X1 U37517 ( .A(n45265), .B(n45266), .Y(n36620) );
  NOR2X1 U37518 ( .A(n42351), .B(n42352), .Y(n36621) );
  OR2X1 U37519 ( .A(n36622), .B(n36623), .Y(n69291) );
  INVX1 U37520 ( .A(n41426), .Y(n36622) );
  OR2X1 U37521 ( .A(n39958), .B(n69849), .Y(n36623) );
  OR2X1 U37522 ( .A(n38283), .B(n36624), .Y(n68908) );
  INVX1 U37523 ( .A(n43670), .Y(n36624) );
  OR2X1 U37524 ( .A(n40539), .B(n40540), .Y(n36625) );
  AND2X1 U37525 ( .A(n66032), .B(n36626), .Y(n66030) );
  INVX1 U37526 ( .A(n66028), .Y(n36626) );
  NAND2X1 U37527 ( .A(n66034), .B(n66033), .Y(n36627) );
  AND2X1 U37528 ( .A(n60563), .B(n60562), .Y(n36628) );
  OR2X1 U37529 ( .A(n36629), .B(n36630), .Y(n63150) );
  INVX1 U37530 ( .A(n63627), .Y(n36629) );
  AND2X1 U37531 ( .A(n41922), .B(n63629), .Y(n36630) );
  XOR2X1 U37532 ( .A(n72686), .B(n39430), .Y(n36631) );
  OR2X1 U37533 ( .A(n36633), .B(n36632), .Y(n64370) );
  INVX1 U37534 ( .A(n64366), .Y(n36632) );
  OR2X1 U37535 ( .A(n41111), .B(n41372), .Y(n36633) );
  OR2X1 U37536 ( .A(n36634), .B(n36635), .Y(n71690) );
  INVX1 U37537 ( .A(n71184), .Y(n36634) );
  AND2X1 U37538 ( .A(n71183), .B(n71182), .Y(n36635) );
  AND2X1 U37539 ( .A(n59130), .B(n59175), .Y(n36636) );
  OR2X1 U37540 ( .A(n36637), .B(n36636), .Y(n59161) );
  INVX1 U37541 ( .A(n41751), .Y(n36637) );
  AND2X1 U37542 ( .A(n66015), .B(n36586), .Y(n36638) );
  INVX1 U37543 ( .A(n36638), .Y(n66475) );
  OR2X1 U37544 ( .A(n71776), .B(n36639), .Y(n72093) );
  NAND2X1 U37545 ( .A(n36640), .B(n71781), .Y(n36639) );
  OR2X1 U37546 ( .A(n71775), .B(n72137), .Y(n36640) );
  AND2X1 U37547 ( .A(n36641), .B(n38623), .Y(n64952) );
  INVX1 U37548 ( .A(n43977), .Y(n36641) );
  XOR2X1 U37549 ( .A(n70163), .B(n70162), .Y(n36642) );
  OR2X1 U37550 ( .A(n36643), .B(n36644), .Y(n62955) );
  AND2X1 U37551 ( .A(n40237), .B(n63250), .Y(n36643) );
  AND2X1 U37552 ( .A(n62954), .B(n63245), .Y(n36644) );
  AND2X1 U37553 ( .A(n63178), .B(n36645), .Y(n63177) );
  INVX1 U37554 ( .A(n63175), .Y(n36645) );
  OR2X1 U37555 ( .A(n36638), .B(n36646), .Y(n66476) );
  OR2X1 U37556 ( .A(n39029), .B(n41257), .Y(n36646) );
  NOR2X1 U37557 ( .A(n66938), .B(n36648), .Y(n36647) );
  INVX1 U37558 ( .A(n36647), .Y(n67282) );
  INVX1 U37559 ( .A(n43625), .Y(n36648) );
  AND2X1 U37560 ( .A(n36649), .B(n36650), .Y(n62437) );
  OR2X1 U37561 ( .A(n62432), .B(n40553), .Y(n36649) );
  OR2X1 U37562 ( .A(n62433), .B(n62432), .Y(n36650) );
  AND2X1 U37563 ( .A(n36652), .B(n36651), .Y(n63176) );
  INVX1 U37564 ( .A(n63175), .Y(n36651) );
  OR2X1 U37565 ( .A(n40419), .B(n40420), .Y(n36652) );
  NAND2X1 U37566 ( .A(n39386), .B(n60941), .Y(n36653) );
  OR2X1 U37567 ( .A(n36655), .B(n36654), .Y(n71711) );
  INVX1 U37568 ( .A(n43692), .Y(n36654) );
  XOR2X1 U37569 ( .A(n71143), .B(n71148), .Y(n36655) );
  AND2X1 U37570 ( .A(n64136), .B(n64137), .Y(n36656) );
  AND2X1 U37571 ( .A(n65715), .B(n40987), .Y(n36657) );
  AND2X1 U37572 ( .A(n64179), .B(n64180), .Y(n36658) );
  NAND2X1 U37573 ( .A(n64379), .B(n64707), .Y(n36659) );
  OR2X1 U37574 ( .A(n36660), .B(n36661), .Y(n65966) );
  AND2X1 U37575 ( .A(n43653), .B(n65932), .Y(n36660) );
  NOR2X1 U37576 ( .A(n38489), .B(n38490), .Y(n36661) );
  OR2X1 U37577 ( .A(n36662), .B(n61151), .Y(n36664) );
  INVX1 U37578 ( .A(n61150), .Y(n36662) );
  INVX1 U37579 ( .A(n61149), .Y(n36663) );
  INVX1 U37580 ( .A(n40534), .Y(n36665) );
  AND2X1 U37581 ( .A(n39798), .B(n36666), .Y(n67194) );
  NOR2X1 U37582 ( .A(n36667), .B(n43573), .Y(n36666) );
  AND2X1 U37583 ( .A(n67556), .B(n67555), .Y(n36667) );
  INVX1 U37584 ( .A(n67646), .Y(n36668) );
  OR2X1 U37585 ( .A(n36669), .B(n66824), .Y(n36671) );
  INVX1 U37586 ( .A(n66823), .Y(n36669) );
  INVX1 U37587 ( .A(n66822), .Y(n36670) );
  AND2X1 U37588 ( .A(n36673), .B(n36672), .Y(n39327) );
  INVX1 U37589 ( .A(n43528), .Y(n36672) );
  NAND2X1 U37590 ( .A(n40123), .B(n70766), .Y(n36673) );
  AND2X1 U37591 ( .A(n67990), .B(n43559), .Y(n36674) );
  INVX1 U37592 ( .A(n36674), .Y(n68583) );
  OR2X1 U37593 ( .A(n36675), .B(n36676), .Y(n68594) );
  AND2X1 U37594 ( .A(n43562), .B(n68582), .Y(n36675) );
  AND2X1 U37595 ( .A(n68589), .B(n68588), .Y(n36676) );
  AND2X1 U37596 ( .A(n65356), .B(n65355), .Y(n36677) );
  INVX1 U37597 ( .A(n68921), .Y(n36678) );
  AND2X1 U37598 ( .A(n36680), .B(n36679), .Y(n68875) );
  INVX1 U37599 ( .A(n43528), .Y(n36679) );
  XOR2X1 U37600 ( .A(n68872), .B(n68871), .Y(n36680) );
  OR2X1 U37601 ( .A(n36681), .B(n66824), .Y(n36683) );
  INVX1 U37602 ( .A(n66320), .Y(n36681) );
  INVX1 U37603 ( .A(n66822), .Y(n36682) );
  NOR2X1 U37604 ( .A(n38393), .B(n39994), .Y(n36684) );
  AND2X1 U37605 ( .A(n59769), .B(n59768), .Y(n36685) );
  NOR2X1 U37606 ( .A(n36687), .B(n36688), .Y(n36686) );
  INVX1 U37607 ( .A(n36686), .Y(n61073) );
  AND2X1 U37608 ( .A(n60719), .B(n39462), .Y(n36687) );
  NOR2X1 U37609 ( .A(n60720), .B(n38724), .Y(n36688) );
  AND2X1 U37610 ( .A(n63885), .B(n63884), .Y(n36689) );
  OR2X1 U37611 ( .A(n36691), .B(n36690), .Y(n65657) );
  INVX1 U37612 ( .A(n65645), .Y(n36690) );
  OR2X1 U37613 ( .A(n41349), .B(n41576), .Y(n36691) );
  AND2X1 U37614 ( .A(n36693), .B(n36692), .Y(n66029) );
  INVX1 U37615 ( .A(n66028), .Y(n36692) );
  OR2X1 U37616 ( .A(n66027), .B(n66026), .Y(n36693) );
  XNOR2X1 U37617 ( .A(n67178), .B(n67177), .Y(n36694) );
  OR2X1 U37618 ( .A(n36696), .B(n36695), .Y(n68582) );
  INVX1 U37619 ( .A(n68584), .Y(n36695) );
  OR2X1 U37620 ( .A(n68497), .B(n68496), .Y(n36696) );
  XNOR2X1 U37621 ( .A(n63629), .B(n63022), .Y(n36697) );
  OR2X1 U37622 ( .A(n36698), .B(n36699), .Y(n64862) );
  INVX1 U37623 ( .A(n42004), .Y(n36698) );
  AND2X1 U37624 ( .A(n64860), .B(n64859), .Y(n36699) );
  OR2X1 U37625 ( .A(n36700), .B(n36701), .Y(n64021) );
  INVX1 U37626 ( .A(n37318), .Y(n36700) );
  NOR2X1 U37627 ( .A(n39467), .B(n39468), .Y(n36701) );
  NOR2X1 U37628 ( .A(n41132), .B(n39101), .Y(n36702) );
  XOR2X1 U37629 ( .A(n41130), .B(n65168), .Y(n36703) );
  XOR2X1 U37630 ( .A(n67663), .B(n36704), .Y(n68264) );
  OR2X1 U37631 ( .A(n67562), .B(n67561), .Y(n36704) );
  XOR2X1 U37632 ( .A(n67571), .B(n67570), .Y(n36705) );
  AND2X1 U37633 ( .A(n39650), .B(n39604), .Y(n36706) );
  AND2X1 U37634 ( .A(opcode_opcode_w[24]), .B(n42761), .Y(n36707) );
  AND2X1 U37635 ( .A(opcode_opcode_w[24]), .B(n42761), .Y(n36708) );
  AND2X1 U37636 ( .A(n36702), .B(n65130), .Y(n36709) );
  OR2X1 U37637 ( .A(n40450), .B(n36713), .Y(n36710) );
  AND2X1 U37638 ( .A(n36710), .B(n36711), .Y(n59727) );
  OR2X1 U37639 ( .A(n36712), .B(n59725), .Y(n36711) );
  INVX1 U37640 ( .A(n59924), .Y(n36712) );
  OR2X1 U37641 ( .A(n40451), .B(n36712), .Y(n36713) );
  OR2X1 U37642 ( .A(n40824), .B(n42798), .Y(n36714) );
  NOR2X1 U37643 ( .A(n46215), .B(n46214), .Y(n36715) );
  AND2X1 U37644 ( .A(n64345), .B(n64346), .Y(n36716) );
  INVX1 U37645 ( .A(n36716), .Y(n64690) );
  OR2X1 U37646 ( .A(n36717), .B(n36718), .Y(n60978) );
  OR2X1 U37647 ( .A(n61203), .B(n62423), .Y(n36717) );
  AND2X1 U37648 ( .A(n39193), .B(n39238), .Y(n36718) );
  AND2X1 U37649 ( .A(n42376), .B(n36714), .Y(n36719) );
  OR2X1 U37650 ( .A(n60938), .B(n36653), .Y(n36720) );
  OR2X1 U37651 ( .A(n38685), .B(n38686), .Y(n36721) );
  AND2X1 U37652 ( .A(n59128), .B(n59134), .Y(n36722) );
  AND2X1 U37653 ( .A(n59672), .B(n59673), .Y(n36723) );
  AND2X1 U37654 ( .A(n68561), .B(n68560), .Y(n36724) );
  OR2X1 U37655 ( .A(n40254), .B(n40255), .Y(n36725) );
  AND2X1 U37656 ( .A(n63767), .B(n63768), .Y(n36726) );
  AND2X1 U37657 ( .A(n65522), .B(n65523), .Y(n36727) );
  OR2X1 U37658 ( .A(n40237), .B(n36728), .Y(n62952) );
  INVX1 U37659 ( .A(n63244), .Y(n36728) );
  OR2X1 U37660 ( .A(n36730), .B(n36729), .Y(n68460) );
  INVX1 U37661 ( .A(n43616), .Y(n36729) );
  OR2X1 U37662 ( .A(n68768), .B(n68189), .Y(n36730) );
  OR2X1 U37663 ( .A(n39544), .B(n39545), .Y(n36731) );
  OR2X1 U37664 ( .A(n67669), .B(n36732), .Y(n68011) );
  INVX1 U37665 ( .A(n42992), .Y(n36732) );
  AND2X1 U37666 ( .A(n42671), .B(n46014), .Y(n36733) );
  XOR2X1 U37667 ( .A(n59710), .B(n59902), .Y(n36734) );
  XOR2X1 U37668 ( .A(n41025), .B(n36678), .Y(n36735) );
  NOR2X1 U37669 ( .A(n46016), .B(n46015), .Y(n36736) );
  OR2X1 U37670 ( .A(n36737), .B(n36738), .Y(n59918) );
  AND2X1 U37671 ( .A(n59917), .B(n59916), .Y(n36737) );
  AND2X1 U37672 ( .A(n59912), .B(n59911), .Y(n36738) );
  AND2X1 U37673 ( .A(n63604), .B(n63605), .Y(n36739) );
  NOR2X1 U37674 ( .A(n64850), .B(n64849), .Y(n36740) );
  OR2X1 U37675 ( .A(n36741), .B(n36742), .Y(n60203) );
  INVX1 U37676 ( .A(n60202), .Y(n36741) );
  NOR2X1 U37677 ( .A(n60200), .B(n41739), .Y(n36742) );
  NOR2X1 U37678 ( .A(n36744), .B(n36745), .Y(n36743) );
  INVX1 U37679 ( .A(n36743), .Y(n61266) );
  AND2X1 U37680 ( .A(n60913), .B(n60912), .Y(n36744) );
  AND2X1 U37681 ( .A(n60924), .B(n60923), .Y(n36745) );
  NOR2X1 U37682 ( .A(n42488), .B(n46382), .Y(n36746) );
  NOR2X1 U37683 ( .A(n45681), .B(n46013), .Y(n36747) );
  NOR2X1 U37684 ( .A(n38798), .B(n37144), .Y(n36748) );
  XOR2X1 U37685 ( .A(n60101), .B(n39458), .Y(n36749) );
  NOR2X1 U37686 ( .A(n67875), .B(n67280), .Y(n36750) );
  NOR2X1 U37687 ( .A(n67647), .B(n67568), .Y(n36751) );
  OR2X1 U37688 ( .A(n61219), .B(n61220), .Y(n61223) );
  XNOR2X1 U37689 ( .A(n69536), .B(n69214), .Y(n36752) );
  XNOR2X1 U37690 ( .A(n36754), .B(n60694), .Y(n36753) );
  INVX1 U37691 ( .A(n36753), .Y(n60576) );
  XOR2X1 U37692 ( .A(n60699), .B(n39205), .Y(n36754) );
  XOR2X1 U37693 ( .A(n71386), .B(n71094), .Y(n71226) );
  OR2X1 U37694 ( .A(n65714), .B(n65719), .Y(n66057) );
  XOR2X1 U37695 ( .A(n68037), .B(n68031), .Y(n68465) );
  XOR2X1 U37696 ( .A(n68560), .B(n68554), .Y(n68557) );
  XNOR2X1 U37697 ( .A(n36756), .B(n39859), .Y(n36755) );
  INVX1 U37698 ( .A(n36755), .Y(n61127) );
  XOR2X1 U37699 ( .A(n61226), .B(n38309), .Y(n36756) );
  OR2X1 U37700 ( .A(n38432), .B(n40014), .Y(n62431) );
  OR2X1 U37701 ( .A(n42335), .B(n42336), .Y(n36757) );
  AND2X1 U37702 ( .A(n35938), .B(n45157), .Y(n36758) );
  AND2X1 U37703 ( .A(opcode_opcode_w[23]), .B(opcode_opcode_w[24]), .Y(n36759)
         );
  AND2X1 U37704 ( .A(n43612), .B(n43810), .Y(n36760) );
  NOR2X1 U37705 ( .A(n71433), .B(n38047), .Y(n36762) );
  AND2X1 U37706 ( .A(n66507), .B(n43625), .Y(n36763) );
  XOR2X1 U37707 ( .A(n59466), .B(n59465), .Y(n36764) );
  AND2X1 U37708 ( .A(n72834), .B(n73503), .Y(n36765) );
  AND2X1 U37709 ( .A(n42308), .B(n73520), .Y(n36766) );
  AND2X1 U37710 ( .A(n37537), .B(n37336), .Y(n36767) );
  AND2X1 U37711 ( .A(n64185), .B(n64372), .Y(n36768) );
  AND2X1 U37712 ( .A(n66317), .B(n66316), .Y(n36769) );
  XOR2X1 U37713 ( .A(n59385), .B(n36437), .Y(n36770) );
  XNOR2X1 U37714 ( .A(n59307), .B(n59306), .Y(n36771) );
  OR2X1 U37715 ( .A(n38642), .B(n38643), .Y(n36772) );
  XOR2X1 U37716 ( .A(n65721), .B(n65722), .Y(n36773) );
  XOR2X1 U37717 ( .A(n65298), .B(n65297), .Y(n36774) );
  AND2X1 U37718 ( .A(n69278), .B(n69277), .Y(n36775) );
  NAND2X1 U37719 ( .A(n40528), .B(n42761), .Y(n36776) );
  XOR2X1 U37720 ( .A(n63577), .B(n63844), .Y(n36777) );
  XOR2X1 U37721 ( .A(n71415), .B(n39866), .Y(n36778) );
  AND2X1 U37722 ( .A(n64076), .B(n64075), .Y(n36779) );
  AND2X1 U37723 ( .A(n70034), .B(n70032), .Y(n36780) );
  AND2X1 U37724 ( .A(n42383), .B(n42227), .Y(n36781) );
  XOR2X1 U37725 ( .A(n62827), .B(n62557), .Y(n36782) );
  AND2X1 U37726 ( .A(n47620), .B(n47619), .Y(n36783) );
  XNOR2X1 U37727 ( .A(n60531), .B(n60533), .Y(n36784) );
  AND2X1 U37728 ( .A(n66207), .B(n66206), .Y(n36785) );
  XOR2X1 U37729 ( .A(n59787), .B(n59786), .Y(n36786) );
  XOR2X1 U37730 ( .A(n60266), .B(n60265), .Y(n36787) );
  AND2X1 U37731 ( .A(n43464), .B(n70371), .Y(n36788) );
  OR2X1 U37732 ( .A(n39706), .B(n39707), .Y(n36789) );
  NOR2X1 U37733 ( .A(n40456), .B(n70500), .Y(n36790) );
  AND2X1 U37734 ( .A(n67606), .B(n43698), .Y(n36791) );
  AND2X1 U37735 ( .A(n64880), .B(n43661), .Y(n36828) );
  AND2X1 U37736 ( .A(n40485), .B(n43943), .Y(n37318) );
  AND2X1 U37737 ( .A(n43724), .B(n43992), .Y(n37319) );
  AND2X1 U37738 ( .A(n42632), .B(n43992), .Y(n37320) );
  AND2X1 U37739 ( .A(n29534), .B(n29535), .Y(n37333) );
  AND2X1 U37740 ( .A(u_csr_writeback_idx_q[1]), .B(n37537), .Y(n37337) );
  AND2X1 U37741 ( .A(n15971), .B(n15972), .Y(n37340) );
  AND2X1 U37742 ( .A(n73524), .B(n73571), .Y(n37341) );
  AND2X1 U37743 ( .A(n37567), .B(n73522), .Y(n37344) );
  AND2X1 U37744 ( .A(n49716), .B(n42876), .Y(n37354) );
  AND2X1 U37745 ( .A(n45544), .B(n42878), .Y(n37355) );
  XNOR2X1 U37746 ( .A(n67826), .B(n67825), .Y(n37356) );
  NOR2X1 U37747 ( .A(n40456), .B(n72646), .Y(n37357) );
  AND2X1 U37748 ( .A(n64028), .B(n64029), .Y(n37358) );
  AND2X1 U37749 ( .A(n64525), .B(n64524), .Y(n37359) );
  AND2X1 U37750 ( .A(n63723), .B(n63985), .Y(n37360) );
  AND2X1 U37751 ( .A(n61193), .B(n63194), .Y(n37361) );
  AND2X1 U37752 ( .A(n43545), .B(n66526), .Y(n37362) );
  NOR2X1 U37753 ( .A(n36694), .B(n67553), .Y(n37363) );
  NOR2X1 U37754 ( .A(n70208), .B(n41417), .Y(n37364) );
  AND2X1 U37755 ( .A(n68160), .B(n68161), .Y(n37365) );
  AND2X1 U37756 ( .A(n64322), .B(n64321), .Y(n37366) );
  AND2X1 U37757 ( .A(n43653), .B(n68821), .Y(n37367) );
  AND2X1 U37758 ( .A(n68162), .B(n68082), .Y(n37368) );
  AND2X1 U37759 ( .A(n66789), .B(n66788), .Y(n37369) );
  AND2X1 U37760 ( .A(n68693), .B(n69024), .Y(n37370) );
  AND2X1 U37761 ( .A(n59939), .B(n59942), .Y(n37371) );
  AND2X1 U37762 ( .A(n69491), .B(n69492), .Y(n37372) );
  XOR2X1 U37763 ( .A(n62938), .B(n42151), .Y(n37373) );
  AND2X1 U37764 ( .A(n43521), .B(n40952), .Y(n37374) );
  AND2X1 U37765 ( .A(n65639), .B(n41313), .Y(n37375) );
  XOR2X1 U37766 ( .A(n68007), .B(n68006), .Y(n37376) );
  XOR2X1 U37767 ( .A(n59897), .B(n38267), .Y(n37377) );
  XNOR2X1 U37768 ( .A(n59363), .B(n59362), .Y(n37378) );
  OR2X1 U37769 ( .A(n39305), .B(n39829), .Y(n37379) );
  AND2X1 U37770 ( .A(n63020), .B(n63019), .Y(n37380) );
  AND2X1 U37771 ( .A(n63716), .B(n63715), .Y(n37381) );
  XOR2X1 U37772 ( .A(n63128), .B(n41616), .Y(n37382) );
  AND2X1 U37773 ( .A(n64938), .B(n41428), .Y(n37383) );
  AND2X1 U37774 ( .A(n68913), .B(n43549), .Y(n37384) );
  AND2X1 U37775 ( .A(n43547), .B(n67208), .Y(n37385) );
  AND2X1 U37776 ( .A(n65112), .B(n65696), .Y(n37386) );
  AND2X1 U37777 ( .A(n68063), .B(n68310), .Y(n37387) );
  AND2X1 U37778 ( .A(n62411), .B(n62412), .Y(n37388) );
  AND2X1 U37779 ( .A(n72200), .B(n41468), .Y(n37389) );
  OR2X1 U37780 ( .A(n39901), .B(n39902), .Y(n37390) );
  AND2X1 U37781 ( .A(n64753), .B(n64752), .Y(n37391) );
  OR2X1 U37782 ( .A(n42833), .B(n42834), .Y(n37392) );
  XOR2X1 U37783 ( .A(n36570), .B(n71118), .Y(n37393) );
  XOR2X1 U37784 ( .A(n39873), .B(n61092), .Y(n37394) );
  OR2X1 U37785 ( .A(n39648), .B(n39649), .Y(n37395) );
  NAND2X1 U37786 ( .A(n40448), .B(n43018), .Y(n37396) );
  AND2X1 U37787 ( .A(n64805), .B(n65053), .Y(n37397) );
  NAND2X1 U37788 ( .A(n38364), .B(n58130), .Y(n37398) );
  NAND2X1 U37789 ( .A(n38364), .B(n39669), .Y(n37399) );
  XNOR2X1 U37790 ( .A(n60436), .B(n41436), .Y(n37400) );
  AND2X1 U37791 ( .A(n65358), .B(n66044), .Y(n37401) );
  AND2X1 U37792 ( .A(n43631), .B(n70532), .Y(n37402) );
  XOR2X1 U37793 ( .A(n60522), .B(n41635), .Y(n37403) );
  AND2X1 U37794 ( .A(n65204), .B(n43512), .Y(n37404) );
  AND2X1 U37795 ( .A(n61651), .B(n61652), .Y(n37405) );
  AND2X1 U37796 ( .A(n43963), .B(n43775), .Y(n37407) );
  AND2X1 U37797 ( .A(n43870), .B(n43487), .Y(n37408) );
  NAND2X1 U37798 ( .A(n8696), .B(n54382), .Y(n37409) );
  NAND2X1 U37799 ( .A(n8696), .B(n51998), .Y(n37410) );
  NAND2X1 U37800 ( .A(n51998), .B(n43309), .Y(n37411) );
  AND2X1 U37801 ( .A(n43909), .B(n42640), .Y(n37412) );
  AND2X1 U37802 ( .A(n38001), .B(n50043), .Y(n37413) );
  AND2X1 U37803 ( .A(n69409), .B(n69408), .Y(n37414) );
  NAND2X1 U37804 ( .A(n59119), .B(n44057), .Y(n37415) );
  AND2X1 U37805 ( .A(n43772), .B(n44048), .Y(n37416) );
  AND2X1 U37806 ( .A(n66974), .B(n44048), .Y(n37417) );
  OR2X1 U37807 ( .A(n42302), .B(n25786), .Y(n37444) );
  NAND2X1 U37808 ( .A(n25631), .B(n25632), .Y(n37449) );
  AND2X1 U37809 ( .A(n25637), .B(n25638), .Y(n37450) );
  AND2X1 U37810 ( .A(n29060), .B(n1062), .Y(n37454) );
  AND2X1 U37811 ( .A(n42582), .B(n42602), .Y(n37455) );
  AND2X1 U37812 ( .A(n29303), .B(n519), .Y(n37456) );
  AND2X1 U37813 ( .A(n42582), .B(n50831), .Y(n37457) );
  AND2X1 U37814 ( .A(n29222), .B(n73406), .Y(n37458) );
  NAND2X1 U37815 ( .A(n28521), .B(n28522), .Y(n37459) );
  NOR2X1 U37816 ( .A(n29062), .B(n24243), .Y(n37460) );
  AND2X1 U37817 ( .A(n29230), .B(n491), .Y(n37462) );
  AND2X1 U37818 ( .A(n50825), .B(n42588), .Y(n37463) );
  NOR2X1 U37819 ( .A(n29305), .B(n24294), .Y(n37464) );
  NOR2X1 U37820 ( .A(n29224), .B(n24122), .Y(n37465) );
  NOR2X1 U37821 ( .A(n29232), .B(n24115), .Y(n37466) );
  NOR2X1 U37822 ( .A(n29140), .B(n24175), .Y(n37467) );
  AND2X1 U37823 ( .A(n29255), .B(n73407), .Y(n37468) );
  AND2X1 U37824 ( .A(n42585), .B(n42600), .Y(n37469) );
  NOR2X1 U37825 ( .A(n29215), .B(n24129), .Y(n37470) );
  NOR2X1 U37826 ( .A(n29284), .B(n24312), .Y(n37471) );
  AND2X1 U37827 ( .A(n43389), .B(n24109), .Y(n37472) );
  AND2X1 U37828 ( .A(n42446), .B(n50831), .Y(n37473) );
  AND2X1 U37829 ( .A(n29151), .B(n37472), .Y(n37474) );
  NOR2X1 U37830 ( .A(n29074), .B(n24200), .Y(n37475) );
  NOR2X1 U37831 ( .A(n29048), .B(n24184), .Y(n37476) );
  NOR2X1 U37832 ( .A(n29100), .B(n24207), .Y(n37477) );
  NOR2X1 U37833 ( .A(n29119), .B(n24214), .Y(n37478) );
  NOR2X1 U37834 ( .A(n29130), .B(n24221), .Y(n37479) );
  AND2X1 U37835 ( .A(n29152), .B(n37472), .Y(n37480) );
  NOR2X1 U37836 ( .A(n29257), .B(n24341), .Y(n37481) );
  AND2X1 U37837 ( .A(u_csr_writeback_idx_q[4]), .B(n58155), .Y(n37482) );
  NOR2X1 U37838 ( .A(n29295), .B(n24302), .Y(n37484) );
  NOR2X1 U37839 ( .A(n29241), .B(n24357), .Y(n37486) );
  NOR2X1 U37840 ( .A(n29249), .B(n24349), .Y(n37487) );
  NOR2X1 U37841 ( .A(n29265), .B(n24333), .Y(n37488) );
  NOR2X1 U37842 ( .A(n29274), .B(n24323), .Y(n37489) );
  NOR2X1 U37843 ( .A(n29194), .B(n24149), .Y(n37490) );
  NOR2X1 U37844 ( .A(n29204), .B(n24140), .Y(n37491) );
  NOR2X1 U37845 ( .A(n29163), .B(n24192), .Y(n37492) );
  NOR2X1 U37846 ( .A(n29174), .B(n24166), .Y(n37493) );
  NOR2X1 U37847 ( .A(n29183), .B(n24158), .Y(n37494) );
  AND2X1 U37848 ( .A(n42582), .B(n42584), .Y(n37495) );
  AND2X1 U37849 ( .A(n42603), .B(n42582), .Y(n37496) );
  AND2X1 U37850 ( .A(n42590), .B(n42584), .Y(n37497) );
  AND2X1 U37851 ( .A(n29072), .B(n550), .Y(n37498) );
  AND2X1 U37852 ( .A(n29117), .B(n551), .Y(n37499) );
  AND2X1 U37853 ( .A(n42603), .B(n42590), .Y(n37500) );
  AND2X1 U37854 ( .A(n29138), .B(n554), .Y(n37501) );
  AND2X1 U37855 ( .A(n42602), .B(n42590), .Y(n37502) );
  AND2X1 U37856 ( .A(n42589), .B(n42585), .Y(n37503) );
  AND2X1 U37857 ( .A(n29098), .B(n548), .Y(n37504) );
  AND2X1 U37858 ( .A(n42601), .B(n42585), .Y(n37505) );
  AND2X1 U37859 ( .A(n29181), .B(n528), .Y(n37506) );
  AND2X1 U37860 ( .A(n29213), .B(n29214), .Y(n37507) );
  AND2X1 U37861 ( .A(n42602), .B(n42446), .Y(n37508) );
  AND2X1 U37862 ( .A(n29282), .B(n29283), .Y(n37509) );
  AND2X1 U37863 ( .A(n42591), .B(n42602), .Y(n37510) );
  AND2X1 U37864 ( .A(n42584), .B(n42446), .Y(n37511) );
  AND2X1 U37865 ( .A(n29192), .B(n572), .Y(n37512) );
  AND2X1 U37866 ( .A(n42603), .B(n42446), .Y(n37513) );
  AND2X1 U37867 ( .A(n29172), .B(n566), .Y(n37514) );
  AND2X1 U37868 ( .A(n42591), .B(n42584), .Y(n37515) );
  AND2X1 U37869 ( .A(n29263), .B(n498), .Y(n37516) );
  AND2X1 U37870 ( .A(n29247), .B(n494), .Y(n37517) );
  AND2X1 U37871 ( .A(n42603), .B(n42591), .Y(n37518) );
  AND2X1 U37872 ( .A(n29046), .B(n546), .Y(n37519) );
  AND2X1 U37873 ( .A(n42592), .B(n42589), .Y(n37520) );
  AND2X1 U37874 ( .A(n29272), .B(n504), .Y(n37521) );
  AND2X1 U37875 ( .A(n42592), .B(n42600), .Y(n37522) );
  AND2X1 U37876 ( .A(n29128), .B(n544), .Y(n37523) );
  AND2X1 U37877 ( .A(n42594), .B(n42589), .Y(n37524) );
  AND2X1 U37878 ( .A(n29239), .B(n502), .Y(n37525) );
  AND2X1 U37879 ( .A(n42594), .B(n42600), .Y(n37526) );
  AND2X1 U37880 ( .A(n42601), .B(n42592), .Y(n37527) );
  AND2X1 U37881 ( .A(n29202), .B(n530), .Y(n37528) );
  AND2X1 U37882 ( .A(n42601), .B(n42594), .Y(n37529) );
  AND2X1 U37883 ( .A(n29161), .B(n526), .Y(n37530) );
  AND2X1 U37884 ( .A(n29293), .B(n512), .Y(n37532) );
  AND2X1 U37885 ( .A(n50753), .B(n42585), .Y(n37534) );
  AND2X1 U37886 ( .A(n50753), .B(n42594), .Y(n37535) );
  AND2X1 U37887 ( .A(n42592), .B(n50753), .Y(n37536) );
  AND2X1 U37888 ( .A(n43415), .B(n58542), .Y(n37539) );
  AND2X1 U37889 ( .A(u_mmu_state_q[1]), .B(u_mmu_state_q[0]), .Y(n37547) );
  AND2X1 U37890 ( .A(n37547), .B(n55819), .Y(n37548) );
  AND2X1 U37891 ( .A(n42947), .B(n15802), .Y(n37552) );
  AND2X1 U37892 ( .A(n57326), .B(n58543), .Y(n37554) );
  AND2X1 U37893 ( .A(n43374), .B(n44844), .Y(n37555) );
  AND2X1 U37894 ( .A(n43415), .B(n15802), .Y(n37556) );
  AND2X1 U37895 ( .A(n51121), .B(n50636), .Y(n37558) );
  AND2X1 U37896 ( .A(n43441), .B(n73513), .Y(n37560) );
  AND2X1 U37897 ( .A(n50498), .B(n50497), .Y(n37561) );
  AND2X1 U37898 ( .A(n8801), .B(n58506), .Y(n37562) );
  OR2X1 U37899 ( .A(n24533), .B(n24473), .Y(n37565) );
  AND2X1 U37900 ( .A(n58266), .B(n27964), .Y(n37567) );
  AND2X1 U37901 ( .A(n57401), .B(n51408), .Y(n37568) );
  AND2X1 U37902 ( .A(n57411), .B(n50633), .Y(n37570) );
  AND2X1 U37903 ( .A(n50633), .B(n50634), .Y(n37572) );
  AND2X1 U37904 ( .A(u_muldiv_invert_res_q), .B(n37333), .Y(n37575) );
  AND2X1 U37905 ( .A(n524), .B(n44600), .Y(n37577) );
  AND2X1 U37906 ( .A(n539), .B(n44558), .Y(n37579) );
  AND2X1 U37907 ( .A(n531), .B(n44570), .Y(n37580) );
  AND2X1 U37908 ( .A(n535), .B(n44582), .Y(n37581) );
  AND2X1 U37909 ( .A(n501), .B(n44471), .Y(n37584) );
  AND2X1 U37910 ( .A(n57921), .B(n57922), .Y(n37587) );
  AND2X1 U37911 ( .A(u_csr_writeback_idx_q[1]), .B(u_csr_writeback_idx_q[0]), 
        .Y(n37597) );
  OR2X1 U37912 ( .A(n47180), .B(n47179), .Y(n37782) );
  OR2X1 U37913 ( .A(n48969), .B(n31922), .Y(n37783) );
  OR2X1 U37914 ( .A(n49103), .B(n32610), .Y(n37784) );
  OR2X1 U37915 ( .A(n49241), .B(n32743), .Y(n37785) );
  OR2X1 U37916 ( .A(n48834), .B(n34625), .Y(n37786) );
  OR2X1 U37917 ( .A(n47475), .B(n32333), .Y(n37787) );
  OR2X1 U37918 ( .A(n49415), .B(n34221), .Y(n37788) );
  OR2X1 U37919 ( .A(n47348), .B(n34356), .Y(n37789) );
  OR2X1 U37920 ( .A(n48697), .B(n48696), .Y(n37790) );
  OR2X1 U37921 ( .A(n47705), .B(n47704), .Y(n37791) );
  AND2X1 U37922 ( .A(n46974), .B(n42876), .Y(n37792) );
  AND2X1 U37923 ( .A(n49507), .B(n42878), .Y(n37793) );
  AND2X1 U37924 ( .A(n45940), .B(n42878), .Y(n37794) );
  AND2X1 U37925 ( .A(n47051), .B(n42877), .Y(n37795) );
  NOR2X1 U37926 ( .A(\clk_gate_u_fetch_skid_buffer_q_reg_1/n2 ), .B(n73546), 
        .Y(n37796) );
  NOR2X1 U37927 ( .A(\clk_gate_u_fetch_skid_buffer_q_reg_2/n2 ), .B(n73546), 
        .Y(n37797) );
  NOR2X1 U37928 ( .A(\clk_gate_u_fetch_skid_buffer_q_reg_0/n2 ), .B(n73546), 
        .Y(n37798) );
  NOR2X1 U37929 ( .A(\clk_gate_u_decode_pc_q_reg/n2 ), .B(n73546), .Y(n37799)
         );
  NOR2X1 U37930 ( .A(\clk_gate_u_decode_pc_q_reg_0/n2 ), .B(n73546), .Y(n37800) );
  NOR2X1 U37931 ( .A(\clk_gate_u_fetch_skid_buffer_q_reg/n2 ), .B(n73546), .Y(
        n37801) );
  NOR2X1 U37932 ( .A(\clk_gate_u_decode_opcode_instr_q_reg_0/n2 ), .B(n73546), 
        .Y(n37802) );
  NOR2X1 U37933 ( .A(\clk_gate_u_mmu_virt_addr_q_reg/n2 ), .B(n73546), .Y(
        n37803) );
  NOR2X1 U37934 ( .A(\clk_gate_u_fetch_pc_d_q_reg/n2 ), .B(n73546), .Y(n37804)
         );
  NOR2X1 U37935 ( .A(\clk_gate_u_fetch_pc_d_q_reg_0/n2 ), .B(n73546), .Y(
        n37805) );
  NOR2X1 U37936 ( .A(\clk_gate_u_decode_opcode_instr_q_reg/n2 ), .B(n73546), 
        .Y(n37806) );
  NOR2X1 U37937 ( .A(\clk_gate_u_decode_opcode_instr_q_reg_1/n2 ), .B(n73546), 
        .Y(n37807) );
  NOR2X1 U37938 ( .A(\clk_gate_u_mmu_pte_addr_q_reg_0/n2 ), .B(n73546), .Y(
        n37808) );
  NOR2X1 U37939 ( .A(\clk_gate_u_decode_u_regfile_reg_r22_q_reg_0/n2 ), .B(
        n73546), .Y(n37809) );
  NOR2X1 U37940 ( .A(\clk_gate_u_decode_u_regfile_reg_r21_q_reg_0/n2 ), .B(
        n73546), .Y(n37810) );
  NOR2X1 U37941 ( .A(\clk_gate_u_decode_u_regfile_reg_r20_q_reg_0/n2 ), .B(
        n73546), .Y(n37811) );
  NOR2X1 U37942 ( .A(\clk_gate_u_decode_u_regfile_reg_r19_q_reg_0/n2 ), .B(
        n73546), .Y(n37812) );
  NOR2X1 U37943 ( .A(\clk_gate_u_decode_u_regfile_reg_r18_q_reg_0/n2 ), .B(
        n73546), .Y(n37813) );
  NOR2X1 U37944 ( .A(\clk_gate_u_decode_u_regfile_reg_r17_q_reg_0/n2 ), .B(
        n73546), .Y(n37814) );
  NOR2X1 U37945 ( .A(\clk_gate_u_decode_u_regfile_reg_r16_q_reg_0/n2 ), .B(
        n73546), .Y(n37815) );
  NOR2X1 U37946 ( .A(\clk_gate_u_decode_u_regfile_reg_r15_q_reg_0/n2 ), .B(
        n73546), .Y(n37816) );
  NOR2X1 U37947 ( .A(\clk_gate_u_decode_u_regfile_reg_r14_q_reg_0/n2 ), .B(
        n73546), .Y(n37817) );
  NOR2X1 U37948 ( .A(\clk_gate_u_decode_u_regfile_reg_r13_q_reg_0/n2 ), .B(
        n73546), .Y(n37818) );
  NOR2X1 U37949 ( .A(\clk_gate_u_decode_u_regfile_reg_r12_q_reg_0/n2 ), .B(
        n73546), .Y(n37819) );
  NOR2X1 U37950 ( .A(\clk_gate_u_decode_u_regfile_reg_r11_q_reg_0/n2 ), .B(
        n73546), .Y(n37820) );
  NOR2X1 U37951 ( .A(\clk_gate_u_decode_u_regfile_reg_r10_q_reg_0/n2 ), .B(
        n73546), .Y(n37821) );
  NOR2X1 U37952 ( .A(\clk_gate_u_decode_u_regfile_reg_r9_q_reg_0/n2 ), .B(
        n73546), .Y(n37822) );
  NOR2X1 U37953 ( .A(\clk_gate_u_decode_u_regfile_reg_r8_q_reg_0/n2 ), .B(
        n73546), .Y(n37823) );
  NOR2X1 U37954 ( .A(\clk_gate_u_decode_u_regfile_reg_r7_q_reg_0/n2 ), .B(
        n73546), .Y(n37824) );
  NOR2X1 U37955 ( .A(\clk_gate_u_decode_u_regfile_reg_r6_q_reg_0/n2 ), .B(
        n73546), .Y(n37825) );
  NOR2X1 U37956 ( .A(\clk_gate_u_decode_u_regfile_reg_r5_q_reg_0/n2 ), .B(
        n73546), .Y(n37826) );
  NOR2X1 U37957 ( .A(\clk_gate_u_decode_u_regfile_reg_r4_q_reg_0/n2 ), .B(
        n73546), .Y(n37827) );
  NOR2X1 U37958 ( .A(\clk_gate_u_decode_u_regfile_reg_r3_q_reg_0/n2 ), .B(
        n73546), .Y(n37828) );
  NOR2X1 U37959 ( .A(\clk_gate_u_decode_u_regfile_reg_r2_q_reg_0/n2 ), .B(
        n73546), .Y(n37829) );
  NOR2X1 U37960 ( .A(\clk_gate_u_decode_u_regfile_reg_r1_q_reg_0/n2 ), .B(
        n73546), .Y(n37830) );
  NOR2X1 U37961 ( .A(\clk_gate_u_decode_u_regfile_reg_r31_q_reg_0/n2 ), .B(
        n73546), .Y(n37831) );
  NOR2X1 U37962 ( .A(\clk_gate_u_decode_u_regfile_reg_r30_q_reg_0/n2 ), .B(
        n73546), .Y(n37832) );
  NOR2X1 U37963 ( .A(\clk_gate_u_decode_u_regfile_reg_r29_q_reg_0/n2 ), .B(
        n73546), .Y(n37833) );
  NOR2X1 U37964 ( .A(\clk_gate_u_decode_u_regfile_reg_r28_q_reg_0/n2 ), .B(
        n73546), .Y(n37834) );
  NOR2X1 U37965 ( .A(\clk_gate_u_decode_u_regfile_reg_r27_q_reg_0/n2 ), .B(
        n73546), .Y(n37835) );
  NOR2X1 U37966 ( .A(\clk_gate_u_decode_u_regfile_reg_r26_q_reg_0/n2 ), .B(
        n73546), .Y(n37836) );
  NOR2X1 U37967 ( .A(\clk_gate_u_decode_u_regfile_reg_r25_q_reg_0/n2 ), .B(
        n73546), .Y(n37837) );
  NOR2X1 U37968 ( .A(\clk_gate_u_decode_u_regfile_reg_r21_q_reg/n2 ), .B(
        n73546), .Y(n37838) );
  NOR2X1 U37969 ( .A(\clk_gate_u_decode_u_regfile_reg_r8_q_reg/n2 ), .B(n73546), .Y(n37839) );
  NOR2X1 U37970 ( .A(\clk_gate_u_decode_u_regfile_reg_r5_q_reg/n2 ), .B(n73546), .Y(n37840) );
  NOR2X1 U37971 ( .A(\clk_gate_u_decode_u_regfile_reg_r22_q_reg/n2 ), .B(
        n73546), .Y(n37841) );
  NOR2X1 U37972 ( .A(\clk_gate_u_decode_u_regfile_reg_r20_q_reg/n2 ), .B(
        n73546), .Y(n37842) );
  NOR2X1 U37973 ( .A(\clk_gate_u_decode_u_regfile_reg_r19_q_reg/n2 ), .B(
        n73546), .Y(n37843) );
  NOR2X1 U37974 ( .A(\clk_gate_u_decode_u_regfile_reg_r18_q_reg/n2 ), .B(
        n73546), .Y(n37844) );
  NOR2X1 U37975 ( .A(\clk_gate_u_decode_u_regfile_reg_r17_q_reg/n2 ), .B(
        n73546), .Y(n37845) );
  NOR2X1 U37976 ( .A(\clk_gate_u_decode_u_regfile_reg_r16_q_reg/n2 ), .B(
        n73546), .Y(n37846) );
  NOR2X1 U37977 ( .A(\clk_gate_u_decode_u_regfile_reg_r15_q_reg/n2 ), .B(
        n73546), .Y(n37847) );
  NOR2X1 U37978 ( .A(\clk_gate_u_decode_u_regfile_reg_r14_q_reg/n2 ), .B(
        n73546), .Y(n37848) );
  NOR2X1 U37979 ( .A(\clk_gate_u_decode_u_regfile_reg_r13_q_reg/n2 ), .B(
        n73546), .Y(n37849) );
  NOR2X1 U37980 ( .A(\clk_gate_u_decode_u_regfile_reg_r12_q_reg/n2 ), .B(
        n73546), .Y(n37850) );
  NOR2X1 U37981 ( .A(\clk_gate_u_decode_u_regfile_reg_r11_q_reg/n2 ), .B(
        n73546), .Y(n37851) );
  NOR2X1 U37982 ( .A(\clk_gate_u_decode_u_regfile_reg_r10_q_reg/n2 ), .B(
        n73546), .Y(n37852) );
  NOR2X1 U37983 ( .A(\clk_gate_u_decode_u_regfile_reg_r9_q_reg/n2 ), .B(n73546), .Y(n37853) );
  NOR2X1 U37984 ( .A(\clk_gate_u_decode_u_regfile_reg_r7_q_reg/n2 ), .B(n73546), .Y(n37854) );
  NOR2X1 U37985 ( .A(\clk_gate_u_decode_u_regfile_reg_r6_q_reg/n2 ), .B(n73546), .Y(n37855) );
  NOR2X1 U37986 ( .A(\clk_gate_u_decode_u_regfile_reg_r4_q_reg/n2 ), .B(n73546), .Y(n37856) );
  NOR2X1 U37987 ( .A(\clk_gate_u_decode_u_regfile_reg_r3_q_reg/n2 ), .B(n73546), .Y(n37857) );
  NOR2X1 U37988 ( .A(\clk_gate_u_decode_u_regfile_reg_r2_q_reg/n2 ), .B(n73546), .Y(n37858) );
  NOR2X1 U37989 ( .A(\clk_gate_u_decode_u_regfile_reg_r31_q_reg/n2 ), .B(
        n73546), .Y(n37859) );
  NOR2X1 U37990 ( .A(\clk_gate_u_decode_u_regfile_reg_r30_q_reg/n2 ), .B(
        n73546), .Y(n37860) );
  NOR2X1 U37991 ( .A(\clk_gate_u_decode_u_regfile_reg_r29_q_reg/n2 ), .B(
        n73546), .Y(n37861) );
  NOR2X1 U37992 ( .A(\clk_gate_u_decode_u_regfile_reg_r28_q_reg/n2 ), .B(
        n73546), .Y(n37862) );
  NOR2X1 U37993 ( .A(\clk_gate_u_decode_u_regfile_reg_r27_q_reg/n2 ), .B(
        n73546), .Y(n37863) );
  NOR2X1 U37994 ( .A(\clk_gate_u_decode_u_regfile_reg_r26_q_reg/n2 ), .B(
        n73546), .Y(n37864) );
  NOR2X1 U37995 ( .A(\clk_gate_u_decode_u_regfile_reg_r1_q_reg/n2 ), .B(n73546), .Y(n37865) );
  NOR2X1 U37996 ( .A(\clk_gate_u_fetch_branch_pc_q_reg_0/n2 ), .B(n73546), .Y(
        n37866) );
  NOR2X1 U37997 ( .A(\clk_gate_u_fetch_branch_pc_q_reg/n2 ), .B(n73546), .Y(
        n37867) );
  NOR2X1 U37998 ( .A(\clk_gate_u_lsu_mem_data_wr_q_reg_0/n2 ), .B(n73546), .Y(
        n37868) );
  NOR2X1 U37999 ( .A(\clk_gate_u_lsu_mem_cacheable_q_reg/n2 ), .B(n73546), .Y(
        n37869) );
  NOR2X1 U38000 ( .A(\clk_gate_u_decode_inst_q_reg/n2 ), .B(n73546), .Y(n37870) );
  NOR2X1 U38001 ( .A(\clk_gate_u_mmu_itlb_entry_q_reg_0/n2 ), .B(n73546), .Y(
        n37871) );
  NOR2X1 U38002 ( .A(\clk_gate_u_mmu_dtlb_entry_q_reg_0/n2 ), .B(n73546), .Y(
        n37872) );
  NOR2X1 U38003 ( .A(\clk_gate_u_mmu_lsu_in_addr_q_reg_0/n2 ), .B(n73546), .Y(
        n37873) );
  NOR2X1 U38004 ( .A(\clk_gate_u_lsu_mem_addr_q_reg_0/n2 ), .B(n73546), .Y(
        n37874) );
  NOR2X1 U38005 ( .A(\clk_gate_u_mmu_lsu_in_addr_q_reg/n2 ), .B(n73546), .Y(
        n37875) );
  NOR2X1 U38006 ( .A(\clk_gate_u_lsu_mem_addr_q_reg/n2 ), .B(n73546), .Y(
        n37876) );
  NOR2X1 U38007 ( .A(\clk_gate_u_decode_u_regfile_reg_r23_q_reg/n2 ), .B(
        n73546), .Y(n37877) );
  NOR2X1 U38008 ( .A(\clk_gate_u_decode_u_regfile_reg_r24_q_reg/n2 ), .B(
        n73546), .Y(n37878) );
  NOR2X1 U38009 ( .A(\clk_gate_u_decode_u_regfile_reg_r25_q_reg/n2 ), .B(
        n73546), .Y(n37879) );
  NOR2X1 U38010 ( .A(\clk_gate_u_decode_u_regfile_reg_r23_q_reg_0/n2 ), .B(
        n73546), .Y(n37880) );
  NOR2X1 U38011 ( .A(\clk_gate_u_decode_u_regfile_reg_r24_q_reg_0/n2 ), .B(
        n73546), .Y(n37881) );
  NOR2X1 U38012 ( .A(\clk_gate_u_fetch_fetch_pc_q_reg/n2 ), .B(n73546), .Y(
        n37882) );
  NOR2X1 U38013 ( .A(\clk_gate_u_fetch_fetch_pc_q_reg_0/n2 ), .B(n73546), .Y(
        n37883) );
  NOR2X1 U38014 ( .A(\clk_gate_u_mmu_pte_addr_q_reg/n2 ), .B(n73546), .Y(
        n37884) );
  NOR2X1 U38015 ( .A(\clk_gate_u_decode_opcode_instr_q_reg_2/n2 ), .B(n73546), 
        .Y(n37885) );
  OR2X1 U38016 ( .A(n40044), .B(n40043), .Y(n37886) );
  OR2X1 U38017 ( .A(n36828), .B(n37887), .Y(n65197) );
  AND2X1 U38018 ( .A(n41154), .B(n64882), .Y(n37887) );
  NOR2X1 U38019 ( .A(n37889), .B(n37890), .Y(n37888) );
  INVX1 U38020 ( .A(n37888), .Y(n60873) );
  AND2X1 U38021 ( .A(n61308), .B(n38456), .Y(n37889) );
  AND2X1 U38022 ( .A(n41982), .B(n60871), .Y(n37890) );
  NOR2X1 U38023 ( .A(n38874), .B(n38875), .Y(n37891) );
  XOR2X1 U38024 ( .A(n37892), .B(n67599), .Y(n67604) );
  OR2X1 U38025 ( .A(n40124), .B(n37921), .Y(n37892) );
  NOR2X1 U38026 ( .A(n37894), .B(n37895), .Y(n37893) );
  INVX1 U38027 ( .A(n37893), .Y(n49925) );
  AND2X1 U38028 ( .A(n54658), .B(n49922), .Y(n37894) );
  AND2X1 U38029 ( .A(n49924), .B(n54657), .Y(n37895) );
  INVX1 U38030 ( .A(n37999), .Y(n37896) );
  OR2X1 U38031 ( .A(n37897), .B(n38000), .Y(n49988) );
  NAND2X1 U38032 ( .A(n37896), .B(n49986), .Y(n37897) );
  NOR2X1 U38033 ( .A(n37899), .B(n37900), .Y(n37898) );
  INVX1 U38034 ( .A(n37898), .Y(n49933) );
  AND2X1 U38035 ( .A(n54823), .B(n49930), .Y(n37899) );
  AND2X1 U38036 ( .A(n49932), .B(n54822), .Y(n37900) );
  INVX1 U38037 ( .A(n54706), .Y(n37901) );
  AND2X1 U38038 ( .A(n54705), .B(n37902), .Y(n54709) );
  NOR2X1 U38039 ( .A(n37901), .B(n54707), .Y(n37902) );
  AND2X1 U38040 ( .A(n62731), .B(n62730), .Y(n37903) );
  AND2X1 U38041 ( .A(n63406), .B(n63405), .Y(n37904) );
  NOR2X1 U38042 ( .A(n40332), .B(n40333), .Y(n37905) );
  XOR2X1 U38043 ( .A(n37905), .B(n64270), .Y(n37906) );
  OR2X1 U38044 ( .A(n66564), .B(n43717), .Y(n66913) );
  AND2X1 U38045 ( .A(n37933), .B(n37934), .Y(n37907) );
  NAND2X1 U38046 ( .A(n66553), .B(n66552), .Y(n37908) );
  XNOR2X1 U38047 ( .A(n67595), .B(n40731), .Y(n37909) );
  XNOR2X1 U38048 ( .A(n37910), .B(n65227), .Y(n65223) );
  XOR2X1 U38049 ( .A(n65226), .B(n43509), .Y(n37910) );
  XNOR2X1 U38050 ( .A(n65937), .B(n65936), .Y(n37911) );
  OR2X1 U38051 ( .A(n37912), .B(n37913), .Y(n65225) );
  OR2X1 U38052 ( .A(n41226), .B(n65218), .Y(n37912) );
  AND2X1 U38053 ( .A(n65222), .B(n65221), .Y(n37913) );
  AND2X1 U38054 ( .A(n65225), .B(n65224), .Y(n37914) );
  NAND2X1 U38055 ( .A(n43706), .B(n66564), .Y(n37915) );
  NOR2X1 U38056 ( .A(n37918), .B(n37917), .Y(n37916) );
  INVX1 U38057 ( .A(n66916), .Y(n37917) );
  AND2X1 U38058 ( .A(n43706), .B(n66564), .Y(n37918) );
  OR2X1 U38059 ( .A(n40263), .B(n37919), .Y(n65937) );
  AND2X1 U38060 ( .A(n41470), .B(n65584), .Y(n37919) );
  OR2X1 U38061 ( .A(n64573), .B(n43717), .Y(n64576) );
  OR2X1 U38062 ( .A(n39143), .B(n39144), .Y(n37920) );
  AND2X1 U38063 ( .A(n37907), .B(n67245), .Y(n37921) );
  XNOR2X1 U38064 ( .A(n66919), .B(n66905), .Y(n37922) );
  OR2X1 U38065 ( .A(n38038), .B(n38039), .Y(n37923) );
  AND2X1 U38066 ( .A(n62325), .B(n62324), .Y(n37924) );
  AND2X1 U38067 ( .A(n61425), .B(n61424), .Y(n37925) );
  OR2X1 U38068 ( .A(n38853), .B(n38854), .Y(n37926) );
  NOR2X1 U38069 ( .A(n65196), .B(n37928), .Y(n37927) );
  INVX1 U38070 ( .A(n43661), .Y(n37928) );
  OR2X1 U38071 ( .A(n40325), .B(n40326), .Y(n37929) );
  XNOR2X1 U38072 ( .A(n37930), .B(n37931), .Y(n65947) );
  AND2X1 U38073 ( .A(n65956), .B(n65953), .Y(n37930) );
  XOR2X1 U38074 ( .A(n37929), .B(n65935), .Y(n37931) );
  NOR2X1 U38075 ( .A(n40263), .B(n65945), .Y(n37932) );
  NAND2X1 U38076 ( .A(n38023), .B(n66915), .Y(n37933) );
  OR2X1 U38077 ( .A(n43707), .B(n66917), .Y(n37934) );
  AND2X1 U38078 ( .A(n67917), .B(n67914), .Y(n37935) );
  OR2X1 U38079 ( .A(n37936), .B(n37935), .Y(n67905) );
  INVX1 U38080 ( .A(n67912), .Y(n37936) );
  AND2X1 U38081 ( .A(n64253), .B(n64252), .Y(n37937) );
  INVX1 U38082 ( .A(n37937), .Y(n64258) );
  XOR2X1 U38083 ( .A(n36393), .B(n37938), .Y(n68228) );
  XOR2X1 U38084 ( .A(n68529), .B(n43708), .Y(n37938) );
  NOR2X1 U38085 ( .A(n37940), .B(n37941), .Y(n37939) );
  INVX1 U38086 ( .A(n37939), .Y(n54395) );
  AND2X1 U38087 ( .A(n51926), .B(n51924), .Y(n37940) );
  AND2X1 U38088 ( .A(n49906), .B(n51923), .Y(n37941) );
  AND2X1 U38089 ( .A(n49910), .B(n49909), .Y(n37942) );
  OR2X1 U38090 ( .A(n37943), .B(n37944), .Y(n54460) );
  AND2X1 U38091 ( .A(n54514), .B(n54516), .Y(n37943) );
  AND2X1 U38092 ( .A(n49912), .B(n54513), .Y(n37944) );
  OR2X1 U38093 ( .A(n37945), .B(n37946), .Y(n54972) );
  AND2X1 U38094 ( .A(n54899), .B(n49938), .Y(n37945) );
  AND2X1 U38095 ( .A(n49940), .B(n54898), .Y(n37946) );
  NOR2X1 U38096 ( .A(n37948), .B(n37949), .Y(n37947) );
  AND2X1 U38097 ( .A(n61422), .B(n40179), .Y(n37948) );
  AND2X1 U38098 ( .A(n41997), .B(n61423), .Y(n37949) );
  AND2X1 U38099 ( .A(n61920), .B(n61919), .Y(n37950) );
  AND2X1 U38100 ( .A(n61940), .B(n61939), .Y(n37951) );
  OR2X1 U38101 ( .A(n68529), .B(n43717), .Y(n68530) );
  AND2X1 U38102 ( .A(n49917), .B(n49916), .Y(n37952) );
  OR2X1 U38103 ( .A(n37953), .B(n37954), .Y(n50293) );
  AND2X1 U38104 ( .A(n50375), .B(n50377), .Y(n37953) );
  AND2X1 U38105 ( .A(n49951), .B(n50374), .Y(n37954) );
  XOR2X1 U38106 ( .A(n68528), .B(n68527), .Y(n37955) );
  OR2X1 U38107 ( .A(n37956), .B(n37957), .Y(n61699) );
  AND2X1 U38108 ( .A(n61792), .B(n61696), .Y(n37956) );
  AND2X1 U38109 ( .A(n41924), .B(n61697), .Y(n37957) );
  OR2X1 U38110 ( .A(n38057), .B(n38058), .Y(n37958) );
  NOR2X1 U38111 ( .A(n37960), .B(n37961), .Y(n37959) );
  INVX1 U38112 ( .A(n37959), .Y(n50357) );
  AND2X1 U38113 ( .A(n49966), .B(n49965), .Y(n37960) );
  AND2X1 U38114 ( .A(n49968), .B(n50078), .Y(n37961) );
  OR2X1 U38115 ( .A(n37962), .B(n37963), .Y(n50451) );
  AND2X1 U38116 ( .A(n50355), .B(n50357), .Y(n37962) );
  AND2X1 U38117 ( .A(n49971), .B(n50354), .Y(n37963) );
  NOR2X1 U38118 ( .A(n37965), .B(n37966), .Y(n37964) );
  INVX1 U38119 ( .A(n37964), .Y(n62107) );
  AND2X1 U38120 ( .A(n62104), .B(n62105), .Y(n37965) );
  AND2X1 U38121 ( .A(n42058), .B(n62106), .Y(n37966) );
  NAND2X1 U38122 ( .A(n40771), .B(n40772), .Y(n37967) );
  AND2X1 U38123 ( .A(n62119), .B(n42098), .Y(n37968) );
  OR2X1 U38124 ( .A(n37968), .B(n37969), .Y(n62121) );
  OR2X1 U38125 ( .A(n37970), .B(n38091), .Y(n37969) );
  INVX1 U38126 ( .A(n62137), .Y(n37970) );
  AND2X1 U38127 ( .A(n62123), .B(n62122), .Y(n37971) );
  AND2X1 U38128 ( .A(n62755), .B(n62754), .Y(n37972) );
  OR2X1 U38129 ( .A(n37973), .B(n37974), .Y(n64562) );
  AND2X1 U38130 ( .A(n43707), .B(n64276), .Y(n37973) );
  AND2X1 U38131 ( .A(n64279), .B(n64278), .Y(n37974) );
  OR2X1 U38132 ( .A(n65557), .B(n37975), .Y(n65595) );
  INVX1 U38133 ( .A(n43683), .Y(n37975) );
  AND2X1 U38134 ( .A(n45535), .B(n42373), .Y(n37976) );
  OR2X1 U38135 ( .A(n61734), .B(n61762), .Y(n61735) );
  OR2X1 U38136 ( .A(n37977), .B(n39091), .Y(n68843) );
  AND2X1 U38137 ( .A(n43505), .B(n68841), .Y(n37977) );
  OR2X1 U38138 ( .A(n37978), .B(n37979), .Y(n49381) );
  AND2X1 U38139 ( .A(n2760), .B(n49674), .Y(n37978) );
  AND2X1 U38140 ( .A(n2774), .B(n42625), .Y(n37979) );
  OR2X1 U38141 ( .A(n61563), .B(n61605), .Y(n61564) );
  OR2X1 U38142 ( .A(n37980), .B(n37981), .Y(n61710) );
  AND2X1 U38143 ( .A(n61706), .B(n61707), .Y(n37980) );
  AND2X1 U38144 ( .A(n41954), .B(n61708), .Y(n37981) );
  OR2X1 U38145 ( .A(n43715), .B(n67605), .Y(n67912) );
  OR2X1 U38146 ( .A(n39459), .B(n39460), .Y(n37982) );
  OR2X1 U38147 ( .A(n38487), .B(n38488), .Y(n37983) );
  NOR2X1 U38148 ( .A(n37985), .B(n37986), .Y(n37984) );
  INVX1 U38149 ( .A(n37984), .Y(n50312) );
  AND2X1 U38150 ( .A(n54971), .B(n54972), .Y(n37985) );
  AND2X1 U38151 ( .A(n49944), .B(n54970), .Y(n37986) );
  OR2X1 U38152 ( .A(n37987), .B(n37988), .Y(n50377) );
  AND2X1 U38153 ( .A(n50311), .B(n50312), .Y(n37987) );
  AND2X1 U38154 ( .A(n49947), .B(n50310), .Y(n37988) );
  NOR2X1 U38155 ( .A(n37990), .B(n37991), .Y(n37989) );
  INVX1 U38156 ( .A(n37989), .Y(n50330) );
  AND2X1 U38157 ( .A(n50291), .B(n50293), .Y(n37990) );
  AND2X1 U38158 ( .A(n49955), .B(n50290), .Y(n37991) );
  OR2X1 U38159 ( .A(n37992), .B(n37993), .Y(n50152) );
  AND2X1 U38160 ( .A(n50328), .B(n50330), .Y(n37992) );
  AND2X1 U38161 ( .A(n49958), .B(n50327), .Y(n37993) );
  NOR2X1 U38162 ( .A(n41161), .B(n41162), .Y(n37994) );
  NOR2X1 U38163 ( .A(n37996), .B(n37997), .Y(n37995) );
  INVX1 U38164 ( .A(n37995), .Y(n50169) );
  AND2X1 U38165 ( .A(n50449), .B(n50451), .Y(n37996) );
  AND2X1 U38166 ( .A(n49975), .B(n50448), .Y(n37997) );
  NOR2X1 U38167 ( .A(n37999), .B(n38000), .Y(n37998) );
  INVX1 U38168 ( .A(n37998), .Y(n49985) );
  AND2X1 U38169 ( .A(n50425), .B(n49981), .Y(n37999) );
  AND2X1 U38170 ( .A(n49984), .B(n50424), .Y(n38000) );
  AND2X1 U38171 ( .A(n8696), .B(n50042), .Y(n38001) );
  AND2X1 U38172 ( .A(n38001), .B(n50043), .Y(n38002) );
  AND2X1 U38173 ( .A(n66926), .B(n43529), .Y(n38003) );
  INVX1 U38174 ( .A(n38003), .Y(n67258) );
  OR2X1 U38175 ( .A(n38004), .B(n38005), .Y(n67617) );
  OR2X1 U38176 ( .A(n67263), .B(n67262), .Y(n38004) );
  AND2X1 U38177 ( .A(n43522), .B(n67264), .Y(n38005) );
  AND2X1 U38178 ( .A(n70186), .B(n69563), .Y(n38006) );
  AND2X1 U38179 ( .A(n66922), .B(n43515), .Y(n66923) );
  OR2X1 U38180 ( .A(n40021), .B(n40022), .Y(n38007) );
  OR2X1 U38181 ( .A(n38008), .B(n38009), .Y(n49404) );
  OR2X1 U38182 ( .A(n49381), .B(n49380), .Y(n38008) );
  OR2X1 U38183 ( .A(n49389), .B(n49388), .Y(n38009) );
  OR2X1 U38184 ( .A(n38010), .B(n38011), .Y(n61741) );
  INVX1 U38185 ( .A(n42065), .Y(n38010) );
  NOR2X1 U38186 ( .A(n61740), .B(n61739), .Y(n38011) );
  OR2X1 U38187 ( .A(n38012), .B(n38013), .Y(n67248) );
  OR2X1 U38188 ( .A(n66575), .B(n66574), .Y(n38012) );
  NOR2X1 U38189 ( .A(n40716), .B(n66579), .Y(n38013) );
  OR2X1 U38190 ( .A(n38014), .B(n36791), .Y(n67611) );
  AND2X1 U38191 ( .A(n67613), .B(n43698), .Y(n38014) );
  OR2X1 U38192 ( .A(n38015), .B(n38016), .Y(n67923) );
  OR2X1 U38193 ( .A(n36507), .B(n67593), .Y(n38015) );
  AND2X1 U38194 ( .A(n66925), .B(n39510), .Y(n38016) );
  NOR2X1 U38195 ( .A(n38018), .B(n38019), .Y(n38017) );
  INVX1 U38196 ( .A(n38017), .Y(n61556) );
  AND2X1 U38197 ( .A(n61554), .B(n39688), .Y(n38018) );
  AND2X1 U38198 ( .A(n41961), .B(n61555), .Y(n38019) );
  NAND2X1 U38199 ( .A(n39258), .B(n65946), .Y(n38020) );
  NAND2X1 U38200 ( .A(n38020), .B(n38021), .Y(n40043) );
  AND2X1 U38201 ( .A(n38022), .B(n39257), .Y(n38021) );
  INVX1 U38202 ( .A(n41465), .Y(n38022) );
  AND2X1 U38203 ( .A(n66914), .B(n37916), .Y(n38023) );
  AND2X1 U38204 ( .A(n38024), .B(n38025), .Y(n68531) );
  OR2X1 U38205 ( .A(n67914), .B(n67913), .Y(n38024) );
  AND2X1 U38206 ( .A(n67917), .B(n67916), .Y(n38025) );
  OR2X1 U38207 ( .A(n38026), .B(n61494), .Y(n61647) );
  AND2X1 U38208 ( .A(n61498), .B(n61497), .Y(n38026) );
  AND2X1 U38209 ( .A(n62311), .B(n62312), .Y(n38027) );
  NAND2X1 U38210 ( .A(n42412), .B(n38084), .Y(n38028) );
  OR2X1 U38211 ( .A(n38028), .B(n38029), .Y(n42410) );
  OR2X1 U38212 ( .A(n38030), .B(n38045), .Y(n38029) );
  INVX1 U38213 ( .A(n38094), .Y(n38030) );
  OR2X1 U38214 ( .A(n68537), .B(n38031), .Y(n38072) );
  NAND2X1 U38215 ( .A(n43710), .B(n40456), .Y(n38031) );
  NOR2X1 U38216 ( .A(n36537), .B(n38033), .Y(n38032) );
  AND2X1 U38217 ( .A(n36436), .B(n38007), .Y(n38033) );
  MX2X1 U38218 ( .A(n70197), .B(n70198), .S0(n43721), .Y(u_muldiv_result_r[24]) );
  NOR2X1 U38219 ( .A(n38035), .B(n38036), .Y(n38034) );
  INVX1 U38220 ( .A(n38034), .Y(n62214) );
  AND2X1 U38221 ( .A(n62651), .B(n62211), .Y(n38035) );
  AND2X1 U38222 ( .A(n41846), .B(n62212), .Y(n38036) );
  NOR2X1 U38223 ( .A(n38038), .B(n38039), .Y(n38037) );
  AND2X1 U38224 ( .A(n62306), .B(n62307), .Y(n38038) );
  AND2X1 U38225 ( .A(n42087), .B(n62308), .Y(n38039) );
  NOR2X1 U38226 ( .A(n38041), .B(n38042), .Y(n38040) );
  INVX1 U38227 ( .A(n38040), .Y(n62017) );
  AND2X1 U38228 ( .A(n62206), .B(n36388), .Y(n38041) );
  AND2X1 U38229 ( .A(n62204), .B(n62015), .Y(n38042) );
  NAND2X1 U38230 ( .A(n42416), .B(n38043), .Y(n42400) );
  AND2X1 U38231 ( .A(mem_i_pc_o[8]), .B(mem_i_pc_o[10]), .Y(n38043) );
  AND2X1 U38232 ( .A(n15), .B(n12), .Y(n38044) );
  NOR2X1 U38233 ( .A(n38045), .B(n42404), .Y(n42413) );
  INVX1 U38234 ( .A(n38044), .Y(n38045) );
  NOR2X1 U38235 ( .A(n38069), .B(n36790), .Y(n38052) );
  INVX1 U38236 ( .A(n43682), .Y(n38047) );
  XNOR2X1 U38237 ( .A(n70171), .B(n38049), .Y(n38048) );
  INVX1 U38238 ( .A(n36559), .Y(n70486) );
  INVX1 U38239 ( .A(n36642), .Y(n38049) );
  NAND2X1 U38240 ( .A(n38052), .B(n70201), .Y(n38050) );
  AND2X1 U38241 ( .A(n38050), .B(n38051), .Y(n70797) );
  OR2X1 U38242 ( .A(n36790), .B(n70812), .Y(n38051) );
  AND2X1 U38243 ( .A(n70200), .B(n43710), .Y(n38053) );
  NAND2X1 U38244 ( .A(n42415), .B(n38054), .Y(n42407) );
  AND2X1 U38245 ( .A(n21), .B(n24), .Y(n38054) );
  NOR2X1 U38246 ( .A(n41159), .B(n41160), .Y(n38055) );
  OR2X1 U38247 ( .A(n69241), .B(n43717), .Y(n69240) );
  NOR2X1 U38248 ( .A(n38057), .B(n38058), .Y(n38056) );
  AND2X1 U38249 ( .A(n61945), .B(n61934), .Y(n38057) );
  AND2X1 U38250 ( .A(n42099), .B(n61936), .Y(n38058) );
  OR2X1 U38251 ( .A(n38059), .B(n38060), .Y(n66552) );
  AND2X1 U38252 ( .A(n66240), .B(n66241), .Y(n38059) );
  AND2X1 U38253 ( .A(n43706), .B(n37911), .Y(n38060) );
  AND2X1 U38254 ( .A(n68837), .B(n69220), .Y(n38061) );
  AND2X1 U38255 ( .A(n43705), .B(n69241), .Y(n38062) );
  AND2X1 U38256 ( .A(n62079), .B(n62078), .Y(n38063) );
  INVX1 U38257 ( .A(n39640), .Y(n38064) );
  OR2X1 U38258 ( .A(n38120), .B(n38121), .Y(n38065) );
  AND2X1 U38259 ( .A(n62774), .B(n62773), .Y(n38066) );
  OR2X1 U38260 ( .A(n38067), .B(n38068), .Y(n72730) );
  AND2X1 U38261 ( .A(n62795), .B(n62794), .Y(n38067) );
  AND2X1 U38262 ( .A(n42130), .B(n62796), .Y(n38068) );
  NOR2X1 U38263 ( .A(n40456), .B(n70200), .Y(n38069) );
  INVX1 U38264 ( .A(n38069), .Y(n70805) );
  NOR2X1 U38265 ( .A(n38238), .B(n38239), .Y(n38070) );
  AND2X1 U38266 ( .A(n62281), .B(n62280), .Y(n38071) );
  NAND2X1 U38267 ( .A(n38072), .B(n38073), .Y(n41410) );
  OR2X1 U38268 ( .A(n43709), .B(n68856), .Y(n38073) );
  OR2X1 U38269 ( .A(n61385), .B(n61476), .Y(n61386) );
  OR2X1 U38270 ( .A(n62817), .B(n62818), .Y(n62820) );
  OR2X1 U38271 ( .A(n69560), .B(n36464), .Y(n69898) );
  AND2X1 U38272 ( .A(n70199), .B(n36436), .Y(n38074) );
  NAND2X1 U38273 ( .A(n42402), .B(n38075), .Y(n42398) );
  AND2X1 U38274 ( .A(n8), .B(n10), .Y(n38075) );
  AND2X1 U38275 ( .A(n42411), .B(n18), .Y(n38076) );
  AND2X1 U38276 ( .A(n38076), .B(n38077), .Y(n56618) );
  AND2X1 U38277 ( .A(n16), .B(n14), .Y(n38077) );
  OR2X1 U38278 ( .A(n38078), .B(n38079), .Y(n72113) );
  AND2X1 U38279 ( .A(n62786), .B(n62787), .Y(n38078) );
  AND2X1 U38280 ( .A(n42125), .B(n62788), .Y(n38079) );
  AND2X1 U38281 ( .A(n70201), .B(n70805), .Y(n38080) );
  OR2X1 U38282 ( .A(n38420), .B(n38421), .Y(n38081) );
  AND2X1 U38283 ( .A(n68263), .B(n68264), .Y(n68260) );
  AND2X1 U38284 ( .A(n65661), .B(n37320), .Y(n65653) );
  XNOR2X1 U38285 ( .A(n67661), .B(n38082), .Y(n67647) );
  NOR2X1 U38286 ( .A(n67195), .B(n67194), .Y(n38082) );
  AND2X1 U38287 ( .A(n54577), .B(n54576), .Y(n38083) );
  NAND2X1 U38288 ( .A(n42412), .B(n38084), .Y(n42404) );
  AND2X1 U38289 ( .A(n7), .B(n17), .Y(n38084) );
  AND2X1 U38290 ( .A(n42882), .B(n40513), .Y(n38085) );
  AND2X1 U38291 ( .A(n62118), .B(n38087), .Y(n38088) );
  INVX1 U38292 ( .A(n38520), .Y(n38086) );
  INVX1 U38293 ( .A(n38521), .Y(n38087) );
  OR2X1 U38294 ( .A(n38520), .B(n38521), .Y(n38089) );
  INVX1 U38295 ( .A(n38089), .Y(n38519) );
  NOR2X1 U38296 ( .A(n38091), .B(n38092), .Y(n38090) );
  INVX1 U38297 ( .A(n38090), .Y(n62120) );
  AND2X1 U38298 ( .A(n62139), .B(n38089), .Y(n38091) );
  AND2X1 U38299 ( .A(n42098), .B(n62119), .Y(n38092) );
  AND2X1 U38300 ( .A(n42401), .B(n38093), .Y(n54771) );
  NOR2X1 U38301 ( .A(n54770), .B(n38083), .Y(n38093) );
  AND2X1 U38302 ( .A(n11), .B(n13), .Y(n38094) );
  OR2X1 U38303 ( .A(n38095), .B(n38096), .Y(n66988) );
  AND2X1 U38304 ( .A(n66991), .B(n66987), .Y(n38095) );
  AND2X1 U38305 ( .A(n66985), .B(n40331), .Y(n38096) );
  AND2X1 U38306 ( .A(n41122), .B(n66078), .Y(n38097) );
  OR2X1 U38307 ( .A(n67290), .B(n39295), .Y(n67288) );
  AND2X1 U38308 ( .A(n61149), .B(n38108), .Y(n38098) );
  OR2X1 U38309 ( .A(n39568), .B(n63462), .Y(n38099) );
  OR2X1 U38310 ( .A(n39033), .B(n37363), .Y(n38100) );
  OR2X1 U38311 ( .A(n38101), .B(n48605), .Y(n47973) );
  OR2X1 U38312 ( .A(n48612), .B(n47972), .Y(n38101) );
  OR2X1 U38313 ( .A(n38454), .B(n38455), .Y(n38102) );
  OR2X1 U38314 ( .A(n38103), .B(n38104), .Y(n61585) );
  AND2X1 U38315 ( .A(n61591), .B(n61582), .Y(n38103) );
  NOR2X1 U38316 ( .A(n39627), .B(n39628), .Y(n38104) );
  NAND2X1 U38317 ( .A(n47860), .B(n47859), .Y(n38105) );
  NAND2X1 U38318 ( .A(n47860), .B(n47859), .Y(n38106) );
  AND2X1 U38319 ( .A(n59687), .B(n59686), .Y(n38107) );
  NAND2X1 U38320 ( .A(n61149), .B(n38108), .Y(n61135) );
  NOR2X1 U38321 ( .A(n38109), .B(n61151), .Y(n38108) );
  INVX1 U38322 ( .A(n61150), .Y(n38109) );
  OR2X1 U38323 ( .A(n42348), .B(n42349), .Y(n38110) );
  OR2X1 U38324 ( .A(n42348), .B(n42349), .Y(n38111) );
  NAND2X1 U38325 ( .A(n62013), .B(n62012), .Y(n38112) );
  OR2X1 U38326 ( .A(n38277), .B(n38278), .Y(n38113) );
  INVX1 U38327 ( .A(opcode_opcode_w[15]), .Y(n38114) );
  INVX1 U38328 ( .A(n38114), .Y(n38115) );
  OR2X1 U38329 ( .A(n38116), .B(n36772), .Y(n59144) );
  OR2X1 U38330 ( .A(n62897), .B(n62896), .Y(n38116) );
  OR2X1 U38331 ( .A(n38117), .B(n38118), .Y(n61740) );
  AND2X1 U38332 ( .A(n61759), .B(n61736), .Y(n38117) );
  AND2X1 U38333 ( .A(n42054), .B(n61738), .Y(n38118) );
  NOR2X1 U38334 ( .A(n38120), .B(n38121), .Y(n38119) );
  AND2X1 U38335 ( .A(n63059), .B(n63060), .Y(n38120) );
  AND2X1 U38336 ( .A(n42117), .B(n63063), .Y(n38121) );
  OR2X1 U38337 ( .A(n38122), .B(n38123), .Y(n69245) );
  OR2X1 U38338 ( .A(n68879), .B(n68878), .Y(n38122) );
  OR2X1 U38339 ( .A(n68875), .B(n68874), .Y(n38123) );
  OR2X1 U38340 ( .A(n38124), .B(n38826), .Y(n70137) );
  AND2X1 U38341 ( .A(n41012), .B(n69616), .Y(n38124) );
  OR2X1 U38342 ( .A(n38125), .B(n38126), .Y(n70447) );
  NAND2X1 U38343 ( .A(n70444), .B(n70445), .Y(n38125) );
  AND2X1 U38344 ( .A(n70446), .B(n43623), .Y(n38126) );
  AND2X1 U38345 ( .A(n39886), .B(n70578), .Y(n38127) );
  INVX1 U38346 ( .A(n38127), .Y(n70572) );
  NAND2X1 U38347 ( .A(n71183), .B(n71182), .Y(n38128) );
  AND2X1 U38348 ( .A(n64635), .B(n64634), .Y(n38129) );
  INVX1 U38349 ( .A(n38129), .Y(n64613) );
  OR2X1 U38350 ( .A(n38130), .B(n38172), .Y(n65244) );
  AND2X1 U38351 ( .A(n65179), .B(n65903), .Y(n38130) );
  AND2X1 U38352 ( .A(n68710), .B(n68429), .Y(n38131) );
  OR2X1 U38353 ( .A(n38307), .B(n38308), .Y(n38132) );
  AND2X1 U38354 ( .A(n38133), .B(n38134), .Y(n70769) );
  OR2X1 U38355 ( .A(n70768), .B(n70767), .Y(n38133) );
  OR2X1 U38356 ( .A(n43523), .B(n36642), .Y(n38134) );
  OR2X1 U38357 ( .A(n38135), .B(n38136), .Y(n69884) );
  OR2X1 U38358 ( .A(n40312), .B(n70158), .Y(n38135) );
  AND2X1 U38359 ( .A(n69883), .B(n69882), .Y(n38136) );
  OR2X1 U38360 ( .A(n38137), .B(n38547), .Y(n64301) );
  AND2X1 U38361 ( .A(n63727), .B(n64247), .Y(n38137) );
  OR2X1 U38362 ( .A(n38138), .B(n59495), .Y(n59569) );
  INVX1 U38363 ( .A(n59535), .Y(n38138) );
  AND2X1 U38364 ( .A(n66832), .B(n66834), .Y(n38139) );
  OR2X1 U38365 ( .A(n38140), .B(n38141), .Y(n68054) );
  AND2X1 U38366 ( .A(n68044), .B(n68043), .Y(n38140) );
  AND2X1 U38367 ( .A(n37416), .B(n68048), .Y(n38141) );
  OR2X1 U38368 ( .A(n38143), .B(n38142), .Y(n70913) );
  INVX1 U38369 ( .A(n70744), .Y(n38142) );
  OR2X1 U38370 ( .A(n70573), .B(n38127), .Y(n38143) );
  AND2X1 U38371 ( .A(n43581), .B(n68602), .Y(n38144) );
  INVX1 U38372 ( .A(n38144), .Y(n69167) );
  OR2X1 U38373 ( .A(n40564), .B(n40565), .Y(n38145) );
  OR2X1 U38374 ( .A(n39376), .B(n39377), .Y(n38146) );
  OR2X1 U38375 ( .A(n38147), .B(n38148), .Y(n63099) );
  AND2X1 U38376 ( .A(n63053), .B(n63054), .Y(n38147) );
  AND2X1 U38377 ( .A(n42093), .B(n63056), .Y(n38148) );
  NOR2X1 U38378 ( .A(n39442), .B(n39443), .Y(n38149) );
  AND2X1 U38379 ( .A(n60854), .B(n60853), .Y(n38150) );
  AND2X1 U38380 ( .A(n68602), .B(n68793), .Y(n38151) );
  OR2X1 U38381 ( .A(n38152), .B(n40052), .Y(n65154) );
  OR2X1 U38382 ( .A(n41562), .B(n41535), .Y(n38152) );
  INVX1 U38383 ( .A(n69916), .Y(n38153) );
  INVX1 U38384 ( .A(n38153), .Y(n38154) );
  AND2X1 U38385 ( .A(n68200), .B(n38155), .Y(n68202) );
  NOR2X1 U38386 ( .A(n39927), .B(n68265), .Y(n38155) );
  AND2X1 U38387 ( .A(n38855), .B(n67056), .Y(n38156) );
  OR2X1 U38388 ( .A(n39280), .B(n38159), .Y(n38157) );
  AND2X1 U38389 ( .A(n38157), .B(n38158), .Y(n69410) );
  OR2X1 U38390 ( .A(n37414), .B(n41239), .Y(n38158) );
  OR2X1 U38391 ( .A(n39500), .B(n37414), .Y(n38159) );
  NOR2X1 U38392 ( .A(n41043), .B(n41044), .Y(n38160) );
  NOR2X1 U38393 ( .A(n38162), .B(n38163), .Y(n38161) );
  INVX1 U38394 ( .A(n38161), .Y(n60408) );
  AND2X1 U38395 ( .A(n60532), .B(n60531), .Y(n38162) );
  AND2X1 U38396 ( .A(n41938), .B(n60406), .Y(n38163) );
  NAND2X1 U38397 ( .A(n62365), .B(n62366), .Y(n38164) );
  AND2X1 U38398 ( .A(n41073), .B(n71441), .Y(n38165) );
  INVX1 U38399 ( .A(n38165), .Y(n71762) );
  OR2X1 U38400 ( .A(n49588), .B(n36873), .Y(n38166) );
  OR2X1 U38401 ( .A(n38823), .B(n42784), .Y(n40851) );
  OR2X1 U38402 ( .A(n39548), .B(n39549), .Y(n38167) );
  OR2X1 U38403 ( .A(n43646), .B(n69916), .Y(n69919) );
  AND2X1 U38404 ( .A(n67128), .B(n67375), .Y(n38168) );
  AND2X1 U38405 ( .A(n71805), .B(n71804), .Y(n38169) );
  OR2X1 U38406 ( .A(n38170), .B(n38171), .Y(n72154) );
  AND2X1 U38407 ( .A(n43544), .B(n71807), .Y(n38170) );
  AND2X1 U38408 ( .A(n71809), .B(n72077), .Y(n38171) );
  NOR2X1 U38409 ( .A(n38173), .B(n65180), .Y(n38172) );
  INVX1 U38410 ( .A(n43631), .Y(n38173) );
  XNOR2X1 U38411 ( .A(n40714), .B(n69540), .Y(n38174) );
  OR2X1 U38412 ( .A(n70453), .B(n39747), .Y(n69926) );
  OR2X1 U38413 ( .A(n38175), .B(n38176), .Y(n71155) );
  INVX1 U38414 ( .A(n71434), .Y(n38175) );
  NOR2X1 U38415 ( .A(n38438), .B(n39011), .Y(n38176) );
  OR2X1 U38416 ( .A(n38177), .B(n38178), .Y(n60368) );
  AND2X1 U38417 ( .A(n60332), .B(n60136), .Y(n38177) );
  AND2X1 U38418 ( .A(n41838), .B(n60137), .Y(n38178) );
  AND2X1 U38419 ( .A(n68788), .B(n68787), .Y(n38179) );
  NOR2X1 U38420 ( .A(n38181), .B(n38182), .Y(n38180) );
  INVX1 U38421 ( .A(n38180), .Y(n60495) );
  AND2X1 U38422 ( .A(n36789), .B(n60364), .Y(n38181) );
  AND2X1 U38423 ( .A(n41840), .B(n60365), .Y(n38182) );
  AND2X1 U38424 ( .A(n60523), .B(n60522), .Y(n38183) );
  INVX1 U38425 ( .A(n38183), .Y(n60400) );
  OR2X1 U38426 ( .A(n38184), .B(n38185), .Y(n68140) );
  OR2X1 U38427 ( .A(n67723), .B(n67722), .Y(n38184) );
  OR2X1 U38428 ( .A(n67728), .B(n67732), .Y(n38185) );
  OR2X1 U38429 ( .A(n38186), .B(n38187), .Y(n67731) );
  INVX1 U38430 ( .A(n67448), .Y(n38186) );
  AND2X1 U38431 ( .A(n41001), .B(n67437), .Y(n38187) );
  OR2X1 U38432 ( .A(n36747), .B(n38188), .Y(n46015) );
  NOR2X1 U38433 ( .A(n38744), .B(n38745), .Y(n38188) );
  OR2X1 U38434 ( .A(n42867), .B(n38768), .Y(n45871) );
  AND2X1 U38435 ( .A(n72106), .B(n40456), .Y(n38189) );
  INVX1 U38436 ( .A(n38189), .Y(n72645) );
  OR2X1 U38437 ( .A(n40187), .B(n40188), .Y(n38190) );
  AND2X1 U38438 ( .A(n69631), .B(n69632), .Y(n38191) );
  NOR2X1 U38439 ( .A(n40746), .B(n40747), .Y(n38192) );
  INVX1 U38440 ( .A(n65998), .Y(n38193) );
  AND2X1 U38441 ( .A(n71762), .B(n40967), .Y(n38194) );
  NAND2X1 U38442 ( .A(n68752), .B(n38195), .Y(n40181) );
  AND2X1 U38443 ( .A(n41729), .B(n68753), .Y(n38195) );
  OR2X1 U38444 ( .A(n70755), .B(n70558), .Y(n70758) );
  NAND2X1 U38445 ( .A(n47701), .B(n38198), .Y(n38196) );
  AND2X1 U38446 ( .A(n38196), .B(n38197), .Y(n63209) );
  OR2X1 U38447 ( .A(n39529), .B(n42804), .Y(n38197) );
  AND2X1 U38448 ( .A(n47702), .B(n36783), .Y(n38198) );
  OR2X1 U38449 ( .A(n38199), .B(n38200), .Y(n66031) );
  OR2X1 U38450 ( .A(n37375), .B(n65643), .Y(n38199) );
  AND2X1 U38451 ( .A(n65644), .B(n41313), .Y(n38200) );
  OR2X1 U38452 ( .A(n70781), .B(n38538), .Y(n38201) );
  NOR2X1 U38453 ( .A(n38201), .B(n38202), .Y(n38595) );
  OR2X1 U38454 ( .A(n41454), .B(n71145), .Y(n38202) );
  NAND2X1 U38455 ( .A(n69606), .B(n69605), .Y(n38203) );
  OR2X1 U38456 ( .A(n38204), .B(n36785), .Y(n66482) );
  OR2X1 U38457 ( .A(n41272), .B(n41276), .Y(n38204) );
  AND2X1 U38458 ( .A(n41770), .B(n62938), .Y(n38205) );
  INVX1 U38459 ( .A(n38205), .Y(n63237) );
  OR2X1 U38460 ( .A(n38206), .B(n38207), .Y(n63541) );
  AND2X1 U38461 ( .A(n63238), .B(n63236), .Y(n38206) );
  AND2X1 U38462 ( .A(n63242), .B(n63241), .Y(n38207) );
  AND2X1 U38463 ( .A(n69928), .B(n69927), .Y(n38208) );
  AND2X1 U38464 ( .A(n38888), .B(n66293), .Y(n38209) );
  INVX1 U38465 ( .A(n42681), .Y(n38210) );
  OR2X1 U38466 ( .A(n38615), .B(n38616), .Y(n38211) );
  NAND2X1 U38467 ( .A(n41319), .B(n43588), .Y(n38212) );
  INVX1 U38468 ( .A(n42224), .Y(n38213) );
  OR2X1 U38469 ( .A(n38214), .B(n38215), .Y(n60994) );
  INVX1 U38470 ( .A(n60992), .Y(n38214) );
  AND2X1 U38471 ( .A(n60991), .B(n61009), .Y(n38215) );
  AND2X1 U38472 ( .A(n39682), .B(n60610), .Y(n60611) );
  XOR2X1 U38473 ( .A(n59485), .B(n59484), .Y(n38216) );
  INVX1 U38474 ( .A(n38216), .Y(n59486) );
  AND2X1 U38475 ( .A(n38217), .B(n38218), .Y(n45187) );
  OR2X1 U38476 ( .A(n36880), .B(n45185), .Y(n38217) );
  OR2X1 U38477 ( .A(n36877), .B(n45186), .Y(n38218) );
  XOR2X1 U38478 ( .A(n65179), .B(n65182), .Y(n65192) );
  XNOR2X1 U38479 ( .A(n38220), .B(n41856), .Y(n38219) );
  INVX1 U38480 ( .A(n38219), .Y(n61333) );
  XOR2X1 U38481 ( .A(n60788), .B(n60787), .Y(n38220) );
  OR2X1 U38482 ( .A(n42799), .B(n38221), .Y(n48399) );
  AND2X1 U38483 ( .A(n63200), .B(n42379), .Y(n38221) );
  XNOR2X1 U38484 ( .A(n69316), .B(n38223), .Y(n38222) );
  INVX1 U38485 ( .A(n38222), .Y(n69639) );
  AND2X1 U38486 ( .A(n68963), .B(n69655), .Y(n38223) );
  XOR2X1 U38487 ( .A(n71098), .B(n71190), .Y(n71099) );
  AND2X1 U38488 ( .A(n65800), .B(n65799), .Y(n38224) );
  AND2X1 U38489 ( .A(n60221), .B(n38225), .Y(n60219) );
  INVX1 U38490 ( .A(n60217), .Y(n38225) );
  OR2X1 U38491 ( .A(n38226), .B(n38227), .Y(n59496) );
  INVX1 U38492 ( .A(n59569), .Y(n38226) );
  AND2X1 U38493 ( .A(n59534), .B(n59572), .Y(n38227) );
  OR2X1 U38494 ( .A(n38228), .B(n38229), .Y(n45248) );
  OR2X1 U38495 ( .A(n45243), .B(n45242), .Y(n38228) );
  OR2X1 U38496 ( .A(n45247), .B(n45246), .Y(n38229) );
  OR2X1 U38497 ( .A(n40606), .B(n38230), .Y(n59397) );
  INVX1 U38498 ( .A(n59394), .Y(n38230) );
  XNOR2X1 U38499 ( .A(n38373), .B(n64852), .Y(n64493) );
  NOR2X1 U38500 ( .A(n42366), .B(n45271), .Y(n38231) );
  INVX1 U38501 ( .A(n38231), .Y(n46367) );
  XOR2X1 U38502 ( .A(n59533), .B(n40580), .Y(n38232) );
  INVX1 U38503 ( .A(n38232), .Y(n59582) );
  NOR2X1 U38504 ( .A(n60938), .B(n39385), .Y(n38233) );
  OR2X1 U38505 ( .A(n38234), .B(n38235), .Y(n61195) );
  AND2X1 U38506 ( .A(n42234), .B(n61186), .Y(n38234) );
  AND2X1 U38507 ( .A(n61191), .B(n42153), .Y(n38235) );
  OR2X1 U38508 ( .A(n38236), .B(n38660), .Y(n63313) );
  OR2X1 U38509 ( .A(n63312), .B(n63773), .Y(n38236) );
  AND2X1 U38510 ( .A(n61135), .B(n61157), .Y(n61154) );
  NOR2X1 U38511 ( .A(n38238), .B(n38239), .Y(n38237) );
  INVX1 U38512 ( .A(n38070), .Y(n62278) );
  AND2X1 U38513 ( .A(n62613), .B(n62274), .Y(n38238) );
  AND2X1 U38514 ( .A(n41996), .B(n62276), .Y(n38239) );
  NOR2X1 U38515 ( .A(n60252), .B(n60643), .Y(n38240) );
  INVX1 U38516 ( .A(n38240), .Y(n61011) );
  XNOR2X1 U38517 ( .A(n64327), .B(n38241), .Y(n64240) );
  XOR2X1 U38518 ( .A(n64008), .B(n64328), .Y(n38241) );
  AND2X1 U38519 ( .A(n60130), .B(n60129), .Y(n38242) );
  INVX1 U38520 ( .A(n38242), .Y(n60362) );
  XOR2X1 U38521 ( .A(n38243), .B(n40765), .Y(n64992) );
  INVX1 U38522 ( .A(n65098), .Y(n38243) );
  XOR2X1 U38523 ( .A(n60445), .B(n41911), .Y(n38244) );
  INVX1 U38524 ( .A(n38244), .Y(n60519) );
  OR2X1 U38525 ( .A(n38245), .B(n38246), .Y(n61169) );
  AND2X1 U38526 ( .A(n60945), .B(n40383), .Y(n38245) );
  AND2X1 U38527 ( .A(n61192), .B(n40391), .Y(n38246) );
  XNOR2X1 U38528 ( .A(n59817), .B(n60018), .Y(n38247) );
  INVX1 U38529 ( .A(n38247), .Y(n60020) );
  OR2X1 U38530 ( .A(n38248), .B(n38249), .Y(n62945) );
  INVX1 U38531 ( .A(n62442), .Y(n38248) );
  AND2X1 U38532 ( .A(n62441), .B(n62440), .Y(n38249) );
  OR2X1 U38533 ( .A(n63250), .B(n63249), .Y(n63533) );
  NOR2X1 U38534 ( .A(n38251), .B(n38252), .Y(n38250) );
  INVX1 U38535 ( .A(n38250), .Y(n62563) );
  AND2X1 U38536 ( .A(n61751), .B(n61748), .Y(n38251) );
  NOR2X1 U38537 ( .A(n39085), .B(n39086), .Y(n38252) );
  OR2X1 U38538 ( .A(n59989), .B(n59805), .Y(n59806) );
  XNOR2X1 U38539 ( .A(n60276), .B(n38254), .Y(n38253) );
  XOR2X1 U38540 ( .A(n60271), .B(n60272), .Y(n38254) );
  OR2X1 U38541 ( .A(n38255), .B(n38256), .Y(n63812) );
  OR2X1 U38542 ( .A(n63228), .B(n63227), .Y(n38255) );
  AND2X1 U38543 ( .A(n63233), .B(n63232), .Y(n38256) );
  XNOR2X1 U38544 ( .A(n38258), .B(n62498), .Y(n38257) );
  INVX1 U38545 ( .A(n38257), .Y(n62875) );
  XOR2X1 U38546 ( .A(n63305), .B(n62881), .Y(n38258) );
  AND2X1 U38547 ( .A(n38793), .B(n38259), .Y(n38271) );
  NAND2X1 U38548 ( .A(n39210), .B(n39612), .Y(n38259) );
  OR2X1 U38549 ( .A(n38260), .B(n38593), .Y(n64151) );
  INVX1 U38550 ( .A(n64149), .Y(n38260) );
  AND2X1 U38551 ( .A(n38261), .B(n38262), .Y(n40191) );
  NOR2X1 U38552 ( .A(n68317), .B(n68316), .Y(n38261) );
  NAND2X1 U38553 ( .A(n68319), .B(n68318), .Y(n38262) );
  XNOR2X1 U38554 ( .A(n66286), .B(n66280), .Y(n38263) );
  INVX1 U38555 ( .A(n38263), .Y(n66282) );
  NOR2X1 U38556 ( .A(n38265), .B(n38266), .Y(n38264) );
  INVX1 U38557 ( .A(n38264), .Y(n70046) );
  AND2X1 U38558 ( .A(n69692), .B(n69691), .Y(n38265) );
  AND2X1 U38559 ( .A(n69696), .B(n69695), .Y(n38266) );
  XOR2X1 U38560 ( .A(n39892), .B(n59896), .Y(n38267) );
  INVX1 U38561 ( .A(n38267), .Y(n60259) );
  NOR2X1 U38562 ( .A(n38269), .B(n38270), .Y(n38268) );
  INVX1 U38563 ( .A(n38268), .Y(n60548) );
  AND2X1 U38564 ( .A(n60541), .B(n60542), .Y(n38269) );
  AND2X1 U38565 ( .A(n60544), .B(n60543), .Y(n38270) );
  OR2X1 U38566 ( .A(n42824), .B(n43461), .Y(n59340) );
  XOR2X1 U38567 ( .A(n67357), .B(n67479), .Y(n66795) );
  XOR2X1 U38568 ( .A(writeback_exec_idx_w[2]), .B(n42814), .Y(n45533) );
  OR2X1 U38569 ( .A(n38397), .B(n62875), .Y(n63169) );
  OR2X1 U38570 ( .A(n38272), .B(n38273), .Y(n63594) );
  AND2X1 U38571 ( .A(n63171), .B(n63170), .Y(n38272) );
  AND2X1 U38572 ( .A(n63174), .B(n63173), .Y(n38273) );
  NOR2X1 U38573 ( .A(n38275), .B(n39571), .Y(n38274) );
  INVX1 U38574 ( .A(n38274), .Y(n60933) );
  INVX1 U38575 ( .A(n60930), .Y(n38275) );
  NOR2X1 U38576 ( .A(n38277), .B(n38278), .Y(n38276) );
  AND2X1 U38577 ( .A(n62073), .B(n62074), .Y(n38277) );
  AND2X1 U38578 ( .A(n41978), .B(n62075), .Y(n38278) );
  XNOR2X1 U38579 ( .A(n60873), .B(n61307), .Y(n38279) );
  INVX1 U38580 ( .A(n38279), .Y(n61447) );
  XNOR2X1 U38581 ( .A(n38281), .B(n40601), .Y(n38280) );
  INVX1 U38582 ( .A(n38280), .Y(n59865) );
  XOR2X1 U38583 ( .A(n59868), .B(n59869), .Y(n38281) );
  OR2X1 U38584 ( .A(n39757), .B(n38282), .Y(n63659) );
  NAND2X1 U38585 ( .A(n63902), .B(n63903), .Y(n38282) );
  XOR2X1 U38586 ( .A(n69209), .B(n68906), .Y(n38283) );
  INVX1 U38587 ( .A(n38283), .Y(n69527) );
  XOR2X1 U38588 ( .A(n38284), .B(n69798), .Y(n69685) );
  XOR2X1 U38589 ( .A(n69796), .B(n69795), .Y(n38284) );
  XNOR2X1 U38590 ( .A(n64627), .B(n40762), .Y(n38285) );
  INVX1 U38591 ( .A(n38285), .Y(n64595) );
  NOR2X1 U38592 ( .A(n38287), .B(n38288), .Y(n38286) );
  INVX1 U38593 ( .A(n38286), .Y(n61841) );
  AND2X1 U38594 ( .A(n62002), .B(n61837), .Y(n38287) );
  AND2X1 U38595 ( .A(n41850), .B(n61839), .Y(n38288) );
  OR2X1 U38596 ( .A(n59561), .B(n59491), .Y(n59492) );
  XNOR2X1 U38597 ( .A(n39552), .B(n38290), .Y(n38289) );
  INVX1 U38598 ( .A(n38289), .Y(n60724) );
  XOR2X1 U38599 ( .A(n69318), .B(n68766), .Y(n69304) );
  XOR2X1 U38600 ( .A(n40553), .B(n61202), .Y(n62481) );
  OR2X1 U38601 ( .A(n38291), .B(n38292), .Y(n48119) );
  AND2X1 U38602 ( .A(n48115), .B(n48370), .Y(n38291) );
  AND2X1 U38603 ( .A(n48118), .B(n48205), .Y(n38292) );
  AND2X1 U38604 ( .A(n64072), .B(n63811), .Y(n38293) );
  INVX1 U38605 ( .A(n38293), .Y(n64113) );
  OR2X1 U38606 ( .A(n61119), .B(n61120), .Y(n61124) );
  XNOR2X1 U38607 ( .A(n59325), .B(n59735), .Y(n38294) );
  INVX1 U38608 ( .A(n38294), .Y(n59668) );
  XNOR2X1 U38609 ( .A(n66519), .B(n65243), .Y(n65245) );
  XNOR2X1 U38610 ( .A(n38851), .B(n38296), .Y(n38295) );
  INVX1 U38611 ( .A(n38295), .Y(n63036) );
  XOR2X1 U38612 ( .A(n63372), .B(n63028), .Y(n38296) );
  XNOR2X1 U38613 ( .A(n36617), .B(n59125), .Y(n59189) );
  AND2X1 U38614 ( .A(n63832), .B(n64090), .Y(n38297) );
  INVX1 U38615 ( .A(n38297), .Y(n64394) );
  OR2X1 U38616 ( .A(n38299), .B(n38298), .Y(n66793) );
  INVX1 U38617 ( .A(n67340), .Y(n38298) );
  OR2X1 U38618 ( .A(n40287), .B(n67344), .Y(n38299) );
  OR2X1 U38619 ( .A(n38300), .B(n38301), .Y(n66108) );
  AND2X1 U38620 ( .A(n65803), .B(n65793), .Y(n38300) );
  AND2X1 U38621 ( .A(n65804), .B(n39102), .Y(n38301) );
  XNOR2X1 U38622 ( .A(n70262), .B(n70095), .Y(n38302) );
  INVX1 U38623 ( .A(n38302), .Y(n70578) );
  OR2X1 U38624 ( .A(n38304), .B(n38303), .Y(n66589) );
  INVX1 U38625 ( .A(n66536), .Y(n38303) );
  OR2X1 U38626 ( .A(n66535), .B(n66534), .Y(n38304) );
  AND2X1 U38627 ( .A(n38592), .B(n43609), .Y(n38305) );
  INVX1 U38628 ( .A(n38305), .Y(n63199) );
  NOR2X1 U38629 ( .A(n38307), .B(n38308), .Y(n38306) );
  AND2X1 U38630 ( .A(n61960), .B(n61906), .Y(n38307) );
  AND2X1 U38631 ( .A(n42023), .B(n61908), .Y(n38308) );
  XNOR2X1 U38632 ( .A(n61025), .B(n61219), .Y(n38309) );
  INVX1 U38633 ( .A(n38309), .Y(n61227) );
  INVX1 U38634 ( .A(n43489), .Y(n38310) );
  INVX1 U38635 ( .A(n43489), .Y(n38311) );
  INVX1 U38636 ( .A(n43485), .Y(n38312) );
  INVX1 U38637 ( .A(n43485), .Y(n38313) );
  INVX1 U38638 ( .A(n44250), .Y(n38314) );
  INVX1 U38639 ( .A(n38314), .Y(n38315) );
  INVX1 U38640 ( .A(n38314), .Y(n38316) );
  INVX1 U38641 ( .A(n38314), .Y(n38317) );
  INVX1 U38642 ( .A(n38314), .Y(n38318) );
  INVX1 U38643 ( .A(n44251), .Y(n38319) );
  INVX1 U38644 ( .A(n38319), .Y(n38320) );
  INVX1 U38645 ( .A(n38319), .Y(n38321) );
  INVX1 U38646 ( .A(n38319), .Y(n38322) );
  INVX1 U38647 ( .A(n38319), .Y(n38323) );
  INVX1 U38648 ( .A(n44250), .Y(n38324) );
  INVX1 U38649 ( .A(n38324), .Y(n38325) );
  INVX1 U38650 ( .A(n38324), .Y(n38326) );
  INVX1 U38651 ( .A(n38324), .Y(n38327) );
  INVX1 U38652 ( .A(n38324), .Y(n38328) );
  INVX1 U38653 ( .A(n44250), .Y(n38329) );
  INVX1 U38654 ( .A(n38329), .Y(n38330) );
  INVX1 U38655 ( .A(n38329), .Y(n38331) );
  INVX1 U38656 ( .A(n38329), .Y(n38332) );
  INVX1 U38657 ( .A(n38329), .Y(n38333) );
  INVX1 U38658 ( .A(n44251), .Y(n38334) );
  INVX1 U38659 ( .A(n38334), .Y(n38335) );
  INVX1 U38660 ( .A(n38334), .Y(n38336) );
  INVX1 U38661 ( .A(n38334), .Y(n38337) );
  INVX1 U38662 ( .A(n38334), .Y(n38338) );
  INVX1 U38663 ( .A(n44251), .Y(n38339) );
  INVX1 U38664 ( .A(n38339), .Y(n38340) );
  INVX1 U38665 ( .A(n38339), .Y(n38341) );
  INVX1 U38666 ( .A(n38339), .Y(n38342) );
  INVX1 U38667 ( .A(n38339), .Y(n38343) );
  INVX1 U38668 ( .A(n44228), .Y(n38344) );
  INVX1 U38669 ( .A(n44226), .Y(n38345) );
  INVX1 U38670 ( .A(n44225), .Y(n38346) );
  INVX1 U38671 ( .A(n44224), .Y(n38347) );
  INVX1 U38672 ( .A(n44201), .Y(n38348) );
  INVX1 U38673 ( .A(n38348), .Y(n38349) );
  INVX1 U38674 ( .A(n38348), .Y(n38350) );
  INVX1 U38675 ( .A(n38348), .Y(n38351) );
  INVX1 U38676 ( .A(n38348), .Y(n38352) );
  INVX1 U38677 ( .A(n44251), .Y(n38353) );
  INVX1 U38678 ( .A(n38353), .Y(n38354) );
  INVX1 U38679 ( .A(n38353), .Y(n38355) );
  INVX1 U38680 ( .A(n38353), .Y(n38356) );
  INVX1 U38681 ( .A(n38353), .Y(n38357) );
  INVX1 U38682 ( .A(n44150), .Y(n38358) );
  INVX1 U38683 ( .A(n38358), .Y(n38359) );
  INVX1 U38684 ( .A(n38358), .Y(n38360) );
  INVX1 U38685 ( .A(n38358), .Y(n38361) );
  INVX1 U38686 ( .A(n38358), .Y(n38362) );
  AND2X1 U38687 ( .A(n38890), .B(n64587), .Y(n38363) );
  INVX1 U38688 ( .A(n36482), .Y(n38364) );
  NAND2X1 U38689 ( .A(n68557), .B(n43670), .Y(n38365) );
  OR2X1 U38690 ( .A(n42364), .B(n42363), .Y(n38366) );
  AND2X1 U38691 ( .A(n65156), .B(n38367), .Y(n65492) );
  AND2X1 U38692 ( .A(n65489), .B(n44000), .Y(n38367) );
  OR2X1 U38693 ( .A(n39927), .B(n70889), .Y(n70559) );
  AND2X1 U38694 ( .A(n66967), .B(n66968), .Y(n38368) );
  OR2X1 U38695 ( .A(n38370), .B(n38369), .Y(n40530) );
  INVX1 U38696 ( .A(n66033), .Y(n38369) );
  OR2X1 U38697 ( .A(n66030), .B(n66029), .Y(n38370) );
  NOR2X1 U38698 ( .A(n64485), .B(n38374), .Y(n38371) );
  OR2X1 U38699 ( .A(n38371), .B(n38372), .Y(n64850) );
  AND2X1 U38700 ( .A(n38373), .B(n64491), .Y(n38372) );
  INVX1 U38701 ( .A(n64851), .Y(n38373) );
  OR2X1 U38702 ( .A(n64486), .B(n64851), .Y(n38374) );
  OR2X1 U38703 ( .A(n61300), .B(n37394), .Y(n61093) );
  OR2X1 U38704 ( .A(n38375), .B(n38376), .Y(n60560) );
  AND2X1 U38705 ( .A(n60752), .B(n60556), .Y(n38375) );
  AND2X1 U38706 ( .A(n41991), .B(n60558), .Y(n38376) );
  XOR2X1 U38707 ( .A(n64500), .B(n64499), .Y(n38377) );
  INVX1 U38708 ( .A(n42235), .Y(n38378) );
  INVX1 U38709 ( .A(n42235), .Y(n38379) );
  INVX1 U38710 ( .A(n42235), .Y(n38380) );
  INVX1 U38711 ( .A(n42235), .Y(n38381) );
  INVX1 U38712 ( .A(n42235), .Y(n38382) );
  INVX1 U38713 ( .A(n42235), .Y(n38383) );
  INVX1 U38714 ( .A(n42235), .Y(n38384) );
  INVX1 U38715 ( .A(n38382), .Y(n38385) );
  INVX1 U38716 ( .A(n38382), .Y(n38386) );
  INVX1 U38717 ( .A(n38383), .Y(n38387) );
  XNOR2X1 U38718 ( .A(n41023), .B(n69531), .Y(n38388) );
  INVX1 U38719 ( .A(n37399), .Y(n38389) );
  INVX1 U38720 ( .A(n37399), .Y(n38390) );
  OR2X1 U38721 ( .A(n38391), .B(n38392), .Y(n63326) );
  OR2X1 U38722 ( .A(n38896), .B(n63321), .Y(n38391) );
  OR2X1 U38723 ( .A(n40480), .B(n63325), .Y(n38392) );
  AND2X1 U38724 ( .A(n66298), .B(n66977), .Y(n38393) );
  INVX1 U38725 ( .A(n38393), .Y(n66950) );
  NAND2X1 U38726 ( .A(n66949), .B(n40331), .Y(n38394) );
  NOR2X1 U38727 ( .A(n42353), .B(n42354), .Y(n38395) );
  OR2X1 U38728 ( .A(n64433), .B(n64755), .Y(n64743) );
  XNOR2X1 U38729 ( .A(n38396), .B(n38472), .Y(n61108) );
  XOR2X1 U38730 ( .A(n60900), .B(n60899), .Y(n38396) );
  AND2X1 U38731 ( .A(n62505), .B(n62504), .Y(n38397) );
  OR2X1 U38732 ( .A(n38398), .B(n37381), .Y(n63978) );
  AND2X1 U38733 ( .A(n63714), .B(n63981), .Y(n38398) );
  XOR2X1 U38734 ( .A(n40143), .B(n71702), .Y(n38399) );
  INVX1 U38735 ( .A(n36424), .Y(n38400) );
  INVX1 U38736 ( .A(n37398), .Y(n38401) );
  INVX1 U38737 ( .A(n37398), .Y(n38402) );
  AND2X1 U38738 ( .A(n67850), .B(n38403), .Y(n67543) );
  AND2X1 U38739 ( .A(n67849), .B(n40670), .Y(n38403) );
  INVX1 U38740 ( .A(n41783), .Y(n38404) );
  INVX1 U38741 ( .A(n41783), .Y(n38405) );
  INVX1 U38742 ( .A(n38404), .Y(n38406) );
  INVX1 U38743 ( .A(n38404), .Y(n38407) );
  INVX1 U38744 ( .A(n38404), .Y(n38408) );
  INVX1 U38745 ( .A(n38404), .Y(n38409) );
  INVX1 U38746 ( .A(n38405), .Y(n38410) );
  INVX1 U38747 ( .A(n38405), .Y(n38411) );
  INVX1 U38748 ( .A(n38405), .Y(n38412) );
  INVX1 U38749 ( .A(n38405), .Y(n38413) );
  NOR2X1 U38750 ( .A(n38415), .B(n38416), .Y(n38414) );
  OR2X1 U38751 ( .A(n46235), .B(n45922), .Y(n38415) );
  OR2X1 U38752 ( .A(n46575), .B(n37038), .Y(n38416) );
  OR2X1 U38753 ( .A(n38417), .B(n38418), .Y(n61707) );
  AND2X1 U38754 ( .A(n61786), .B(n61703), .Y(n38417) );
  AND2X1 U38755 ( .A(n41945), .B(n61705), .Y(n38418) );
  NOR2X1 U38756 ( .A(n38420), .B(n38421), .Y(n38419) );
  AND2X1 U38757 ( .A(n62584), .B(n38442), .Y(n38420) );
  AND2X1 U38758 ( .A(n42114), .B(n62322), .Y(n38421) );
  NOR2X1 U38759 ( .A(n39145), .B(n38423), .Y(n38422) );
  INVX1 U38760 ( .A(n38422), .Y(n70459) );
  AND2X1 U38761 ( .A(n69935), .B(n69934), .Y(n38423) );
  NOR2X1 U38762 ( .A(n68592), .B(n68591), .Y(n38424) );
  NOR2X1 U38763 ( .A(n38426), .B(n38427), .Y(n38425) );
  INVX1 U38764 ( .A(n38425), .Y(n63284) );
  OR2X1 U38765 ( .A(n63277), .B(n63276), .Y(n38426) );
  AND2X1 U38766 ( .A(n63279), .B(n63278), .Y(n38427) );
  OR2X1 U38767 ( .A(n38428), .B(n37383), .Y(n65280) );
  NAND2X1 U38768 ( .A(n41612), .B(n64942), .Y(n38428) );
  NOR2X1 U38769 ( .A(n38430), .B(n38431), .Y(n38429) );
  AND2X1 U38770 ( .A(n61878), .B(n61879), .Y(n38430) );
  AND2X1 U38771 ( .A(n41951), .B(n61880), .Y(n38431) );
  AND2X1 U38772 ( .A(n62430), .B(n62429), .Y(n38432) );
  OR2X1 U38773 ( .A(n38433), .B(n38434), .Y(n71662) );
  AND2X1 U38774 ( .A(n71214), .B(n39629), .Y(n38433) );
  AND2X1 U38775 ( .A(n71213), .B(n71212), .Y(n38434) );
  XNOR2X1 U38776 ( .A(n71150), .B(n38145), .Y(n38435) );
  AND2X1 U38777 ( .A(n43538), .B(n68265), .Y(n68262) );
  AND2X1 U38778 ( .A(n63732), .B(n63733), .Y(n63734) );
  OR2X1 U38779 ( .A(n38436), .B(n38437), .Y(n69947) );
  OR2X1 U38780 ( .A(n69638), .B(n69637), .Y(n38436) );
  AND2X1 U38781 ( .A(n69640), .B(n39306), .Y(n38437) );
  AND2X1 U38782 ( .A(n43676), .B(n71116), .Y(n38438) );
  OR2X1 U38783 ( .A(n72040), .B(n43562), .Y(n72042) );
  OR2X1 U38784 ( .A(n38439), .B(n38440), .Y(n61674) );
  AND2X1 U38785 ( .A(n61810), .B(n61670), .Y(n38439) );
  AND2X1 U38786 ( .A(n41861), .B(n61672), .Y(n38440) );
  INVX1 U38787 ( .A(n40401), .Y(n38441) );
  OR2X1 U38788 ( .A(n38755), .B(n38756), .Y(n38442) );
  NAND2X1 U38789 ( .A(n60256), .B(n38961), .Y(n38443) );
  AND2X1 U38790 ( .A(n59682), .B(n59681), .Y(n38444) );
  NOR2X1 U38791 ( .A(n38446), .B(n38447), .Y(n38445) );
  INVX1 U38792 ( .A(n38445), .Y(n61666) );
  AND2X1 U38793 ( .A(n61815), .B(n61662), .Y(n38446) );
  AND2X1 U38794 ( .A(n61814), .B(n61664), .Y(n38447) );
  OR2X1 U38795 ( .A(n38448), .B(n38449), .Y(n66485) );
  AND2X1 U38796 ( .A(n66474), .B(n66014), .Y(n38448) );
  AND2X1 U38797 ( .A(n40781), .B(n66020), .Y(n38449) );
  NAND2X1 U38798 ( .A(n38676), .B(n41553), .Y(n38450) );
  OR2X1 U38799 ( .A(n38451), .B(n38452), .Y(n63165) );
  AND2X1 U38800 ( .A(n63155), .B(n63161), .Y(n38451) );
  AND2X1 U38801 ( .A(n63160), .B(n63159), .Y(n38452) );
  OR2X1 U38802 ( .A(n43657), .B(n68517), .Y(n68885) );
  NOR2X1 U38803 ( .A(n38454), .B(n38455), .Y(n38453) );
  AND2X1 U38804 ( .A(n61545), .B(n39409), .Y(n38454) );
  AND2X1 U38805 ( .A(n41931), .B(n61546), .Y(n38455) );
  OR2X1 U38806 ( .A(n38888), .B(n66293), .Y(n66626) );
  OR2X1 U38807 ( .A(n40358), .B(n40359), .Y(n38456) );
  OR2X1 U38808 ( .A(n71778), .B(n43663), .Y(n71779) );
  OR2X1 U38809 ( .A(n65288), .B(n38457), .Y(n66018) );
  NAND2X1 U38810 ( .A(n38458), .B(n65292), .Y(n38457) );
  OR2X1 U38811 ( .A(n41037), .B(n65289), .Y(n38458) );
  INVX1 U38812 ( .A(n63551), .Y(n38459) );
  NOR2X1 U38813 ( .A(n66026), .B(n38463), .Y(n38460) );
  OR2X1 U38814 ( .A(n38460), .B(n38461), .Y(n66034) );
  AND2X1 U38815 ( .A(n38462), .B(n66028), .Y(n38461) );
  INVX1 U38816 ( .A(n66030), .Y(n38462) );
  OR2X1 U38817 ( .A(n66030), .B(n66027), .Y(n38463) );
  INVX1 U38818 ( .A(n51983), .Y(n38464) );
  AND2X1 U38819 ( .A(n62482), .B(n62481), .Y(n38465) );
  AND2X1 U38820 ( .A(n66272), .B(n66273), .Y(n38466) );
  OR2X1 U38821 ( .A(n38467), .B(n38468), .Y(n60448) );
  AND2X1 U38822 ( .A(n60376), .B(n60377), .Y(n38467) );
  NOR2X1 U38823 ( .A(n39711), .B(n39712), .Y(n38468) );
  OR2X1 U38824 ( .A(n38469), .B(n38470), .Y(n64345) );
  AND2X1 U38825 ( .A(n41513), .B(n64221), .Y(n38469) );
  AND2X1 U38826 ( .A(n64229), .B(n64228), .Y(n38470) );
  AND2X1 U38827 ( .A(n59201), .B(n44071), .Y(n38471) );
  OR2X1 U38828 ( .A(n39751), .B(n39752), .Y(n38472) );
  INVX1 U38829 ( .A(n45176), .Y(n38473) );
  OR2X1 U38830 ( .A(n38474), .B(n38475), .Y(n61731) );
  AND2X1 U38831 ( .A(n61768), .B(n61728), .Y(n38474) );
  NOR2X1 U38832 ( .A(n39406), .B(n39407), .Y(n38475) );
  AND2X1 U38833 ( .A(n65992), .B(n65991), .Y(n38476) );
  NAND2X1 U38834 ( .A(n61269), .B(n38480), .Y(n38477) );
  AND2X1 U38835 ( .A(n38477), .B(n38478), .Y(n61274) );
  OR2X1 U38836 ( .A(n38479), .B(n61273), .Y(n38478) );
  INVX1 U38837 ( .A(n62522), .Y(n38479) );
  AND2X1 U38838 ( .A(n61268), .B(n62522), .Y(n38480) );
  AND2X1 U38839 ( .A(n68339), .B(n68089), .Y(n38481) );
  OR2X1 U38840 ( .A(n38482), .B(n38483), .Y(n59819) );
  AND2X1 U38841 ( .A(n59782), .B(n59629), .Y(n38482) );
  AND2X1 U38842 ( .A(n41828), .B(n59631), .Y(n38483) );
  AND2X1 U38843 ( .A(n65533), .B(n65532), .Y(n38484) );
  AND2X1 U38844 ( .A(n59129), .B(n36722), .Y(n38485) );
  NOR2X1 U38845 ( .A(n38487), .B(n38488), .Y(n38486) );
  AND2X1 U38846 ( .A(n60171), .B(n60172), .Y(n38487) );
  AND2X1 U38847 ( .A(n60174), .B(n60173), .Y(n38488) );
  OR2X1 U38848 ( .A(n65931), .B(n41398), .Y(n38489) );
  AND2X1 U38849 ( .A(n65933), .B(n43659), .Y(n38490) );
  OR2X1 U38850 ( .A(n41533), .B(n41534), .Y(n38491) );
  INVX1 U38851 ( .A(n42875), .Y(n38492) );
  AND2X1 U38852 ( .A(n62909), .B(n48108), .Y(n38493) );
  OR2X1 U38853 ( .A(n38495), .B(n38494), .Y(n65086) );
  INVX1 U38854 ( .A(n65039), .Y(n38494) );
  AND2X1 U38855 ( .A(n64767), .B(n65413), .Y(n38495) );
  AND2X1 U38856 ( .A(n38496), .B(n62338), .Y(n38498) );
  INVX1 U38857 ( .A(n40315), .Y(n38496) );
  INVX1 U38858 ( .A(n40316), .Y(n38497) );
  OR2X1 U38859 ( .A(n40315), .B(n40316), .Y(n38499) );
  INVX1 U38860 ( .A(n38499), .Y(n40314) );
  OR2X1 U38861 ( .A(n63562), .B(n43611), .Y(n38500) );
  INVX1 U38862 ( .A(n38802), .Y(n38501) );
  OR2X1 U38863 ( .A(n40650), .B(n40651), .Y(n38502) );
  OR2X1 U38864 ( .A(n40149), .B(n40150), .Y(n38503) );
  AND2X1 U38865 ( .A(n63810), .B(n63809), .Y(n38504) );
  INVX1 U38866 ( .A(n38504), .Y(n64427) );
  AND2X1 U38867 ( .A(n59534), .B(n59572), .Y(n38505) );
  OR2X1 U38868 ( .A(n38506), .B(n38507), .Y(n64419) );
  INVX1 U38869 ( .A(n64426), .Y(n38506) );
  AND2X1 U38870 ( .A(n39207), .B(n64120), .Y(n38507) );
  AND2X1 U38871 ( .A(n61041), .B(n61040), .Y(n38508) );
  NAND2X1 U38872 ( .A(n63987), .B(n38512), .Y(n38509) );
  AND2X1 U38873 ( .A(n38509), .B(n38510), .Y(n64588) );
  OR2X1 U38874 ( .A(n38511), .B(n63985), .Y(n38510) );
  INVX1 U38875 ( .A(n63986), .Y(n38511) );
  AND2X1 U38876 ( .A(n63720), .B(n63986), .Y(n38512) );
  OR2X1 U38877 ( .A(n38513), .B(n37375), .Y(n66026) );
  AND2X1 U38878 ( .A(n66025), .B(n41313), .Y(n38513) );
  NOR2X1 U38879 ( .A(n43470), .B(n43519), .Y(n38514) );
  INVX1 U38880 ( .A(n38514), .Y(n63226) );
  AND2X1 U38881 ( .A(n65268), .B(n41558), .Y(n38515) );
  NOR2X1 U38882 ( .A(n60641), .B(n60640), .Y(n38516) );
  NOR2X1 U38883 ( .A(n60641), .B(n60640), .Y(n38517) );
  AND2X1 U38884 ( .A(n38493), .B(n38636), .Y(n38518) );
  AND2X1 U38885 ( .A(n62141), .B(n62115), .Y(n38520) );
  AND2X1 U38886 ( .A(n42090), .B(n62117), .Y(n38521) );
  NOR2X1 U38887 ( .A(n39471), .B(n36785), .Y(n38522) );
  AND2X1 U38888 ( .A(n64030), .B(n38523), .Y(n63748) );
  INVX1 U38889 ( .A(n63746), .Y(n38523) );
  NOR2X1 U38890 ( .A(n40321), .B(n40322), .Y(n38524) );
  AND2X1 U38891 ( .A(n38525), .B(n38526), .Y(n41025) );
  NAND2X1 U38892 ( .A(n68507), .B(n68508), .Y(n38525) );
  NAND2X1 U38893 ( .A(n39084), .B(n68509), .Y(n38526) );
  NAND2X1 U38894 ( .A(n38652), .B(n62460), .Y(n38527) );
  INVX1 U38895 ( .A(n48361), .Y(n38528) );
  AND2X1 U38896 ( .A(n59467), .B(n59469), .Y(n38530) );
  NOR2X1 U38897 ( .A(n38726), .B(n38727), .Y(n38531) );
  OR2X1 U38898 ( .A(n38532), .B(n38533), .Y(n61725) );
  AND2X1 U38899 ( .A(n61721), .B(n61722), .Y(n38532) );
  AND2X1 U38900 ( .A(n41995), .B(n61723), .Y(n38533) );
  INVX1 U38901 ( .A(n47675), .Y(n38534) );
  OR2X1 U38902 ( .A(n38535), .B(n38536), .Y(n68868) );
  OR2X1 U38903 ( .A(n69547), .B(n68833), .Y(n38535) );
  NOR2X1 U38904 ( .A(n40215), .B(n40214), .Y(n38536) );
  INVX1 U38905 ( .A(n58469), .Y(n38537) );
  OR2X1 U38906 ( .A(n37364), .B(n38601), .Y(n38538) );
  NAND2X1 U38907 ( .A(n38538), .B(n38539), .Y(n70820) );
  AND2X1 U38908 ( .A(n70783), .B(n38540), .Y(n38539) );
  INVX1 U38909 ( .A(n40213), .Y(n38540) );
  OR2X1 U38910 ( .A(n60948), .B(n60949), .Y(n63823) );
  AND2X1 U38911 ( .A(n63721), .B(n63722), .Y(n38541) );
  INVX1 U38912 ( .A(n38541), .Y(n63985) );
  OR2X1 U38913 ( .A(n38542), .B(n38543), .Y(n62491) );
  AND2X1 U38914 ( .A(n61216), .B(n61215), .Y(n38542) );
  NOR2X1 U38915 ( .A(n61217), .B(n38812), .Y(n38543) );
  AND2X1 U38916 ( .A(n68985), .B(n68984), .Y(n38544) );
  OR2X1 U38917 ( .A(n38545), .B(n38546), .Y(n63702) );
  AND2X1 U38918 ( .A(n63423), .B(n63424), .Y(n38545) );
  AND2X1 U38919 ( .A(n42106), .B(n63426), .Y(n38546) );
  OR2X1 U38920 ( .A(n63598), .B(n42842), .Y(n63604) );
  AND2X1 U38921 ( .A(n63729), .B(n63730), .Y(n38547) );
  OR2X1 U38922 ( .A(n38548), .B(n38549), .Y(n60451) );
  AND2X1 U38923 ( .A(n60494), .B(n60495), .Y(n38548) );
  AND2X1 U38924 ( .A(n41855), .B(n60367), .Y(n38549) );
  OR2X1 U38925 ( .A(n59960), .B(n59961), .Y(n59964) );
  XOR2X1 U38926 ( .A(n71687), .B(n71782), .Y(n71695) );
  OR2X1 U38927 ( .A(n60618), .B(n60619), .Y(n60930) );
  OR2X1 U38928 ( .A(n38550), .B(n38551), .Y(n66832) );
  AND2X1 U38929 ( .A(n66315), .B(n66314), .Y(n38550) );
  OR2X1 U38930 ( .A(n66313), .B(n66837), .Y(n38551) );
  AND2X1 U38931 ( .A(n68572), .B(n43626), .Y(n38552) );
  INVX1 U38932 ( .A(n38552), .Y(n68571) );
  OR2X1 U38933 ( .A(n38553), .B(n38554), .Y(n70206) );
  NAND2X1 U38934 ( .A(n39103), .B(n39104), .Y(n38553) );
  AND2X1 U38935 ( .A(n69583), .B(n69582), .Y(n38554) );
  OR2X1 U38936 ( .A(n38555), .B(n70460), .Y(n70770) );
  INVX1 U38937 ( .A(n43665), .Y(n38555) );
  AND2X1 U38938 ( .A(n65143), .B(n65142), .Y(n38556) );
  AND2X1 U38939 ( .A(n70472), .B(n70161), .Y(n38557) );
  XNOR2X1 U38940 ( .A(n41010), .B(n40705), .Y(n38558) );
  OR2X1 U38941 ( .A(n38559), .B(n38560), .Y(n64587) );
  INVX1 U38942 ( .A(n42083), .Y(n38559) );
  NOR2X1 U38943 ( .A(n39382), .B(n39383), .Y(n38560) );
  INVX1 U38944 ( .A(n40503), .Y(n38561) );
  OR2X1 U38945 ( .A(n38563), .B(n38562), .Y(n65479) );
  INVX1 U38946 ( .A(n65645), .Y(n38562) );
  OR2X1 U38947 ( .A(n41349), .B(n41576), .Y(n38563) );
  OR2X1 U38948 ( .A(n43710), .B(n71126), .Y(n72107) );
  AND2X1 U38949 ( .A(n64365), .B(n64364), .Y(n38564) );
  AND2X1 U38950 ( .A(n63180), .B(n63179), .Y(n38565) );
  OR2X1 U38951 ( .A(n39141), .B(n39142), .Y(n38566) );
  OR2X1 U38952 ( .A(n38567), .B(n38568), .Y(n63681) );
  AND2X1 U38953 ( .A(n63387), .B(n63388), .Y(n38567) );
  AND2X1 U38954 ( .A(n42107), .B(n63391), .Y(n38568) );
  INVX1 U38955 ( .A(n60148), .Y(n38569) );
  NAND2X1 U38956 ( .A(n38570), .B(n60147), .Y(n60150) );
  NOR2X1 U38957 ( .A(n38569), .B(n36749), .Y(n38570) );
  NAND2X1 U38958 ( .A(n62476), .B(n62475), .Y(n38571) );
  OR2X1 U38959 ( .A(n48109), .B(n36820), .Y(n38572) );
  NOR2X1 U38960 ( .A(n48210), .B(n42854), .Y(n38573) );
  OR2X1 U38961 ( .A(n38574), .B(n38575), .Y(n67550) );
  OR2X1 U38962 ( .A(n67547), .B(n67546), .Y(n38574) );
  AND2X1 U38963 ( .A(n43581), .B(n67548), .Y(n38575) );
  AND2X1 U38964 ( .A(n63978), .B(n63979), .Y(n38576) );
  INVX1 U38965 ( .A(n48381), .Y(n38577) );
  OR2X1 U38966 ( .A(n38578), .B(n38579), .Y(n64638) );
  AND2X1 U38967 ( .A(n64640), .B(n64641), .Y(n38578) );
  AND2X1 U38968 ( .A(n42040), .B(n64314), .Y(n38579) );
  INVX1 U38969 ( .A(n38628), .Y(n38580) );
  OR2X1 U38970 ( .A(n58469), .B(n42783), .Y(n46207) );
  OR2X1 U38971 ( .A(n38581), .B(n36724), .Y(n40707) );
  OR2X1 U38972 ( .A(n69523), .B(n69208), .Y(n38581) );
  INVX1 U38973 ( .A(n43808), .Y(n38582) );
  NOR2X1 U38974 ( .A(n38585), .B(n38584), .Y(n38583) );
  INVX1 U38975 ( .A(n38583), .Y(n64946) );
  INVX1 U38976 ( .A(n64960), .Y(n38584) );
  OR2X1 U38977 ( .A(n41572), .B(n41579), .Y(n38585) );
  OR2X1 U38978 ( .A(n43756), .B(n38586), .Y(n62655) );
  INVX1 U38979 ( .A(n42720), .Y(n38586) );
  OR2X1 U38980 ( .A(n38587), .B(n38588), .Y(n72686) );
  AND2X1 U38981 ( .A(n38399), .B(n43513), .Y(n38587) );
  AND2X1 U38982 ( .A(n71731), .B(n71732), .Y(n38588) );
  INVX1 U38983 ( .A(n41927), .Y(n38589) );
  AND2X1 U38984 ( .A(n62181), .B(n62052), .Y(n38590) );
  OR2X1 U38985 ( .A(n70787), .B(n70782), .Y(n38591) );
  NAND2X1 U38986 ( .A(n36783), .B(n63825), .Y(n38592) );
  OR2X1 U38987 ( .A(n36777), .B(n38593), .Y(n64150) );
  AND2X1 U38988 ( .A(n63527), .B(n63526), .Y(n38593) );
  AND2X1 U38989 ( .A(n36564), .B(n38596), .Y(n38594) );
  NOR2X1 U38990 ( .A(n38594), .B(n38595), .Y(n39269) );
  AND2X1 U38991 ( .A(n70788), .B(n43696), .Y(n38596) );
  AND2X1 U38992 ( .A(n38597), .B(n67515), .Y(n67832) );
  OR2X1 U38993 ( .A(n67166), .B(n67511), .Y(n38597) );
  XNOR2X1 U38994 ( .A(n61297), .B(n62372), .Y(n38598) );
  INVX1 U38995 ( .A(n47624), .Y(n38599) );
  AND2X1 U38996 ( .A(n65111), .B(n65110), .Y(n38600) );
  INVX1 U38997 ( .A(n38600), .Y(n65696) );
  OR2X1 U38998 ( .A(n37364), .B(n38601), .Y(n70785) );
  OR2X1 U38999 ( .A(n41339), .B(n70207), .Y(n38601) );
  INVX1 U39000 ( .A(n45317), .Y(n38602) );
  OR2X1 U39001 ( .A(n38603), .B(n67018), .Y(n67022) );
  INVX1 U39002 ( .A(n67329), .Y(n38603) );
  OR2X1 U39003 ( .A(n58469), .B(n40510), .Y(n46206) );
  AND2X1 U39004 ( .A(n46019), .B(n42671), .Y(n38604) );
  AND2X1 U39005 ( .A(n36625), .B(n69243), .Y(n38605) );
  NOR2X1 U39006 ( .A(n38607), .B(n38608), .Y(n38606) );
  AND2X1 U39007 ( .A(n43536), .B(n66284), .Y(n38607) );
  AND2X1 U39008 ( .A(n66287), .B(n66286), .Y(n38608) );
  INVX1 U39009 ( .A(n36608), .Y(n38609) );
  NOR2X1 U39010 ( .A(n63562), .B(n43611), .Y(n38610) );
  INVX1 U39011 ( .A(n43747), .Y(n38611) );
  OR2X1 U39012 ( .A(n40550), .B(n40551), .Y(n38612) );
  OR2X1 U39013 ( .A(n68264), .B(n39927), .Y(n67651) );
  AND2X1 U39014 ( .A(n40390), .B(n61192), .Y(n60956) );
  OR2X1 U39015 ( .A(n38613), .B(n36757), .Y(n59168) );
  OR2X1 U39016 ( .A(n59127), .B(n59126), .Y(n38613) );
  NOR2X1 U39017 ( .A(n38615), .B(n38616), .Y(n38614) );
  OR2X1 U39018 ( .A(n45866), .B(n45865), .Y(n38615) );
  AND2X1 U39019 ( .A(n40490), .B(n45916), .Y(n38616) );
  AND2X1 U39020 ( .A(n69168), .B(n69167), .Y(n38617) );
  OR2X1 U39021 ( .A(n40068), .B(n40069), .Y(n38618) );
  XOR2X1 U39022 ( .A(n63578), .B(n36777), .Y(n38619) );
  OR2X1 U39023 ( .A(n38621), .B(n38620), .Y(n64844) );
  INVX1 U39024 ( .A(n64357), .Y(n38620) );
  OR2X1 U39025 ( .A(n64353), .B(n64352), .Y(n38621) );
  NAND2X1 U39026 ( .A(n65715), .B(n40987), .Y(n38622) );
  OR2X1 U39027 ( .A(n39027), .B(n39028), .Y(n38623) );
  NAND2X1 U39028 ( .A(n68557), .B(n38626), .Y(n38624) );
  NAND2X1 U39029 ( .A(n38624), .B(n38625), .Y(n40167) );
  OR2X1 U39030 ( .A(n39747), .B(n68892), .Y(n38625) );
  AND2X1 U39031 ( .A(n43670), .B(n43670), .Y(n38626) );
  OR2X1 U39032 ( .A(n37097), .B(n40479), .Y(n38627) );
  OR2X1 U39033 ( .A(n42881), .B(n40479), .Y(n49665) );
  OR2X1 U39034 ( .A(n40456), .B(n38628), .Y(n72721) );
  XOR2X1 U39035 ( .A(n36631), .B(n72104), .Y(n38628) );
  NOR2X1 U39036 ( .A(n61725), .B(n61724), .Y(n39404) );
  XOR2X1 U39037 ( .A(n39655), .B(n70453), .Y(n69916) );
  NAND2X1 U39038 ( .A(n38631), .B(n38630), .Y(n38629) );
  INVX1 U39039 ( .A(n38629), .Y(n62837) );
  INVX1 U39040 ( .A(n62838), .Y(n38630) );
  OR2X1 U39041 ( .A(n41269), .B(n41270), .Y(n38631) );
  OR2X1 U39042 ( .A(n38632), .B(n38633), .Y(n49401) );
  NAND2X1 U39043 ( .A(n42472), .B(n42473), .Y(n38632) );
  AND2X1 U39044 ( .A(n2767), .B(n57613), .Y(n38633) );
  OR2X1 U39045 ( .A(n38634), .B(n36746), .Y(n46214) );
  OR2X1 U39046 ( .A(n46213), .B(n46212), .Y(n38634) );
  OR2X1 U39047 ( .A(n38977), .B(n38978), .Y(n38635) );
  INVX1 U39048 ( .A(n38700), .Y(n38636) );
  XNOR2X1 U39049 ( .A(n50720), .B(opcode_opcode_w[21]), .Y(n38637) );
  INVX1 U39050 ( .A(n38637), .Y(n45267) );
  NOR2X1 U39051 ( .A(n39345), .B(n39346), .Y(n38638) );
  NAND2X1 U39052 ( .A(n63651), .B(n38639), .Y(n63744) );
  NOR2X1 U39053 ( .A(n63648), .B(n63647), .Y(n38639) );
  OR2X1 U39054 ( .A(n38640), .B(n38641), .Y(n66761) );
  AND2X1 U39055 ( .A(n66359), .B(n66358), .Y(n38640) );
  AND2X1 U39056 ( .A(n66364), .B(n66363), .Y(n38641) );
  OR2X1 U39057 ( .A(n48193), .B(n48192), .Y(n38642) );
  OR2X1 U39058 ( .A(n48223), .B(n48222), .Y(n38643) );
  OR2X1 U39059 ( .A(n38644), .B(n42720), .Y(n63826) );
  NAND2X1 U39060 ( .A(n36783), .B(n63825), .Y(n38644) );
  OR2X1 U39061 ( .A(n46006), .B(n46206), .Y(n49624) );
  NOR2X1 U39062 ( .A(n38646), .B(n38647), .Y(n38645) );
  AND2X1 U39063 ( .A(n60887), .B(n60886), .Y(n38646) );
  AND2X1 U39064 ( .A(n60891), .B(n60890), .Y(n38647) );
  AND2X1 U39065 ( .A(n38648), .B(n38649), .Y(n45618) );
  AND2X1 U39066 ( .A(n2956), .B(n45614), .Y(n38648) );
  AND2X1 U39067 ( .A(n45615), .B(n45176), .Y(n38649) );
  OR2X1 U39068 ( .A(n38650), .B(n38651), .Y(n63157) );
  INVX1 U39069 ( .A(n62422), .Y(n38650) );
  OR2X1 U39070 ( .A(n39422), .B(n62871), .Y(n38651) );
  NOR2X1 U39071 ( .A(n38653), .B(n38654), .Y(n38652) );
  INVX1 U39072 ( .A(n38652), .Y(n63190) );
  AND2X1 U39073 ( .A(writeback_exec_value_w[2]), .B(n43025), .Y(n38653) );
  AND2X1 U39074 ( .A(n47707), .B(n62907), .Y(n38654) );
  OR2X1 U39075 ( .A(n39345), .B(n39346), .Y(n38655) );
  INVX1 U39076 ( .A(n38815), .Y(n38656) );
  OR2X1 U39077 ( .A(n38657), .B(n38816), .Y(n61890) );
  NAND2X1 U39078 ( .A(n38656), .B(n61889), .Y(n38657) );
  XNOR2X1 U39079 ( .A(n71439), .B(n38658), .Y(n71689) );
  XOR2X1 U39080 ( .A(n71660), .B(n71399), .Y(n38658) );
  AND2X1 U39081 ( .A(opcode_opcode_w[23]), .B(n42750), .Y(n38659) );
  NOR2X1 U39082 ( .A(n63302), .B(n37407), .Y(n38660) );
  OR2X1 U39083 ( .A(n60525), .B(n37403), .Y(n60526) );
  OR2X1 U39084 ( .A(n42329), .B(n42328), .Y(n38661) );
  OR2X1 U39085 ( .A(n42329), .B(n42328), .Y(n38662) );
  XOR2X1 U39086 ( .A(n63629), .B(n63022), .Y(n63642) );
  XNOR2X1 U39087 ( .A(opcode_opcode_w[24]), .B(n45299), .Y(n38663) );
  XNOR2X1 U39088 ( .A(n41284), .B(n63366), .Y(n38664) );
  NOR2X1 U39089 ( .A(n40412), .B(n40413), .Y(n38665) );
  OR2X1 U39090 ( .A(n38666), .B(n42622), .Y(n49378) );
  AND2X1 U39091 ( .A(n38668), .B(n38667), .Y(n63647) );
  INVX1 U39092 ( .A(n63646), .Y(n38667) );
  OR2X1 U39093 ( .A(n63645), .B(n63644), .Y(n38668) );
  AND2X1 U39094 ( .A(n64330), .B(n64329), .Y(n38669) );
  OR2X1 U39095 ( .A(n65019), .B(n37408), .Y(n65011) );
  INVX1 U39096 ( .A(n38829), .Y(n38670) );
  OR2X1 U39097 ( .A(n38671), .B(n38830), .Y(n62117) );
  NAND2X1 U39098 ( .A(n38670), .B(n62116), .Y(n38671) );
  OR2X1 U39099 ( .A(n39480), .B(n39481), .Y(n38672) );
  INVX1 U39100 ( .A(n64811), .Y(n38673) );
  AND2X1 U39101 ( .A(n39207), .B(n64120), .Y(n38674) );
  AND2X1 U39102 ( .A(n69926), .B(n38208), .Y(n39748) );
  NOR2X1 U39103 ( .A(n40109), .B(n40110), .Y(n38675) );
  XNOR2X1 U39104 ( .A(n62514), .B(n41561), .Y(n38676) );
  OR2X1 U39105 ( .A(n46577), .B(n38677), .Y(n46396) );
  OR2X1 U39106 ( .A(n46726), .B(n38678), .Y(n38677) );
  AND2X1 U39107 ( .A(n66107), .B(n66415), .Y(n38679) );
  XOR2X1 U39108 ( .A(n64317), .B(n38681), .Y(n38680) );
  INVX1 U39109 ( .A(n38680), .Y(n64322) );
  XOR2X1 U39110 ( .A(n64318), .B(n64669), .Y(n38681) );
  AND2X1 U39111 ( .A(n64061), .B(n38682), .Y(n64063) );
  AND2X1 U39112 ( .A(n64150), .B(n64448), .Y(n38682) );
  AND2X1 U39113 ( .A(n71801), .B(n71800), .Y(n38683) );
  INVX1 U39114 ( .A(n38683), .Y(n72041) );
  NOR2X1 U39115 ( .A(n46326), .B(n42768), .Y(n42821) );
  NOR2X1 U39116 ( .A(n38685), .B(n38686), .Y(n38684) );
  AND2X1 U39117 ( .A(n61043), .B(n61042), .Y(n38685) );
  AND2X1 U39118 ( .A(n61047), .B(n61046), .Y(n38686) );
  OR2X1 U39119 ( .A(n39915), .B(n39916), .Y(n38687) );
  NOR2X1 U39120 ( .A(n40239), .B(n40240), .Y(n38688) );
  OR2X1 U39121 ( .A(n42887), .B(n38689), .Y(n46362) );
  AND2X1 U39122 ( .A(n46361), .B(n46360), .Y(n38689) );
  AND2X1 U39123 ( .A(n46585), .B(n46584), .Y(n38690) );
  AND2X1 U39124 ( .A(n40392), .B(n39844), .Y(n38691) );
  INVX1 U39125 ( .A(n38691), .Y(n62929) );
  OR2X1 U39126 ( .A(n40014), .B(n38432), .Y(n62971) );
  OR2X1 U39127 ( .A(n40126), .B(n40127), .Y(n38692) );
  AND2X1 U39128 ( .A(n61000), .B(n60999), .Y(n38693) );
  XNOR2X1 U39129 ( .A(n68549), .B(n41072), .Y(n38694) );
  OR2X1 U39130 ( .A(n39618), .B(n39619), .Y(n38695) );
  OR2X1 U39131 ( .A(n38750), .B(n38749), .Y(n38696) );
  AND2X1 U39132 ( .A(n64495), .B(n64497), .Y(n38697) );
  NOR2X1 U39133 ( .A(n64389), .B(n38698), .Y(n40133) );
  NAND2X1 U39134 ( .A(n38699), .B(n64392), .Y(n38698) );
  OR2X1 U39135 ( .A(n39836), .B(n64388), .Y(n38699) );
  OR2X1 U39136 ( .A(n62455), .B(n38700), .Y(n40228) );
  AND2X1 U39137 ( .A(n42801), .B(n62453), .Y(n38700) );
  INVX1 U39138 ( .A(n39645), .Y(n38701) );
  OR2X1 U39139 ( .A(n38702), .B(n38703), .Y(n62988) );
  AND2X1 U39140 ( .A(n63275), .B(n62981), .Y(n38702) );
  OR2X1 U39141 ( .A(n63274), .B(n63280), .Y(n38703) );
  NOR2X1 U39142 ( .A(n62836), .B(n38704), .Y(n39782) );
  NAND2X1 U39143 ( .A(n38629), .B(n62840), .Y(n38704) );
  XNOR2X1 U39144 ( .A(n38706), .B(n59462), .Y(n38705) );
  INVX1 U39145 ( .A(n38705), .Y(n59515) );
  XOR2X1 U39146 ( .A(n59461), .B(n59460), .Y(n38706) );
  OR2X1 U39147 ( .A(n62538), .B(n62539), .Y(n62536) );
  XNOR2X1 U39148 ( .A(n38707), .B(n61126), .Y(n61235) );
  XOR2X1 U39149 ( .A(n61128), .B(n36755), .Y(n38707) );
  INVX1 U39150 ( .A(n38944), .Y(n38708) );
  INVX1 U39151 ( .A(n38944), .Y(n38709) );
  INVX1 U39152 ( .A(n38944), .Y(n38710) );
  INVX1 U39153 ( .A(n42819), .Y(n38711) );
  INVX1 U39154 ( .A(n42819), .Y(n38712) );
  NOR2X1 U39155 ( .A(n38714), .B(n38713), .Y(n41637) );
  INVX1 U39156 ( .A(n69633), .Y(n38713) );
  AND2X1 U39157 ( .A(n69488), .B(n69487), .Y(n38714) );
  OR2X1 U39158 ( .A(n38715), .B(n38716), .Y(n45894) );
  OR2X1 U39159 ( .A(n39809), .B(n42881), .Y(n38715) );
  INVX1 U39160 ( .A(n42885), .Y(n38717) );
  OR2X1 U39161 ( .A(n38718), .B(n38719), .Y(n45923) );
  AND2X1 U39162 ( .A(n45921), .B(n42149), .Y(n38718) );
  NOR2X1 U39163 ( .A(n38819), .B(n38820), .Y(n38719) );
  INVX1 U39164 ( .A(n63141), .Y(n38720) );
  OR2X1 U39165 ( .A(n38722), .B(n38723), .Y(n59891) );
  OR2X1 U39166 ( .A(n60942), .B(n59889), .Y(n38722) );
  OR2X1 U39167 ( .A(n62458), .B(n39192), .Y(n38723) );
  AND2X1 U39168 ( .A(n39552), .B(n60721), .Y(n38724) );
  XNOR2X1 U39169 ( .A(n67628), .B(n36705), .Y(n38725) );
  INVX1 U39170 ( .A(n42155), .Y(n38726) );
  AND2X1 U39171 ( .A(n42839), .B(n59420), .Y(n38727) );
  XOR2X1 U39172 ( .A(n59929), .B(n40663), .Y(n38728) );
  OR2X1 U39173 ( .A(n64063), .B(n38732), .Y(n38729) );
  AND2X1 U39174 ( .A(n38729), .B(n38730), .Y(n65025) );
  OR2X1 U39175 ( .A(n38731), .B(n64729), .Y(n38730) );
  INVX1 U39176 ( .A(n64732), .Y(n38731) );
  OR2X1 U39177 ( .A(n64062), .B(n38731), .Y(n38732) );
  OR2X1 U39178 ( .A(n59381), .B(n38733), .Y(n59384) );
  NAND2X1 U39179 ( .A(n59382), .B(n59383), .Y(n38733) );
  AND2X1 U39180 ( .A(n38734), .B(n38735), .Y(n71776) );
  OR2X1 U39181 ( .A(n43654), .B(n71778), .Y(n38734) );
  AND2X1 U39182 ( .A(n71774), .B(n41392), .Y(n38735) );
  NOR2X1 U39183 ( .A(n61731), .B(n61730), .Y(n40102) );
  AND2X1 U39184 ( .A(n67436), .B(n67437), .Y(n38736) );
  OR2X1 U39185 ( .A(n38737), .B(n38738), .Y(n49403) );
  OR2X1 U39186 ( .A(n49397), .B(n49396), .Y(n38737) );
  OR2X1 U39187 ( .A(n49402), .B(n49401), .Y(n38738) );
  AND2X1 U39188 ( .A(n44994), .B(n42686), .Y(n38739) );
  AND2X1 U39189 ( .A(n40523), .B(n42772), .Y(n38740) );
  OR2X1 U39190 ( .A(n38741), .B(n38742), .Y(n63698) );
  AND2X1 U39191 ( .A(n43676), .B(n63419), .Y(n38741) );
  AND2X1 U39192 ( .A(n63422), .B(n63421), .Y(n38742) );
  OR2X1 U39193 ( .A(n49630), .B(n38743), .Y(n46227) );
  OR2X1 U39194 ( .A(n42793), .B(n42669), .Y(n48612) );
  OR2X1 U39195 ( .A(n46577), .B(n46726), .Y(n38745) );
  NOR2X1 U39196 ( .A(n38747), .B(n38748), .Y(n38746) );
  INVX1 U39197 ( .A(n38746), .Y(n61418) );
  AND2X1 U39198 ( .A(n39823), .B(n61415), .Y(n38747) );
  AND2X1 U39199 ( .A(n41965), .B(n61416), .Y(n38748) );
  OR2X1 U39200 ( .A(n38749), .B(n38750), .Y(n64812) );
  NOR2X1 U39201 ( .A(n39935), .B(n39934), .Y(n38749) );
  AND2X1 U39202 ( .A(n64461), .B(n64460), .Y(n38750) );
  OR2X1 U39203 ( .A(n62455), .B(n38751), .Y(n61193) );
  AND2X1 U39204 ( .A(n42803), .B(n59144), .Y(n38751) );
  NAND2X1 U39205 ( .A(n38947), .B(n42770), .Y(n38752) );
  OR2X1 U39206 ( .A(n38821), .B(n39770), .Y(n38753) );
  NOR2X1 U39207 ( .A(n38755), .B(n38756), .Y(n38754) );
  AND2X1 U39208 ( .A(n62318), .B(n62319), .Y(n38755) );
  AND2X1 U39209 ( .A(n42108), .B(n62320), .Y(n38756) );
  NAND2X1 U39210 ( .A(n62915), .B(n38760), .Y(n38757) );
  NAND2X1 U39211 ( .A(n38757), .B(n38758), .Y(n39626) );
  OR2X1 U39212 ( .A(n38759), .B(n42802), .Y(n38758) );
  INVX1 U39213 ( .A(n38652), .Y(n38759) );
  AND2X1 U39214 ( .A(n62916), .B(n38652), .Y(n38760) );
  NOR2X1 U39215 ( .A(n38762), .B(n38763), .Y(n38761) );
  INVX1 U39216 ( .A(n38761), .Y(n61517) );
  AND2X1 U39217 ( .A(n61514), .B(n61515), .Y(n38762) );
  AND2X1 U39218 ( .A(n41837), .B(n61516), .Y(n38763) );
  NOR2X1 U39219 ( .A(n42738), .B(n48109), .Y(n38764) );
  XNOR2X1 U39220 ( .A(n59277), .B(n59725), .Y(n38765) );
  OR2X1 U39221 ( .A(n38766), .B(n38767), .Y(n70733) );
  OR2X1 U39222 ( .A(n70268), .B(n70267), .Y(n38766) );
  AND2X1 U39223 ( .A(n70271), .B(n70578), .Y(n38767) );
  OR2X1 U39224 ( .A(opcode_opcode_w[20]), .B(n38960), .Y(n38768) );
  NAND2X1 U39225 ( .A(n59225), .B(n38772), .Y(n38769) );
  AND2X1 U39226 ( .A(n38769), .B(n38770), .Y(n59681) );
  OR2X1 U39227 ( .A(n38771), .B(n59678), .Y(n38770) );
  INVX1 U39228 ( .A(n59680), .Y(n38771) );
  AND2X1 U39229 ( .A(n42816), .B(n59680), .Y(n38772) );
  AND2X1 U39230 ( .A(n63127), .B(n63128), .Y(n38773) );
  INVX1 U39231 ( .A(n38773), .Y(n63670) );
  OR2X1 U39232 ( .A(n38775), .B(n38774), .Y(n64321) );
  INVX1 U39233 ( .A(n64319), .Y(n38774) );
  OR2X1 U39234 ( .A(n41564), .B(n41606), .Y(n38775) );
  OR2X1 U39235 ( .A(n38907), .B(n38908), .Y(n38776) );
  OR2X1 U39236 ( .A(n42366), .B(n45271), .Y(n38777) );
  OR2X1 U39237 ( .A(n38778), .B(n38779), .Y(n61178) );
  OR2X1 U39238 ( .A(n47960), .B(n47959), .Y(n38778) );
  OR2X1 U39239 ( .A(n47984), .B(n47983), .Y(n38779) );
  AND2X1 U39240 ( .A(n63117), .B(n37382), .Y(n38780) );
  INVX1 U39241 ( .A(n38780), .Y(n63673) );
  AND2X1 U39242 ( .A(n65987), .B(n65875), .Y(n38781) );
  OR2X1 U39243 ( .A(n39936), .B(n39903), .Y(n38782) );
  OR2X1 U39244 ( .A(n39936), .B(n39903), .Y(n38783) );
  OR2X1 U39245 ( .A(n63015), .B(n63016), .Y(n63330) );
  NOR2X1 U39246 ( .A(n39339), .B(n39340), .Y(n38784) );
  OR2X1 U39247 ( .A(n38785), .B(n42689), .Y(n48186) );
  OR2X1 U39248 ( .A(n42728), .B(n42726), .Y(n38785) );
  OR2X1 U39249 ( .A(n38773), .B(n38786), .Y(n39223) );
  AND2X1 U39250 ( .A(n63669), .B(n43984), .Y(n38786) );
  NOR2X1 U39251 ( .A(n38787), .B(n38598), .Y(n41601) );
  NAND2X1 U39252 ( .A(n63033), .B(n63035), .Y(n38787) );
  AND2X1 U39253 ( .A(n68338), .B(n68341), .Y(n38788) );
  XNOR2X1 U39254 ( .A(n38789), .B(n38790), .Y(n67632) );
  INVX1 U39255 ( .A(n41300), .Y(n38789) );
  OR2X1 U39256 ( .A(n67874), .B(n40504), .Y(n38790) );
  AND2X1 U39257 ( .A(n59410), .B(n59407), .Y(n38791) );
  INVX1 U39258 ( .A(n38791), .Y(n59347) );
  AND2X1 U39259 ( .A(n64511), .B(n64510), .Y(n38792) );
  AND2X1 U39260 ( .A(n45311), .B(n45310), .Y(n38793) );
  INVX1 U39261 ( .A(n38793), .Y(n47706) );
  OR2X1 U39262 ( .A(n38794), .B(n38795), .Y(n65060) );
  AND2X1 U39263 ( .A(n64798), .B(n64414), .Y(n38794) );
  AND2X1 U39264 ( .A(n64416), .B(n64415), .Y(n38795) );
  OR2X1 U39265 ( .A(n40363), .B(n40364), .Y(n38796) );
  OR2X1 U39266 ( .A(n45255), .B(n38661), .Y(n45615) );
  OR2X1 U39267 ( .A(n38780), .B(n38797), .Y(n63674) );
  AND2X1 U39268 ( .A(n63672), .B(n43993), .Y(n38797) );
  OR2X1 U39269 ( .A(n40532), .B(n46007), .Y(n38798) );
  AND2X1 U39270 ( .A(n48157), .B(n48156), .Y(n38799) );
  OR2X1 U39271 ( .A(n38800), .B(n38801), .Y(n45525) );
  AND2X1 U39272 ( .A(n45523), .B(n38604), .Y(n38800) );
  AND2X1 U39273 ( .A(n45524), .B(n40499), .Y(n38801) );
  INVX1 U39274 ( .A(n58458), .Y(n38802) );
  NAND2X1 U39275 ( .A(n59464), .B(n59437), .Y(n38803) );
  AND2X1 U39276 ( .A(n48145), .B(n48144), .Y(n38804) );
  INVX1 U39277 ( .A(n42645), .Y(n38805) );
  NOR2X1 U39278 ( .A(n42808), .B(n42688), .Y(n38806) );
  OR2X1 U39279 ( .A(n38807), .B(n45619), .Y(n45610) );
  OR2X1 U39280 ( .A(n68089), .B(n68339), .Y(n68635) );
  NAND2X1 U39281 ( .A(n45276), .B(n45533), .Y(n38807) );
  NAND2X1 U39282 ( .A(n38179), .B(n38811), .Y(n38808) );
  AND2X1 U39283 ( .A(n38808), .B(n38809), .Y(n69302) );
  OR2X1 U39284 ( .A(n38810), .B(n69161), .Y(n38809) );
  INVX1 U39285 ( .A(n69301), .Y(n38810) );
  AND2X1 U39286 ( .A(n69159), .B(n69301), .Y(n38811) );
  AND2X1 U39287 ( .A(n40595), .B(n61218), .Y(n38812) );
  INVX1 U39288 ( .A(n38518), .Y(n38813) );
  NOR2X1 U39289 ( .A(n38815), .B(n38816), .Y(n38814) );
  INVX1 U39290 ( .A(n38814), .Y(n61888) );
  AND2X1 U39291 ( .A(n61885), .B(n61886), .Y(n38815) );
  AND2X1 U39292 ( .A(n41970), .B(n61887), .Y(n38816) );
  OR2X1 U39293 ( .A(n38817), .B(n38792), .Y(n64632) );
  AND2X1 U39294 ( .A(n64631), .B(n44018), .Y(n38817) );
  XOR2X1 U39295 ( .A(n36631), .B(n72104), .Y(n38818) );
  OR2X1 U39296 ( .A(n60916), .B(n60917), .Y(n60712) );
  OR2X1 U39297 ( .A(n46009), .B(n46526), .Y(n38819) );
  OR2X1 U39298 ( .A(n46577), .B(n37064), .Y(n38820) );
  INVX1 U39299 ( .A(n38848), .Y(n38821) );
  INVX1 U39300 ( .A(n38848), .Y(n38822) );
  INVX1 U39301 ( .A(n38848), .Y(n38823) );
  INVX1 U39302 ( .A(n49588), .Y(n38824) );
  INVX1 U39303 ( .A(n49588), .Y(n38825) );
  NAND2X1 U39304 ( .A(n42803), .B(n59144), .Y(n38827) );
  NOR2X1 U39305 ( .A(n38829), .B(n38830), .Y(n38828) );
  INVX1 U39306 ( .A(n38828), .Y(n62115) );
  AND2X1 U39307 ( .A(n62112), .B(n62113), .Y(n38829) );
  AND2X1 U39308 ( .A(n42080), .B(n62114), .Y(n38830) );
  OR2X1 U39309 ( .A(n58469), .B(n40866), .Y(n46372) );
  NOR2X1 U39310 ( .A(n42368), .B(n42369), .Y(n38831) );
  OR2X1 U39311 ( .A(n38832), .B(n38833), .Y(n62404) );
  AND2X1 U39312 ( .A(n36721), .B(n61233), .Y(n38832) );
  AND2X1 U39313 ( .A(n61237), .B(n61236), .Y(n38833) );
  OR2X1 U39314 ( .A(n38835), .B(n38834), .Y(n70720) );
  INVX1 U39315 ( .A(n71045), .Y(n38834) );
  AND2X1 U39316 ( .A(n71042), .B(n70718), .Y(n38835) );
  OR2X1 U39317 ( .A(n38836), .B(n38837), .Y(n62890) );
  AND2X1 U39318 ( .A(n40960), .B(n62885), .Y(n38836) );
  OR2X1 U39319 ( .A(n63290), .B(n63295), .Y(n38837) );
  OR2X1 U39320 ( .A(n38838), .B(n38839), .Y(n45916) );
  OR2X1 U39321 ( .A(n45891), .B(n45890), .Y(n38838) );
  OR2X1 U39322 ( .A(n45915), .B(n45914), .Y(n38839) );
  AND2X1 U39323 ( .A(n71645), .B(n71233), .Y(n38840) );
  INVX1 U39324 ( .A(n38840), .Y(n71663) );
  OR2X1 U39325 ( .A(n38841), .B(n37385), .Y(n67217) );
  AND2X1 U39326 ( .A(n66892), .B(n66891), .Y(n38841) );
  XNOR2X1 U39327 ( .A(n40710), .B(n68924), .Y(n38842) );
  INVX1 U39328 ( .A(n38842), .Y(n69207) );
  OR2X1 U39329 ( .A(n38843), .B(n37391), .Y(n65088) );
  OR2X1 U39330 ( .A(n64749), .B(n64748), .Y(n38843) );
  OR2X1 U39331 ( .A(n58820), .B(n42783), .Y(n46575) );
  INVX1 U39332 ( .A(n42894), .Y(n38844) );
  OR2X1 U39333 ( .A(n39231), .B(n39232), .Y(n38845) );
  NOR2X1 U39334 ( .A(n38807), .B(n45181), .Y(n38846) );
  NAND2X1 U39335 ( .A(n38847), .B(n45522), .Y(n39683) );
  NOR2X1 U39336 ( .A(n38414), .B(n45525), .Y(n38847) );
  NOR2X1 U39337 ( .A(n40516), .B(n42814), .Y(n38848) );
  NAND2X1 U39338 ( .A(n47164), .B(n38849), .Y(n42348) );
  NOR2X1 U39339 ( .A(n38850), .B(n47165), .Y(n38849) );
  OR2X1 U39340 ( .A(n47163), .B(n47162), .Y(n38850) );
  NOR2X1 U39341 ( .A(n63681), .B(n63682), .Y(n40330) );
  AND2X1 U39342 ( .A(n62374), .B(n62373), .Y(n38851) );
  NOR2X1 U39343 ( .A(n38853), .B(n38854), .Y(n38852) );
  AND2X1 U39344 ( .A(n63104), .B(n63105), .Y(n38853) );
  AND2X1 U39345 ( .A(n42085), .B(n63108), .Y(n38854) );
  AND2X1 U39346 ( .A(n66098), .B(n66097), .Y(n38855) );
  INVX1 U39347 ( .A(n38855), .Y(n66338) );
  XOR2X1 U39348 ( .A(n39682), .B(n60242), .Y(n38856) );
  NOR2X1 U39349 ( .A(n38858), .B(n66098), .Y(n38857) );
  INVX1 U39350 ( .A(n38857), .Y(n67058) );
  OR2X1 U39351 ( .A(n66345), .B(n66344), .Y(n38858) );
  AND2X1 U39352 ( .A(n59176), .B(n59175), .Y(n38859) );
  NOR2X1 U39353 ( .A(n38862), .B(n38861), .Y(n38860) );
  INVX1 U39354 ( .A(n38860), .Y(n71736) );
  INVX1 U39355 ( .A(n71436), .Y(n38861) );
  AND2X1 U39356 ( .A(n43676), .B(n71433), .Y(n38862) );
  AND2X1 U39357 ( .A(n71469), .B(n71468), .Y(n38863) );
  NOR2X1 U39358 ( .A(n64182), .B(n64057), .Y(n38864) );
  INVX1 U39359 ( .A(n38864), .Y(n64464) );
  OR2X1 U39360 ( .A(n38865), .B(n38866), .Y(n69605) );
  OR2X1 U39361 ( .A(n69266), .B(n69265), .Y(n38865) );
  AND2X1 U39362 ( .A(n69267), .B(n43549), .Y(n38866) );
  XNOR2X1 U39363 ( .A(n64996), .B(n41389), .Y(n38867) );
  INVX1 U39364 ( .A(n38867), .Y(n65106) );
  OR2X1 U39365 ( .A(n43585), .B(n69293), .Y(n69299) );
  OR2X1 U39366 ( .A(n38868), .B(n38869), .Y(n68748) );
  OR2X1 U39367 ( .A(n68747), .B(n68746), .Y(n38868) );
  XOR2X1 U39368 ( .A(n68977), .B(n41118), .Y(n38869) );
  OR2X1 U39369 ( .A(n38870), .B(n38871), .Y(n69548) );
  OR2X1 U39370 ( .A(n68863), .B(n68862), .Y(n38870) );
  AND2X1 U39371 ( .A(n36523), .B(n43683), .Y(n38871) );
  OR2X1 U39372 ( .A(n38872), .B(n68767), .Y(n68461) );
  OR2X1 U39373 ( .A(n43615), .B(n39731), .Y(n38872) );
  NOR2X1 U39374 ( .A(n69972), .B(n69971), .Y(n38873) );
  OR2X1 U39375 ( .A(n43462), .B(n38395), .Y(n59394) );
  AND2X1 U39376 ( .A(n61302), .B(n60877), .Y(n38874) );
  AND2X1 U39377 ( .A(n42016), .B(n60879), .Y(n38875) );
  OR2X1 U39378 ( .A(n38876), .B(n38877), .Y(n66286) );
  OR2X1 U39379 ( .A(n65997), .B(n65996), .Y(n38876) );
  AND2X1 U39380 ( .A(n66004), .B(n66003), .Y(n38877) );
  OR2X1 U39381 ( .A(n38878), .B(n38879), .Y(n65258) );
  AND2X1 U39382 ( .A(n65253), .B(n65252), .Y(n38878) );
  AND2X1 U39383 ( .A(n65257), .B(n41559), .Y(n38879) );
  NAND2X1 U39384 ( .A(n64168), .B(n38619), .Y(n38880) );
  NAND2X1 U39385 ( .A(n64168), .B(n38619), .Y(n38881) );
  OR2X1 U39386 ( .A(n68275), .B(n38882), .Y(n68793) );
  NAND2X1 U39387 ( .A(n38883), .B(n68600), .Y(n38882) );
  OR2X1 U39388 ( .A(n68274), .B(n43588), .Y(n38883) );
  AND2X1 U39389 ( .A(n66309), .B(n66308), .Y(n38884) );
  INVX1 U39390 ( .A(n38884), .Y(n66665) );
  OR2X1 U39391 ( .A(n70789), .B(n41417), .Y(n70821) );
  AND2X1 U39392 ( .A(n41594), .B(n41595), .Y(n38885) );
  AND2X1 U39393 ( .A(n43682), .B(n38886), .Y(n71431) );
  OR2X1 U39394 ( .A(n36762), .B(n71430), .Y(n38886) );
  OR2X1 U39395 ( .A(n40396), .B(n40397), .Y(n38887) );
  AND2X1 U39396 ( .A(n65991), .B(n65992), .Y(n38888) );
  INVX1 U39397 ( .A(n70241), .Y(n38889) );
  AND2X1 U39398 ( .A(n64588), .B(n64589), .Y(n38890) );
  OR2X1 U39399 ( .A(n38891), .B(n38892), .Y(n63988) );
  OR2X1 U39400 ( .A(n41308), .B(n63735), .Y(n38891) );
  AND2X1 U39401 ( .A(n63737), .B(n63991), .Y(n38892) );
  AND2X1 U39402 ( .A(n38893), .B(n68750), .Y(n68454) );
  AND2X1 U39403 ( .A(n40166), .B(n68448), .Y(n38893) );
  NAND2X1 U39404 ( .A(n62997), .B(n38897), .Y(n38894) );
  AND2X1 U39405 ( .A(n38894), .B(n38895), .Y(n62999) );
  OR2X1 U39406 ( .A(n38896), .B(n38902), .Y(n38895) );
  INVX1 U39407 ( .A(n63000), .Y(n38896) );
  AND2X1 U39408 ( .A(n62998), .B(n63000), .Y(n38897) );
  AND2X1 U39409 ( .A(n70228), .B(n70227), .Y(n38898) );
  XOR2X1 U39410 ( .A(n69818), .B(n41638), .Y(n38899) );
  NAND2X1 U39411 ( .A(n62412), .B(n38903), .Y(n38900) );
  AND2X1 U39412 ( .A(n38900), .B(n38901), .Y(n39277) );
  OR2X1 U39413 ( .A(n38902), .B(n62415), .Y(n38901) );
  INVX1 U39414 ( .A(n63320), .Y(n38902) );
  AND2X1 U39415 ( .A(n62413), .B(n63320), .Y(n38903) );
  OR2X1 U39416 ( .A(n38904), .B(n38905), .Y(n72120) );
  AND2X1 U39417 ( .A(n39222), .B(n72119), .Y(n38904) );
  NOR2X1 U39418 ( .A(n38969), .B(n38968), .Y(n38905) );
  NOR2X1 U39419 ( .A(n38907), .B(n38908), .Y(n38906) );
  AND2X1 U39420 ( .A(n62326), .B(n62327), .Y(n38907) );
  AND2X1 U39421 ( .A(n42124), .B(n62328), .Y(n38908) );
  NOR2X1 U39422 ( .A(n38909), .B(n38910), .Y(n40033) );
  OR2X1 U39423 ( .A(n72664), .B(n72663), .Y(n38909) );
  AND2X1 U39424 ( .A(n72714), .B(n72713), .Y(n38910) );
  AND2X1 U39425 ( .A(n62379), .B(n38911), .Y(n38912) );
  INVX1 U39426 ( .A(n62377), .Y(n38911) );
  AND2X1 U39427 ( .A(n67973), .B(n67972), .Y(n38913) );
  NAND2X1 U39428 ( .A(n65112), .B(n65696), .Y(n38914) );
  NOR2X1 U39429 ( .A(n38916), .B(n38917), .Y(n38915) );
  INVX1 U39430 ( .A(n38915), .Y(n60821) );
  AND2X1 U39431 ( .A(n61344), .B(n60817), .Y(n38916) );
  AND2X1 U39432 ( .A(n41816), .B(n60819), .Y(n38917) );
  OR2X1 U39433 ( .A(n38918), .B(n42622), .Y(n48771) );
  INVX1 U39434 ( .A(n39639), .Y(n38919) );
  OR2X1 U39435 ( .A(n61674), .B(n61673), .Y(n61675) );
  INVX1 U39436 ( .A(n39063), .Y(n38920) );
  OR2X1 U39437 ( .A(n38921), .B(n39064), .Y(n61903) );
  NAND2X1 U39438 ( .A(n38920), .B(n61902), .Y(n38921) );
  XNOR2X1 U39439 ( .A(n66077), .B(n38923), .Y(n38922) );
  AND2X1 U39440 ( .A(n66055), .B(n66091), .Y(n38923) );
  NAND2X1 U39441 ( .A(n67586), .B(n67939), .Y(n38924) );
  INVX1 U39442 ( .A(n69501), .Y(n38926) );
  AND2X1 U39443 ( .A(n69626), .B(n38927), .Y(n69625) );
  NOR2X1 U39444 ( .A(n38926), .B(n38962), .Y(n38927) );
  XOR2X1 U39445 ( .A(n67677), .B(n67678), .Y(n38928) );
  INVX1 U39446 ( .A(n38928), .Y(n68046) );
  NAND2X1 U39447 ( .A(n65506), .B(n65172), .Y(n38929) );
  AND2X1 U39448 ( .A(n71104), .B(n43657), .Y(n38930) );
  AND2X1 U39449 ( .A(n71171), .B(n71170), .Y(n38931) );
  INVX1 U39450 ( .A(n41740), .Y(n38932) );
  NOR2X1 U39451 ( .A(n38934), .B(n38935), .Y(n38933) );
  INVX1 U39452 ( .A(n38933), .Y(n71814) );
  AND2X1 U39453 ( .A(n43592), .B(n71605), .Y(n38934) );
  AND2X1 U39454 ( .A(n41664), .B(n71613), .Y(n38935) );
  INVX1 U39455 ( .A(n39075), .Y(n38936) );
  OR2X1 U39456 ( .A(n38937), .B(n39076), .Y(n62129) );
  NAND2X1 U39457 ( .A(n38936), .B(n62128), .Y(n38937) );
  NOR2X1 U39458 ( .A(n38939), .B(n38940), .Y(n38938) );
  INVX1 U39459 ( .A(n38938), .Y(n70592) );
  AND2X1 U39460 ( .A(n43600), .B(n70420), .Y(n38939) );
  AND2X1 U39461 ( .A(n70423), .B(n70422), .Y(n38940) );
  AND2X1 U39462 ( .A(n43653), .B(n71778), .Y(n38941) );
  INVX1 U39463 ( .A(n38941), .Y(n72137) );
  OR2X1 U39464 ( .A(n38942), .B(n38943), .Y(n64314) );
  OR2X1 U39465 ( .A(n38989), .B(n64315), .Y(n38942) );
  NAND2X1 U39466 ( .A(n40200), .B(n64650), .Y(n38943) );
  OR2X1 U39467 ( .A(n42881), .B(n45199), .Y(n38944) );
  AND2X1 U39468 ( .A(n68820), .B(n43657), .Y(n38945) );
  INVX1 U39469 ( .A(n38945), .Y(n68883) );
  NOR2X1 U39470 ( .A(n67958), .B(n39747), .Y(n38946) );
  INVX1 U39471 ( .A(n38946), .Y(n68248) );
  NOR2X1 U39472 ( .A(n40604), .B(n42739), .Y(n38947) );
  OR2X1 U39473 ( .A(n38821), .B(n39770), .Y(n49678) );
  OR2X1 U39474 ( .A(n38948), .B(n38949), .Y(n68165) );
  OR2X1 U39475 ( .A(n67701), .B(n67700), .Y(n38948) );
  AND2X1 U39476 ( .A(n67704), .B(n67703), .Y(n38949) );
  OR2X1 U39477 ( .A(n39048), .B(n39049), .Y(n38950) );
  AND2X1 U39478 ( .A(n68418), .B(n68427), .Y(n38951) );
  OR2X1 U39479 ( .A(n39057), .B(n38952), .Y(n67624) );
  OR2X1 U39480 ( .A(n40741), .B(n40742), .Y(n38952) );
  NOR2X1 U39481 ( .A(n71773), .B(n38953), .Y(n40139) );
  NAND2X1 U39482 ( .A(n71695), .B(n71692), .Y(n38953) );
  NOR2X1 U39483 ( .A(n38956), .B(n38955), .Y(n38954) );
  INVX1 U39484 ( .A(n38954), .Y(n68621) );
  INVX1 U39485 ( .A(n68435), .Y(n38955) );
  OR2X1 U39486 ( .A(n41439), .B(n41384), .Y(n38956) );
  XOR2X1 U39487 ( .A(n66631), .B(n41347), .Y(n66285) );
  NOR2X1 U39488 ( .A(n39864), .B(n39865), .Y(n38957) );
  OR2X1 U39489 ( .A(n38958), .B(n67281), .Y(n38959) );
  INVX1 U39490 ( .A(n67878), .Y(n38958) );
  OR2X1 U39491 ( .A(opcode_opcode_w[20]), .B(n38960), .Y(n40498) );
  OR2X1 U39492 ( .A(n42814), .B(n42763), .Y(n38960) );
  OR2X1 U39493 ( .A(n39893), .B(n39894), .Y(n38961) );
  AND2X1 U39494 ( .A(n41740), .B(n2612), .Y(n48818) );
  XOR2X1 U39495 ( .A(n38963), .B(n69311), .Y(n38962) );
  INVX1 U39496 ( .A(n38962), .Y(n69627) );
  OR2X1 U39497 ( .A(n68952), .B(n68951), .Y(n38963) );
  NOR2X1 U39498 ( .A(n38964), .B(n38965), .Y(n69644) );
  AND2X1 U39499 ( .A(n38222), .B(n43598), .Y(n38964) );
  NAND2X1 U39500 ( .A(n69642), .B(n69641), .Y(n38965) );
  OR2X1 U39501 ( .A(n67679), .B(n38966), .Y(n68037) );
  NAND2X1 U39502 ( .A(n38967), .B(n67681), .Y(n38966) );
  OR2X1 U39503 ( .A(n41377), .B(n38928), .Y(n38967) );
  INVX1 U39504 ( .A(n72123), .Y(n38968) );
  AND2X1 U39505 ( .A(n39689), .B(n39690), .Y(n38970) );
  NAND2X1 U39506 ( .A(n38970), .B(n38971), .Y(n39317) );
  AND2X1 U39507 ( .A(n65499), .B(n65630), .Y(n38971) );
  OR2X1 U39508 ( .A(n65814), .B(n65819), .Y(n66168) );
  OR2X1 U39509 ( .A(n43696), .B(n38973), .Y(n71130) );
  AND2X1 U39510 ( .A(n70189), .B(n70188), .Y(n38973) );
  NAND2X1 U39511 ( .A(n70814), .B(n38591), .Y(n38974) );
  OR2X1 U39512 ( .A(n38974), .B(n38975), .Y(n71141) );
  OR2X1 U39513 ( .A(n43697), .B(n40566), .Y(n38975) );
  NOR2X1 U39514 ( .A(n38977), .B(n38978), .Y(n38976) );
  OR2X1 U39515 ( .A(n63289), .B(n63288), .Y(n38977) );
  AND2X1 U39516 ( .A(n63292), .B(n63291), .Y(n38978) );
  OR2X1 U39517 ( .A(n38979), .B(n38980), .Y(n65445) );
  INVX1 U39518 ( .A(n65710), .Y(n38979) );
  AND2X1 U39519 ( .A(n39016), .B(n65699), .Y(n38980) );
  XOR2X1 U39520 ( .A(n62870), .B(n62507), .Y(n38981) );
  INVX1 U39521 ( .A(n40518), .Y(n38982) );
  XNOR2X1 U39522 ( .A(n70790), .B(n38983), .Y(n71137) );
  XOR2X1 U39523 ( .A(n70492), .B(n41281), .Y(n38983) );
  OR2X1 U39524 ( .A(n38984), .B(n38985), .Y(n68738) );
  OR2X1 U39525 ( .A(n67800), .B(n67799), .Y(n38984) );
  AND2X1 U39526 ( .A(n67802), .B(n67801), .Y(n38985) );
  AND2X1 U39527 ( .A(n68719), .B(n68720), .Y(n38986) );
  OR2X1 U39528 ( .A(n43656), .B(n71104), .Y(n71106) );
  OR2X1 U39529 ( .A(n38987), .B(n38988), .Y(n70444) );
  AND2X1 U39530 ( .A(n43619), .B(n69939), .Y(n38987) );
  AND2X1 U39531 ( .A(n69942), .B(n70147), .Y(n38988) );
  AND2X1 U39532 ( .A(n64642), .B(n64005), .Y(n38989) );
  OR2X1 U39533 ( .A(n59749), .B(n38991), .Y(n38992) );
  INVX1 U39534 ( .A(n59526), .Y(n38990) );
  INVX1 U39535 ( .A(n59525), .Y(n38991) );
  AND2X1 U39536 ( .A(n61534), .B(n61533), .Y(n38993) );
  AND2X1 U39537 ( .A(n40278), .B(n59136), .Y(n38994) );
  AND2X1 U39538 ( .A(n38995), .B(n38996), .Y(n39372) );
  NOR2X1 U39539 ( .A(n69844), .B(n69845), .Y(n38995) );
  AND2X1 U39540 ( .A(n39981), .B(n39982), .Y(n38996) );
  NAND2X1 U39541 ( .A(n66455), .B(n38999), .Y(n38997) );
  AND2X1 U39542 ( .A(n38997), .B(n38998), .Y(n67020) );
  OR2X1 U39543 ( .A(n66798), .B(n66460), .Y(n38998) );
  AND2X1 U39544 ( .A(n66454), .B(n66800), .Y(n38999) );
  OR2X1 U39545 ( .A(n62523), .B(n39000), .Y(n62859) );
  NAND2X1 U39546 ( .A(n39001), .B(n62524), .Y(n39000) );
  OR2X1 U39547 ( .A(n62849), .B(n62522), .Y(n39001) );
  OR2X1 U39548 ( .A(n39002), .B(n39003), .Y(n68495) );
  AND2X1 U39549 ( .A(n43561), .B(n67646), .Y(n39002) );
  AND2X1 U39550 ( .A(n40953), .B(n67648), .Y(n39003) );
  AND2X1 U39551 ( .A(n68914), .B(n68920), .Y(n39004) );
  AND2X1 U39552 ( .A(n69562), .B(n43691), .Y(n39005) );
  INVX1 U39553 ( .A(n39005), .Y(n70186) );
  INVX1 U39554 ( .A(n39593), .Y(n39006) );
  NOR2X1 U39555 ( .A(n39007), .B(n39594), .Y(n41587) );
  NAND2X1 U39556 ( .A(n39006), .B(n59592), .Y(n39007) );
  OR2X1 U39557 ( .A(n40458), .B(n40459), .Y(n39008) );
  OR2X1 U39558 ( .A(n39009), .B(n39010), .Y(n46058) );
  OR2X1 U39559 ( .A(n46052), .B(n46051), .Y(n39009) );
  OR2X1 U39560 ( .A(n46057), .B(n46056), .Y(n39010) );
  NAND2X1 U39561 ( .A(n71152), .B(n71153), .Y(n39011) );
  AND2X1 U39562 ( .A(n69551), .B(n43682), .Y(n39012) );
  INVX1 U39563 ( .A(n39012), .Y(n70172) );
  INVX1 U39564 ( .A(n39891), .Y(n39013) );
  XNOR2X1 U39565 ( .A(n64970), .B(n64695), .Y(n39014) );
  OR2X1 U39566 ( .A(n43514), .B(n70787), .Y(n70822) );
  OR2X1 U39567 ( .A(n62381), .B(n62380), .Y(n62390) );
  OR2X1 U39568 ( .A(n63772), .B(n39015), .Y(n63314) );
  INVX1 U39569 ( .A(n63502), .Y(n39015) );
  NAND2X1 U39570 ( .A(n65112), .B(n65696), .Y(n39016) );
  OR2X1 U39571 ( .A(n61585), .B(n61584), .Y(n61586) );
  OR2X1 U39572 ( .A(n40065), .B(n40066), .Y(n39017) );
  XOR2X1 U39573 ( .A(n39019), .B(n39020), .Y(n39018) );
  INVX1 U39574 ( .A(n39018), .Y(n66535) );
  INVX1 U39575 ( .A(n65969), .Y(n39019) );
  XOR2X1 U39576 ( .A(n65970), .B(n43666), .Y(n39020) );
  OR2X1 U39577 ( .A(n63438), .B(n39021), .Y(n63726) );
  NOR2X1 U39578 ( .A(n63675), .B(n63674), .Y(n39021) );
  AND2X1 U39579 ( .A(n40392), .B(n42709), .Y(n39022) );
  INVX1 U39580 ( .A(n39022), .Y(n59157) );
  AND2X1 U39581 ( .A(n39023), .B(n39024), .Y(n69855) );
  OR2X1 U39582 ( .A(n39985), .B(n39958), .Y(n39023) );
  OR2X1 U39583 ( .A(n41426), .B(n43574), .Y(n39024) );
  OR2X1 U39584 ( .A(n68562), .B(n39391), .Y(n68258) );
  OR2X1 U39585 ( .A(n65506), .B(n65172), .Y(n65171) );
  AND2X1 U39586 ( .A(n68700), .B(n68702), .Y(n39025) );
  INVX1 U39587 ( .A(n38697), .Y(n39026) );
  OR2X1 U39588 ( .A(n39027), .B(n39028), .Y(n64953) );
  INVX1 U39589 ( .A(n64689), .Y(n39027) );
  NAND2X1 U39590 ( .A(n39026), .B(n64688), .Y(n39028) );
  AND2X1 U39591 ( .A(n65858), .B(n66015), .Y(n39029) );
  INVX1 U39592 ( .A(n39029), .Y(n66020) );
  NAND2X1 U39593 ( .A(n43619), .B(n69611), .Y(n39030) );
  OR2X1 U39594 ( .A(n39031), .B(n39032), .Y(n63474) );
  OR2X1 U39595 ( .A(n63138), .B(n63137), .Y(n39031) );
  AND2X1 U39596 ( .A(n63139), .B(n63467), .Y(n39032) );
  OR2X1 U39597 ( .A(n39033), .B(n37363), .Y(n67855) );
  OR2X1 U39598 ( .A(n67552), .B(n67551), .Y(n39033) );
  NAND2X1 U39599 ( .A(n70137), .B(n39037), .Y(n39034) );
  NAND2X1 U39600 ( .A(n39034), .B(n39035), .Y(n41104) );
  OR2X1 U39601 ( .A(n39036), .B(n70140), .Y(n39035) );
  INVX1 U39602 ( .A(n70141), .Y(n39036) );
  AND2X1 U39603 ( .A(n70138), .B(n70141), .Y(n39037) );
  OR2X1 U39604 ( .A(n39307), .B(n39040), .Y(n39038) );
  AND2X1 U39605 ( .A(n39038), .B(n39039), .Y(n70127) );
  OR2X1 U39606 ( .A(n39927), .B(n70126), .Y(n39039) );
  OR2X1 U39607 ( .A(n39927), .B(n39927), .Y(n39040) );
  XOR2X1 U39608 ( .A(n41299), .B(n39041), .Y(n71735) );
  XOR2X1 U39609 ( .A(n71429), .B(n71699), .Y(n39041) );
  NOR2X1 U39610 ( .A(n39388), .B(n39389), .Y(n39042) );
  OR2X1 U39611 ( .A(n39285), .B(n39286), .Y(n39043) );
  NOR2X1 U39612 ( .A(n39045), .B(n39046), .Y(n39044) );
  INVX1 U39613 ( .A(n39044), .Y(n59309) );
  INVX1 U39614 ( .A(n59368), .Y(n39045) );
  AND2X1 U39615 ( .A(n59335), .B(n59371), .Y(n39046) );
  NOR2X1 U39616 ( .A(n39048), .B(n39049), .Y(n39047) );
  OR2X1 U39617 ( .A(n69683), .B(n69682), .Y(n39048) );
  AND2X1 U39618 ( .A(n69685), .B(n69684), .Y(n39049) );
  OR2X1 U39619 ( .A(n43632), .B(n71185), .Y(n39050) );
  OR2X1 U39620 ( .A(n69611), .B(n39295), .Y(n70147) );
  NOR2X1 U39621 ( .A(n39052), .B(n39053), .Y(n39051) );
  INVX1 U39622 ( .A(n39051), .Y(n59180) );
  AND2X1 U39623 ( .A(n59196), .B(n38859), .Y(n39052) );
  AND2X1 U39624 ( .A(n59179), .B(n59178), .Y(n39053) );
  OR2X1 U39625 ( .A(n39054), .B(n39055), .Y(n69040) );
  INVX1 U39626 ( .A(n41521), .Y(n39054) );
  AND2X1 U39627 ( .A(n68411), .B(n68410), .Y(n39055) );
  OR2X1 U39628 ( .A(n59764), .B(n39056), .Y(n59768) );
  AND2X1 U39629 ( .A(n59765), .B(n41328), .Y(n39056) );
  AND2X1 U39630 ( .A(n67632), .B(n41045), .Y(n39057) );
  AND2X1 U39631 ( .A(n41319), .B(n39058), .Y(n66948) );
  NOR2X1 U39632 ( .A(n43587), .B(n67546), .Y(n39058) );
  OR2X1 U39633 ( .A(n39059), .B(n39060), .Y(n68996) );
  INVX1 U39634 ( .A(n68999), .Y(n39059) );
  AND2X1 U39635 ( .A(n42026), .B(n68997), .Y(n39060) );
  OR2X1 U39636 ( .A(n36719), .B(n43770), .Y(n60111) );
  OR2X1 U39637 ( .A(n60974), .B(n39193), .Y(n39061) );
  OR2X1 U39638 ( .A(n37395), .B(n60007), .Y(n60008) );
  NOR2X1 U39639 ( .A(n39063), .B(n39064), .Y(n39062) );
  INVX1 U39640 ( .A(n39062), .Y(n61901) );
  AND2X1 U39641 ( .A(n61898), .B(n61899), .Y(n39063) );
  AND2X1 U39642 ( .A(n42002), .B(n61900), .Y(n39064) );
  NOR2X1 U39643 ( .A(n40566), .B(n39065), .Y(n41019) );
  NAND2X1 U39644 ( .A(n38591), .B(n70814), .Y(n39065) );
  AND2X1 U39645 ( .A(n70715), .B(n70714), .Y(n39066) );
  OR2X1 U39646 ( .A(n39794), .B(n42825), .Y(n59128) );
  NAND2X1 U39647 ( .A(n37914), .B(n65584), .Y(n39067) );
  OR2X1 U39648 ( .A(n61666), .B(n61665), .Y(n61667) );
  OR2X1 U39649 ( .A(n39068), .B(n39069), .Y(n63732) );
  INVX1 U39650 ( .A(n42032), .Y(n39068) );
  NOR2X1 U39651 ( .A(n63666), .B(n39223), .Y(n39069) );
  OR2X1 U39652 ( .A(n39070), .B(n39071), .Y(n62566) );
  INVX1 U39653 ( .A(n42095), .Y(n39070) );
  AND2X1 U39654 ( .A(n38250), .B(n62565), .Y(n39071) );
  OR2X1 U39655 ( .A(n39072), .B(n39073), .Y(n70940) );
  OR2X1 U39656 ( .A(n70695), .B(n70694), .Y(n39072) );
  AND2X1 U39657 ( .A(n70697), .B(n70704), .Y(n39073) );
  NOR2X1 U39658 ( .A(n39075), .B(n39076), .Y(n39074) );
  INVX1 U39659 ( .A(n39074), .Y(n62127) );
  AND2X1 U39660 ( .A(n62124), .B(n62125), .Y(n39075) );
  AND2X1 U39661 ( .A(n42110), .B(n62126), .Y(n39076) );
  OR2X1 U39662 ( .A(n39077), .B(n39078), .Y(n65581) );
  AND2X1 U39663 ( .A(n65567), .B(n43713), .Y(n39077) );
  AND2X1 U39664 ( .A(n65572), .B(n65571), .Y(n39078) );
  OR2X1 U39665 ( .A(n37402), .B(n40088), .Y(n70851) );
  OR2X1 U39666 ( .A(n39079), .B(n39080), .Y(n70771) );
  OR2X1 U39667 ( .A(n70457), .B(n70456), .Y(n39079) );
  AND2X1 U39668 ( .A(n70460), .B(n43669), .Y(n39080) );
  AND2X1 U39669 ( .A(n65245), .B(n43638), .Y(n39081) );
  NOR2X1 U39670 ( .A(n42226), .B(n39083), .Y(n39082) );
  INVX1 U39671 ( .A(n39082), .Y(n64066) );
  INVX1 U39672 ( .A(n43609), .Y(n39083) );
  AND2X1 U39673 ( .A(n39363), .B(n39092), .Y(n39084) );
  INVX1 U39674 ( .A(n42086), .Y(n39085) );
  OR2X1 U39675 ( .A(n39119), .B(n39087), .Y(n67712) );
  AND2X1 U39676 ( .A(n67718), .B(n67461), .Y(n39087) );
  AND2X1 U39677 ( .A(n61440), .B(n61439), .Y(n39088) );
  AND2X1 U39678 ( .A(n42053), .B(n61437), .Y(n39089) );
  OR2X1 U39679 ( .A(n39876), .B(n39877), .Y(n39090) );
  NOR2X1 U39680 ( .A(n43514), .B(n68842), .Y(n39091) );
  NAND2X1 U39681 ( .A(n39363), .B(n39092), .Y(n68507) );
  NOR2X1 U39682 ( .A(n39093), .B(n38552), .Y(n39092) );
  AND2X1 U39683 ( .A(n40303), .B(n68572), .Y(n39093) );
  OR2X1 U39684 ( .A(n39094), .B(n39095), .Y(n64593) );
  OR2X1 U39685 ( .A(n64590), .B(n64589), .Y(n39094) );
  AND2X1 U39686 ( .A(n38285), .B(n64591), .Y(n39095) );
  NAND2X1 U39687 ( .A(n39725), .B(n39096), .Y(n71763) );
  AND2X1 U39688 ( .A(n71688), .B(n43643), .Y(n39096) );
  OR2X1 U39689 ( .A(n39097), .B(n37357), .Y(n72658) );
  AND2X1 U39690 ( .A(n72656), .B(n72655), .Y(n39097) );
  NOR2X1 U39691 ( .A(n39099), .B(n39100), .Y(n39098) );
  AND2X1 U39692 ( .A(n61329), .B(n39450), .Y(n39099) );
  AND2X1 U39693 ( .A(n41890), .B(n60839), .Y(n39100) );
  OR2X1 U39694 ( .A(n59859), .B(n59860), .Y(n59861) );
  NOR2X1 U39695 ( .A(n64825), .B(n64826), .Y(n39101) );
  INVX1 U39696 ( .A(n39101), .Y(n64828) );
  AND2X1 U39697 ( .A(n65427), .B(n65426), .Y(n39102) );
  OR2X1 U39698 ( .A(n39091), .B(n69220), .Y(n39595) );
  OR2X1 U39699 ( .A(n43508), .B(n69578), .Y(n39103) );
  OR2X1 U39700 ( .A(n43507), .B(n69581), .Y(n39104) );
  OR2X1 U39701 ( .A(n60649), .B(n60648), .Y(n60652) );
  OR2X1 U39702 ( .A(n39105), .B(n36768), .Y(n64472) );
  AND2X1 U39703 ( .A(n64699), .B(n64700), .Y(n39105) );
  OR2X1 U39704 ( .A(n71194), .B(n39106), .Y(n71439) );
  NAND2X1 U39705 ( .A(n39050), .B(n71197), .Y(n39106) );
  OR2X1 U39706 ( .A(n72060), .B(n43577), .Y(n72062) );
  OR2X1 U39707 ( .A(n39107), .B(n37384), .Y(n69267) );
  AND2X1 U39708 ( .A(n41034), .B(n38842), .Y(n39107) );
  AND2X1 U39709 ( .A(n65697), .B(n39108), .Y(n65701) );
  NOR2X1 U39710 ( .A(n38600), .B(n65698), .Y(n39108) );
  AND2X1 U39711 ( .A(n65019), .B(n40272), .Y(n39109) );
  XNOR2X1 U39712 ( .A(n71150), .B(n71151), .Y(n71433) );
  NOR2X1 U39713 ( .A(n62375), .B(n62376), .Y(n39110) );
  NOR2X1 U39714 ( .A(n39110), .B(n39111), .Y(n40452) );
  OR2X1 U39715 ( .A(n39112), .B(n62377), .Y(n39111) );
  INVX1 U39716 ( .A(n62379), .Y(n39112) );
  NOR2X1 U39717 ( .A(n65446), .B(n65445), .Y(n39113) );
  OR2X1 U39718 ( .A(n39755), .B(n39756), .Y(n39114) );
  INVX1 U39719 ( .A(n42740), .Y(n39115) );
  INVX1 U39720 ( .A(n39115), .Y(n39116) );
  NOR2X1 U39721 ( .A(n39118), .B(n37401), .Y(n39117) );
  INVX1 U39722 ( .A(n39117), .Y(n65687) );
  AND2X1 U39723 ( .A(n65357), .B(n66043), .Y(n39118) );
  AND2X1 U39724 ( .A(n67457), .B(n67714), .Y(n39119) );
  AND2X1 U39725 ( .A(n61124), .B(n39122), .Y(n39120) );
  OR2X1 U39726 ( .A(n39120), .B(n39121), .Y(n62395) );
  AND2X1 U39727 ( .A(n40185), .B(n40045), .Y(n39121) );
  AND2X1 U39728 ( .A(n61125), .B(n40185), .Y(n39122) );
  OR2X1 U39729 ( .A(n39123), .B(n37389), .Y(n70696) );
  AND2X1 U39730 ( .A(n70693), .B(n70692), .Y(n39123) );
  OR2X1 U39731 ( .A(n39124), .B(n39125), .Y(n71080) );
  AND2X1 U39732 ( .A(n70912), .B(n42993), .Y(n39124) );
  AND2X1 U39733 ( .A(n70581), .B(n70580), .Y(n39125) );
  AND2X1 U39734 ( .A(n39704), .B(n39556), .Y(n39126) );
  AND2X1 U39735 ( .A(n65290), .B(n39127), .Y(n65288) );
  INVX1 U39736 ( .A(n41037), .Y(n39127) );
  OR2X1 U39737 ( .A(n37387), .B(n39567), .Y(n39128) );
  NAND2X1 U39738 ( .A(n40313), .B(n65763), .Y(n39129) );
  INVX1 U39739 ( .A(n42154), .Y(n39130) );
  INVX1 U39740 ( .A(n42154), .Y(n39131) );
  INVX1 U39741 ( .A(n39130), .Y(n39132) );
  INVX1 U39742 ( .A(n39130), .Y(n39133) );
  INVX1 U39743 ( .A(n39130), .Y(n39134) );
  INVX1 U39744 ( .A(n39130), .Y(n39135) );
  INVX1 U39745 ( .A(n39131), .Y(n39136) );
  INVX1 U39746 ( .A(n39131), .Y(n39137) );
  INVX1 U39747 ( .A(n39131), .Y(n39138) );
  INVX1 U39748 ( .A(n39131), .Y(n39139) );
  NOR2X1 U39749 ( .A(n39141), .B(n39142), .Y(n39140) );
  AND2X1 U39750 ( .A(n60413), .B(n60412), .Y(n39141) );
  AND2X1 U39751 ( .A(n60415), .B(n60414), .Y(n39142) );
  AND2X1 U39752 ( .A(n43705), .B(n64573), .Y(n39143) );
  AND2X1 U39753 ( .A(n64576), .B(n64575), .Y(n39144) );
  AND2X1 U39754 ( .A(n69933), .B(n43636), .Y(n39145) );
  XNOR2X1 U39755 ( .A(n40764), .B(n64990), .Y(n39146) );
  NAND2X1 U39756 ( .A(n40172), .B(n65273), .Y(n39147) );
  OR2X1 U39757 ( .A(n68940), .B(n39148), .Y(n69626) );
  AND2X1 U39758 ( .A(n43592), .B(n69499), .Y(n39148) );
  OR2X1 U39759 ( .A(n60534), .B(n36784), .Y(n60535) );
  NOR2X1 U39760 ( .A(n39150), .B(n39151), .Y(n39149) );
  INVX1 U39761 ( .A(n39149), .Y(n60836) );
  AND2X1 U39762 ( .A(n61333), .B(n60833), .Y(n39150) );
  AND2X1 U39763 ( .A(n41870), .B(n60834), .Y(n39151) );
  OR2X1 U39764 ( .A(n38293), .B(n39152), .Y(n65067) );
  AND2X1 U39765 ( .A(n64112), .B(n63815), .Y(n39152) );
  AND2X1 U39766 ( .A(n70137), .B(n70138), .Y(n39153) );
  INVX1 U39767 ( .A(n39153), .Y(n69936) );
  AND2X1 U39768 ( .A(n66548), .B(n43691), .Y(n39154) );
  OR2X1 U39769 ( .A(n60755), .B(n39155), .Y(n60554) );
  AND2X1 U39770 ( .A(n60756), .B(n60754), .Y(n39155) );
  OR2X1 U39771 ( .A(n39156), .B(n68020), .Y(n68277) );
  OR2X1 U39772 ( .A(n68019), .B(n68018), .Y(n39156) );
  OR2X1 U39773 ( .A(n70187), .B(n69231), .Y(n39157) );
  OR2X1 U39774 ( .A(n39158), .B(n39568), .Y(n63461) );
  OR2X1 U39775 ( .A(n41599), .B(n41639), .Y(n39158) );
  XNOR2X1 U39776 ( .A(n68753), .B(n40980), .Y(n39159) );
  AND2X1 U39777 ( .A(n67973), .B(n67972), .Y(n39160) );
  INVX1 U39778 ( .A(n38913), .Y(n67952) );
  OR2X1 U39779 ( .A(n43627), .B(n66214), .Y(n66608) );
  AND2X1 U39780 ( .A(n65144), .B(n39161), .Y(n66181) );
  INVX1 U39781 ( .A(n66179), .Y(n39161) );
  AND2X1 U39782 ( .A(n63437), .B(n63436), .Y(n39162) );
  INVX1 U39783 ( .A(n43783), .Y(n39163) );
  INVX1 U39784 ( .A(n43785), .Y(n39164) );
  NOR2X1 U39785 ( .A(n65718), .B(n39165), .Y(n40246) );
  NAND2X1 U39786 ( .A(n39166), .B(n66088), .Y(n39165) );
  AND2X1 U39787 ( .A(n65717), .B(n65716), .Y(n39166) );
  OR2X1 U39788 ( .A(n39167), .B(n39168), .Y(n39476) );
  OR2X1 U39789 ( .A(n38283), .B(n69530), .Y(n39167) );
  OR2X1 U39790 ( .A(n69867), .B(n43672), .Y(n39168) );
  OR2X1 U39791 ( .A(n39169), .B(n39170), .Y(n59336) );
  AND2X1 U39792 ( .A(n59289), .B(n59290), .Y(n39169) );
  AND2X1 U39793 ( .A(n59292), .B(n59291), .Y(n39170) );
  XNOR2X1 U39794 ( .A(n66478), .B(n66010), .Y(n39171) );
  OR2X1 U39795 ( .A(n63099), .B(n63100), .Y(n63103) );
  NOR2X1 U39796 ( .A(n39173), .B(n39174), .Y(n39172) );
  INVX1 U39797 ( .A(n39172), .Y(n60793) );
  AND2X1 U39798 ( .A(n60796), .B(n60477), .Y(n39173) );
  AND2X1 U39799 ( .A(n41814), .B(n60479), .Y(n39174) );
  INVX1 U39800 ( .A(n39290), .Y(n39175) );
  OR2X1 U39801 ( .A(n39176), .B(n39291), .Y(n61918) );
  NAND2X1 U39802 ( .A(n39175), .B(n61917), .Y(n39176) );
  XOR2X1 U39803 ( .A(n71733), .B(n39412), .Y(n39177) );
  OR2X1 U39804 ( .A(n39178), .B(n39179), .Y(n45522) );
  OR2X1 U39805 ( .A(n46526), .B(n38473), .Y(n39178) );
  OR2X1 U39806 ( .A(n46577), .B(n37094), .Y(n39179) );
  INVX1 U39807 ( .A(n39303), .Y(n39180) );
  OR2X1 U39808 ( .A(n39181), .B(n39304), .Y(n62814) );
  NAND2X1 U39809 ( .A(n39180), .B(n62813), .Y(n39181) );
  OR2X1 U39810 ( .A(n39182), .B(n43771), .Y(n59994) );
  INVX1 U39811 ( .A(n42717), .Y(n39182) );
  OR2X1 U39812 ( .A(n39401), .B(n39402), .Y(n39183) );
  OR2X1 U39813 ( .A(n39464), .B(n39465), .Y(n39184) );
  OR2X1 U39814 ( .A(n39467), .B(n39468), .Y(n39185) );
  AND2X1 U39815 ( .A(n39186), .B(n69524), .Y(n69521) );
  INVX1 U39816 ( .A(n43632), .Y(n39186) );
  XOR2X1 U39817 ( .A(n68927), .B(n40745), .Y(n39187) );
  AND2X1 U39818 ( .A(n39189), .B(n39188), .Y(n47341) );
  INVX1 U39819 ( .A(n42888), .Y(n39188) );
  OR2X1 U39820 ( .A(n47339), .B(n47338), .Y(n39189) );
  OR2X1 U39821 ( .A(n39190), .B(n39191), .Y(n45780) );
  OR2X1 U39822 ( .A(n46577), .B(n37043), .Y(n39190) );
  OR2X1 U39823 ( .A(n46024), .B(n45612), .Y(n39191) );
  AND2X1 U39824 ( .A(n38493), .B(n38827), .Y(n39192) );
  OR2X1 U39825 ( .A(n42700), .B(n39770), .Y(n49677) );
  NOR2X1 U39826 ( .A(n39615), .B(n39616), .Y(n39193) );
  NOR2X1 U39827 ( .A(n39956), .B(n39957), .Y(n39194) );
  INVX1 U39828 ( .A(n42490), .Y(n39195) );
  INVX1 U39829 ( .A(n42490), .Y(n39196) );
  INVX1 U39830 ( .A(n36601), .Y(n39197) );
  INVX1 U39831 ( .A(n36601), .Y(n39198) );
  NAND2X1 U39832 ( .A(n61143), .B(n39202), .Y(n39199) );
  AND2X1 U39833 ( .A(n39199), .B(n39200), .Y(n62972) );
  OR2X1 U39834 ( .A(n39201), .B(n61146), .Y(n39200) );
  INVX1 U39835 ( .A(n62482), .Y(n39201) );
  AND2X1 U39836 ( .A(n61144), .B(n62482), .Y(n39202) );
  OR2X1 U39837 ( .A(n39203), .B(n39204), .Y(n59252) );
  AND2X1 U39838 ( .A(n59165), .B(n59131), .Y(n39203) );
  AND2X1 U39839 ( .A(n39022), .B(n59133), .Y(n39204) );
  AND2X1 U39840 ( .A(n60204), .B(n60203), .Y(n39205) );
  NAND2X1 U39841 ( .A(n39680), .B(n40390), .Y(n39206) );
  AND2X1 U39842 ( .A(n63807), .B(n63808), .Y(n39207) );
  OR2X1 U39843 ( .A(n36719), .B(n40444), .Y(n59199) );
  OR2X1 U39844 ( .A(n39209), .B(n39208), .Y(n62886) );
  INVX1 U39845 ( .A(n62883), .Y(n39208) );
  OR2X1 U39846 ( .A(n41061), .B(n41085), .Y(n39209) );
  AND2X1 U39847 ( .A(n45313), .B(n45312), .Y(n39210) );
  INVX1 U39848 ( .A(n39210), .Y(n48104) );
  NOR2X1 U39849 ( .A(n45521), .B(n39214), .Y(n39211) );
  OR2X1 U39850 ( .A(n39211), .B(n39212), .Y(n45626) );
  AND2X1 U39851 ( .A(n39213), .B(n45613), .Y(n39212) );
  INVX1 U39852 ( .A(n45922), .Y(n39213) );
  OR2X1 U39853 ( .A(n45611), .B(n45922), .Y(n39214) );
  NOR2X1 U39854 ( .A(n39216), .B(n39217), .Y(n39215) );
  INVX1 U39855 ( .A(n39215), .Y(n61241) );
  OR2X1 U39856 ( .A(n61065), .B(n61064), .Y(n39216) );
  AND2X1 U39857 ( .A(n61067), .B(n61066), .Y(n39217) );
  XNOR2X1 U39858 ( .A(n39218), .B(n41134), .Y(n39985) );
  INVX1 U39859 ( .A(n69294), .Y(n39218) );
  NOR2X1 U39860 ( .A(n39220), .B(n39221), .Y(n39219) );
  INVX1 U39861 ( .A(n39219), .Y(n61042) );
  AND2X1 U39862 ( .A(n60582), .B(n38687), .Y(n39220) );
  AND2X1 U39863 ( .A(n41678), .B(n60583), .Y(n39221) );
  AND2X1 U39864 ( .A(n40192), .B(n40456), .Y(n39222) );
  OR2X1 U39865 ( .A(n39224), .B(n39225), .Y(n61106) );
  OR2X1 U39866 ( .A(n41337), .B(n61108), .Y(n39224) );
  AND2X1 U39867 ( .A(n60895), .B(n60894), .Y(n39225) );
  XOR2X1 U39868 ( .A(n41124), .B(n69218), .Y(n39226) );
  OR2X1 U39869 ( .A(n61699), .B(n61698), .Y(n61700) );
  AND2X1 U39870 ( .A(n39177), .B(n39227), .Y(n71740) );
  NOR2X1 U39871 ( .A(n43682), .B(n43511), .Y(n39227) );
  OR2X1 U39872 ( .A(n39228), .B(n39229), .Y(n60159) );
  INVX1 U39873 ( .A(n41894), .Y(n39228) );
  AND2X1 U39874 ( .A(n36493), .B(n60158), .Y(n39229) );
  NOR2X1 U39875 ( .A(n39231), .B(n39232), .Y(n39230) );
  AND2X1 U39876 ( .A(n38502), .B(n59979), .Y(n39231) );
  AND2X1 U39877 ( .A(n59836), .B(n59835), .Y(n39232) );
  OR2X1 U39878 ( .A(n39233), .B(n39234), .Y(n45709) );
  OR2X1 U39879 ( .A(n45612), .B(n45922), .Y(n39233) );
  OR2X1 U39880 ( .A(n46206), .B(n37057), .Y(n39234) );
  AND2X1 U39881 ( .A(n39235), .B(n70704), .Y(n70694) );
  INVX1 U39882 ( .A(n72200), .Y(n39235) );
  OR2X1 U39883 ( .A(n39789), .B(n39790), .Y(n39236) );
  NAND2X1 U39884 ( .A(n69039), .B(n69040), .Y(n39237) );
  XNOR2X1 U39885 ( .A(n41574), .B(n60934), .Y(n39238) );
  OR2X1 U39886 ( .A(n39239), .B(n39240), .Y(n71142) );
  OR2X1 U39887 ( .A(n39922), .B(n71140), .Y(n39239) );
  NAND2X1 U39888 ( .A(n39268), .B(n39269), .Y(n39240) );
  NAND2X1 U39889 ( .A(n70167), .B(n43528), .Y(n39241) );
  OR2X1 U39890 ( .A(n39242), .B(n39243), .Y(n71742) );
  OR2X1 U39891 ( .A(n43507), .B(n40304), .Y(n39242) );
  AND2X1 U39892 ( .A(n39576), .B(n71741), .Y(n39243) );
  OR2X1 U39893 ( .A(n39244), .B(n39245), .Y(n60155) );
  INVX1 U39894 ( .A(n60325), .Y(n39244) );
  AND2X1 U39895 ( .A(n36490), .B(n60326), .Y(n39245) );
  OR2X1 U39896 ( .A(n41038), .B(n39249), .Y(n39246) );
  AND2X1 U39897 ( .A(n39246), .B(n39247), .Y(n62998) );
  OR2X1 U39898 ( .A(n39248), .B(n62411), .Y(n39247) );
  INVX1 U39899 ( .A(n41506), .Y(n39248) );
  OR2X1 U39900 ( .A(n61128), .B(n39248), .Y(n39249) );
  OR2X1 U39901 ( .A(n39250), .B(n39251), .Y(n61424) );
  INVX1 U39902 ( .A(n42010), .Y(n39250) );
  AND2X1 U39903 ( .A(n37947), .B(n38279), .Y(n39251) );
  NOR2X1 U39904 ( .A(n39253), .B(n39254), .Y(n39252) );
  INVX1 U39905 ( .A(n39252), .Y(n72689) );
  AND2X1 U39906 ( .A(n72676), .B(n43684), .Y(n39253) );
  AND2X1 U39907 ( .A(n72683), .B(n72682), .Y(n39254) );
  XNOR2X1 U39908 ( .A(n71436), .B(n71149), .Y(n39255) );
  OR2X1 U39909 ( .A(n39107), .B(n37384), .Y(n69513) );
  NAND2X1 U39910 ( .A(n65946), .B(n39258), .Y(n39256) );
  NAND2X1 U39911 ( .A(n39257), .B(n39256), .Y(n41219) );
  OR2X1 U39912 ( .A(n39154), .B(n65948), .Y(n39257) );
  AND2X1 U39913 ( .A(n66547), .B(n37932), .Y(n39258) );
  AND2X1 U39914 ( .A(n64639), .B(n64638), .Y(n39259) );
  AND2X1 U39915 ( .A(n69443), .B(n69442), .Y(n39260) );
  INVX1 U39916 ( .A(n40112), .Y(n39261) );
  NOR2X1 U39917 ( .A(n39262), .B(n40113), .Y(n41286) );
  NAND2X1 U39918 ( .A(n39261), .B(n38267), .Y(n39262) );
  OR2X1 U39919 ( .A(n39263), .B(n39264), .Y(n68857) );
  OR2X1 U39920 ( .A(n68827), .B(n68828), .Y(n39263) );
  AND2X1 U39921 ( .A(n39841), .B(n68877), .Y(n39264) );
  OR2X1 U39922 ( .A(n40252), .B(n39265), .Y(n70472) );
  OR2X1 U39923 ( .A(n40312), .B(n43656), .Y(n39265) );
  AND2X1 U39924 ( .A(n65180), .B(n43635), .Y(n39266) );
  AND2X1 U39925 ( .A(n63521), .B(n39267), .Y(n63523) );
  INVX1 U39926 ( .A(n63524), .Y(n39267) );
  NAND2X1 U39927 ( .A(n70792), .B(n39270), .Y(n39268) );
  AND2X1 U39928 ( .A(n70791), .B(n43696), .Y(n39270) );
  OR2X1 U39929 ( .A(n40112), .B(n40113), .Y(n39271) );
  OR2X1 U39930 ( .A(n39272), .B(n39273), .Y(n65098) );
  OR2X1 U39931 ( .A(n64719), .B(n64718), .Y(n39272) );
  AND2X1 U39932 ( .A(n65106), .B(n64720), .Y(n39273) );
  AND2X1 U39933 ( .A(n69673), .B(n43000), .Y(n39274) );
  INVX1 U39934 ( .A(n39274), .Y(n69966) );
  AND2X1 U39935 ( .A(n61127), .B(n61126), .Y(n39275) );
  INVX1 U39936 ( .A(n39275), .Y(n62411) );
  OR2X1 U39937 ( .A(n39277), .B(n39276), .Y(n39423) );
  INVX1 U39938 ( .A(n62998), .Y(n39276) );
  OR2X1 U39939 ( .A(n39278), .B(n39279), .Y(n66463) );
  AND2X1 U39940 ( .A(n66166), .B(n66163), .Y(n39278) );
  AND2X1 U39941 ( .A(n66172), .B(n66171), .Y(n39279) );
  OR2X1 U39942 ( .A(n39280), .B(n39500), .Y(n69417) );
  AND2X1 U39943 ( .A(n69406), .B(n69405), .Y(n39280) );
  AND2X1 U39944 ( .A(n65309), .B(n65310), .Y(n39281) );
  OR2X1 U39945 ( .A(n39282), .B(n39283), .Y(n65849) );
  OR2X1 U39946 ( .A(n41375), .B(n65848), .Y(n39282) );
  AND2X1 U39947 ( .A(n66184), .B(n66183), .Y(n39283) );
  AND2X1 U39948 ( .A(n69293), .B(n43585), .Y(n39284) );
  INVX1 U39949 ( .A(n39284), .Y(n69839) );
  OR2X1 U39950 ( .A(n39285), .B(n39286), .Y(n70856) );
  AND2X1 U39951 ( .A(n43544), .B(n70544), .Y(n39285) );
  AND2X1 U39952 ( .A(n70547), .B(n70546), .Y(n39286) );
  OR2X1 U39953 ( .A(n39287), .B(n39288), .Y(n70470) );
  AND2X1 U39954 ( .A(n38154), .B(n43646), .Y(n39287) );
  AND2X1 U39955 ( .A(n69919), .B(n69918), .Y(n39288) );
  NOR2X1 U39956 ( .A(n39290), .B(n39291), .Y(n39289) );
  INVX1 U39957 ( .A(n39289), .Y(n61916) );
  AND2X1 U39958 ( .A(n61913), .B(n61914), .Y(n39290) );
  AND2X1 U39959 ( .A(n42050), .B(n61915), .Y(n39291) );
  NOR2X1 U39960 ( .A(n39293), .B(n39294), .Y(n39292) );
  INVX1 U39961 ( .A(n39292), .Y(n67539) );
  AND2X1 U39962 ( .A(n37417), .B(n66971), .Y(n39293) );
  AND2X1 U39963 ( .A(n37417), .B(n66972), .Y(n39294) );
  OR2X1 U39964 ( .A(n70557), .B(n39295), .Y(n70556) );
  INVX1 U39965 ( .A(n43623), .Y(n39295) );
  AND2X1 U39966 ( .A(n62877), .B(n41083), .Y(n39296) );
  NAND2X1 U39967 ( .A(n67674), .B(n67673), .Y(n39297) );
  AND2X1 U39968 ( .A(n39297), .B(n39298), .Y(n68467) );
  AND2X1 U39969 ( .A(n39299), .B(n67675), .Y(n39298) );
  INVX1 U39970 ( .A(n43617), .Y(n39299) );
  OR2X1 U39971 ( .A(n69304), .B(n43616), .Y(n69633) );
  AND2X1 U39972 ( .A(n66483), .B(n66968), .Y(n39300) );
  INVX1 U39973 ( .A(n39300), .Y(n66852) );
  OR2X1 U39974 ( .A(n39301), .B(n69878), .Y(n69920) );
  INVX1 U39975 ( .A(n43642), .Y(n39301) );
  NOR2X1 U39976 ( .A(n39303), .B(n39304), .Y(n39302) );
  INVX1 U39977 ( .A(n39302), .Y(n62811) );
  AND2X1 U39978 ( .A(n62571), .B(n62570), .Y(n39303) );
  AND2X1 U39979 ( .A(n42119), .B(n62574), .Y(n39304) );
  OR2X1 U39980 ( .A(n62513), .B(n62512), .Y(n39305) );
  XOR2X1 U39981 ( .A(n69486), .B(n69485), .Y(n39306) );
  OR2X1 U39982 ( .A(n39307), .B(n39927), .Y(n70131) );
  AND2X1 U39983 ( .A(n41182), .B(n70125), .Y(n39307) );
  NOR2X1 U39984 ( .A(n39308), .B(n71722), .Y(n40367) );
  NAND2X1 U39985 ( .A(n43514), .B(n71705), .Y(n39308) );
  XOR2X1 U39986 ( .A(n66488), .B(n39845), .Y(n39309) );
  XNOR2X1 U39987 ( .A(n66984), .B(n40737), .Y(n39310) );
  OR2X1 U39988 ( .A(n39311), .B(n39312), .Y(n63511) );
  OR2X1 U39989 ( .A(n63297), .B(n63296), .Y(n39311) );
  AND2X1 U39990 ( .A(n63298), .B(n38635), .Y(n39312) );
  NOR2X1 U39991 ( .A(n39314), .B(n39315), .Y(n39313) );
  AND2X1 U39992 ( .A(n59665), .B(n59853), .Y(n39314) );
  AND2X1 U39993 ( .A(n59852), .B(n59666), .Y(n39315) );
  AND2X1 U39994 ( .A(n39316), .B(n39317), .Y(n65992) );
  OR2X1 U39995 ( .A(n65618), .B(n65617), .Y(n39316) );
  AND2X1 U39996 ( .A(n41274), .B(n68876), .Y(n68879) );
  AND2X1 U39997 ( .A(n38947), .B(n42770), .Y(n39318) );
  AND2X1 U39998 ( .A(n38947), .B(n42770), .Y(n39319) );
  OR2X1 U39999 ( .A(n42997), .B(n69311), .Y(n69310) );
  NOR2X1 U40000 ( .A(n39321), .B(n38363), .Y(n39320) );
  INVX1 U40001 ( .A(n39320), .Y(n65901) );
  AND2X1 U40002 ( .A(n64599), .B(n64598), .Y(n39321) );
  INVX1 U40003 ( .A(n42019), .Y(n39322) );
  AND2X1 U40004 ( .A(n37925), .B(n61427), .Y(n39323) );
  OR2X1 U40005 ( .A(n39324), .B(n39325), .Y(n67807) );
  INVX1 U40006 ( .A(n67321), .Y(n39324) );
  AND2X1 U40007 ( .A(n67320), .B(n67319), .Y(n39325) );
  OR2X1 U40008 ( .A(n39326), .B(n39327), .Y(n70838) );
  INVX1 U40009 ( .A(n70837), .Y(n39326) );
  OR2X1 U40010 ( .A(n39328), .B(n39329), .Y(n72703) );
  OR2X1 U40011 ( .A(n72691), .B(n72690), .Y(n39328) );
  AND2X1 U40012 ( .A(n72695), .B(n72694), .Y(n39329) );
  OR2X1 U40013 ( .A(n37368), .B(n39330), .Y(n68427) );
  AND2X1 U40014 ( .A(n68421), .B(n68083), .Y(n39330) );
  AND2X1 U40015 ( .A(n70209), .B(n43658), .Y(n39331) );
  AND2X1 U40016 ( .A(n68324), .B(n68086), .Y(n39332) );
  INVX1 U40017 ( .A(n39332), .Y(n68149) );
  AND2X1 U40018 ( .A(n40405), .B(n36642), .Y(n70839) );
  INVX1 U40019 ( .A(n39473), .Y(n39333) );
  OR2X1 U40020 ( .A(n39334), .B(n39474), .Y(n61931) );
  NAND2X1 U40021 ( .A(n39333), .B(n61930), .Y(n39334) );
  XOR2X1 U40022 ( .A(n68507), .B(n68205), .Y(n68567) );
  OR2X1 U40023 ( .A(n42832), .B(n42831), .Y(n39335) );
  XOR2X1 U40024 ( .A(n71104), .B(n70835), .Y(n71157) );
  AND2X1 U40025 ( .A(n60695), .B(n60700), .Y(n39336) );
  OR2X1 U40026 ( .A(n39337), .B(n59232), .Y(n59685) );
  AND2X1 U40027 ( .A(n59146), .B(n59678), .Y(n39337) );
  NOR2X1 U40028 ( .A(n39339), .B(n39340), .Y(n39338) );
  INVX1 U40029 ( .A(n38784), .Y(n64362) );
  AND2X1 U40030 ( .A(n64216), .B(n64215), .Y(n39339) );
  AND2X1 U40031 ( .A(n64218), .B(n64217), .Y(n39340) );
  AND2X1 U40032 ( .A(n60580), .B(n60581), .Y(n39341) );
  XOR2X1 U40033 ( .A(n40191), .B(n39434), .Y(n39342) );
  NAND2X1 U40034 ( .A(n41122), .B(n66078), .Y(n39343) );
  NOR2X1 U40035 ( .A(n39345), .B(n39346), .Y(n39344) );
  AND2X1 U40036 ( .A(n39435), .B(n38309), .Y(n39345) );
  AND2X1 U40037 ( .A(n61229), .B(n61228), .Y(n39346) );
  NOR2X1 U40038 ( .A(n39348), .B(n39349), .Y(n39347) );
  INVX1 U40039 ( .A(n39347), .Y(n63487) );
  INVX1 U40040 ( .A(n38896), .Y(n39348) );
  AND2X1 U40041 ( .A(n63319), .B(n63318), .Y(n39349) );
  OR2X1 U40042 ( .A(n39350), .B(n40561), .Y(n40713) );
  OR2X1 U40043 ( .A(n71148), .B(n71147), .Y(n39350) );
  OR2X1 U40044 ( .A(n39351), .B(n39352), .Y(n64297) );
  OR2X1 U40045 ( .A(n38547), .B(n64299), .Y(n39351) );
  AND2X1 U40046 ( .A(n64247), .B(n44009), .Y(n39352) );
  OR2X1 U40047 ( .A(n39191), .B(n40526), .Y(n39353) );
  OR2X1 U40048 ( .A(n39191), .B(n40526), .Y(n39354) );
  OR2X1 U40049 ( .A(n39355), .B(n39356), .Y(n64198) );
  OR2X1 U40050 ( .A(n63867), .B(n64189), .Y(n39355) );
  AND2X1 U40051 ( .A(n63868), .B(n64192), .Y(n39356) );
  AND2X1 U40052 ( .A(n68907), .B(n69527), .Y(n39357) );
  AND2X1 U40053 ( .A(n42376), .B(n62895), .Y(n39358) );
  INVX1 U40054 ( .A(n39358), .Y(n73384) );
  OR2X1 U40055 ( .A(n39359), .B(n39360), .Y(n63608) );
  AND2X1 U40056 ( .A(n63615), .B(n63363), .Y(n39359) );
  AND2X1 U40057 ( .A(n63364), .B(n63612), .Y(n39360) );
  NOR2X1 U40058 ( .A(n59607), .B(n59606), .Y(n39361) );
  AND2X1 U40059 ( .A(n40743), .B(n40744), .Y(n39362) );
  OR2X1 U40060 ( .A(n61696), .B(n61792), .Y(n61697) );
  AND2X1 U40061 ( .A(n2935), .B(n40423), .Y(n45246) );
  OR2X1 U40062 ( .A(n67865), .B(n40302), .Y(n39363) );
  OR2X1 U40063 ( .A(n39954), .B(n39366), .Y(n39364) );
  AND2X1 U40064 ( .A(n39364), .B(n39365), .Y(n69846) );
  OR2X1 U40065 ( .A(n39284), .B(n69299), .Y(n39365) );
  OR2X1 U40066 ( .A(n39953), .B(n39284), .Y(n39366) );
  AND2X1 U40067 ( .A(n68259), .B(n68258), .Y(n39367) );
  NAND2X1 U40068 ( .A(n64734), .B(n39371), .Y(n39368) );
  AND2X1 U40069 ( .A(n39368), .B(n39369), .Y(n65364) );
  OR2X1 U40070 ( .A(n39370), .B(n64736), .Y(n39369) );
  INVX1 U40071 ( .A(n65036), .Y(n39370) );
  AND2X1 U40072 ( .A(n41508), .B(n65036), .Y(n39371) );
  OR2X1 U40073 ( .A(n39374), .B(n39373), .Y(n64631) );
  INVX1 U40074 ( .A(n64508), .Y(n39373) );
  NAND2X1 U40075 ( .A(n41309), .B(n64507), .Y(n39374) );
  NOR2X1 U40076 ( .A(n39376), .B(n39377), .Y(n39375) );
  AND2X1 U40077 ( .A(n61466), .B(n61398), .Y(n39376) );
  AND2X1 U40078 ( .A(n41916), .B(n61400), .Y(n39377) );
  NOR2X1 U40079 ( .A(n39587), .B(n39588), .Y(n39378) );
  AND2X1 U40080 ( .A(n43581), .B(n67856), .Y(n39379) );
  OR2X1 U40081 ( .A(n60560), .B(n60559), .Y(n60561) );
  NOR2X1 U40082 ( .A(n63757), .B(n64205), .Y(n39380) );
  INVX1 U40083 ( .A(n39380), .Y(n64213) );
  OR2X1 U40084 ( .A(n39381), .B(n65338), .Y(n65326) );
  INVX1 U40085 ( .A(n65312), .Y(n39381) );
  OR2X1 U40086 ( .A(n38541), .B(n63986), .Y(n39382) );
  AND2X1 U40087 ( .A(n63987), .B(n44018), .Y(n39383) );
  AND2X1 U40088 ( .A(n65312), .B(n65311), .Y(n39384) );
  INVX1 U40089 ( .A(n39384), .Y(n65327) );
  NAND2X1 U40090 ( .A(n39386), .B(n60941), .Y(n39385) );
  OR2X1 U40091 ( .A(n60937), .B(n60939), .Y(n39386) );
  NOR2X1 U40092 ( .A(n39388), .B(n39389), .Y(n39387) );
  INVX1 U40093 ( .A(n39042), .Y(n60887) );
  AND2X1 U40094 ( .A(n60736), .B(n60735), .Y(n39388) );
  AND2X1 U40095 ( .A(n41977), .B(n60747), .Y(n39389) );
  OR2X1 U40096 ( .A(n60759), .B(n39390), .Y(n60550) );
  AND2X1 U40097 ( .A(n38268), .B(n60549), .Y(n39390) );
  AND2X1 U40098 ( .A(n68567), .B(n43550), .Y(n39391) );
  AND2X1 U40099 ( .A(n71422), .B(n41454), .Y(n72099) );
  AND2X1 U40100 ( .A(n59816), .B(n59815), .Y(n39392) );
  NOR2X1 U40101 ( .A(n39523), .B(n39524), .Y(n39393) );
  OR2X1 U40102 ( .A(n39394), .B(n39395), .Y(n64578) );
  AND2X1 U40103 ( .A(n43507), .B(n64287), .Y(n39394) );
  AND2X1 U40104 ( .A(n64289), .B(n64288), .Y(n39395) );
  AND2X1 U40105 ( .A(n68149), .B(n68151), .Y(n39396) );
  NOR2X1 U40106 ( .A(n39398), .B(n39399), .Y(n39397) );
  AND2X1 U40107 ( .A(n60089), .B(n60040), .Y(n39398) );
  AND2X1 U40108 ( .A(n41895), .B(n60042), .Y(n39399) );
  NOR2X1 U40109 ( .A(n39401), .B(n39402), .Y(n39400) );
  AND2X1 U40110 ( .A(n61625), .B(n61535), .Y(n39401) );
  AND2X1 U40111 ( .A(n41899), .B(n61537), .Y(n39402) );
  OR2X1 U40112 ( .A(n39403), .B(n39404), .Y(n61726) );
  INVX1 U40113 ( .A(n42008), .Y(n39403) );
  OR2X1 U40114 ( .A(n40562), .B(n39405), .Y(n71114) );
  AND2X1 U40115 ( .A(n70779), .B(n70840), .Y(n39405) );
  INVX1 U40116 ( .A(n42018), .Y(n39406) );
  AND2X1 U40117 ( .A(n61767), .B(n61729), .Y(n39407) );
  OR2X1 U40118 ( .A(n37366), .B(n39408), .Y(n64667) );
  AND2X1 U40119 ( .A(n64663), .B(n64323), .Y(n39408) );
  OR2X1 U40120 ( .A(n43748), .B(n36719), .Y(n59995) );
  OR2X1 U40121 ( .A(n39643), .B(n39644), .Y(n39409) );
  OR2X1 U40122 ( .A(n39410), .B(n39411), .Y(n63615) );
  OR2X1 U40123 ( .A(n63364), .B(n63354), .Y(n39410) );
  OR2X1 U40124 ( .A(n37380), .B(n63357), .Y(n39411) );
  NOR2X1 U40125 ( .A(n39413), .B(n37374), .Y(n39412) );
  INVX1 U40126 ( .A(n39412), .Y(n71757) );
  OR2X1 U40127 ( .A(n41047), .B(n40944), .Y(n39413) );
  XOR2X1 U40128 ( .A(n65867), .B(n40077), .Y(n39414) );
  AND2X1 U40129 ( .A(n63481), .B(n39415), .Y(n63479) );
  INVX1 U40130 ( .A(n63477), .Y(n39415) );
  INVX1 U40131 ( .A(n39538), .Y(n39416) );
  OR2X1 U40132 ( .A(n39538), .B(n39539), .Y(n39417) );
  INVX1 U40133 ( .A(n39417), .Y(n39537) );
  OR2X1 U40134 ( .A(n39418), .B(n39419), .Y(n71131) );
  OR2X1 U40135 ( .A(n70184), .B(n70190), .Y(n39418) );
  AND2X1 U40136 ( .A(n70185), .B(n70186), .Y(n39419) );
  OR2X1 U40137 ( .A(n61203), .B(n40496), .Y(n61204) );
  OR2X1 U40138 ( .A(n39956), .B(n39957), .Y(n39420) );
  AND2X1 U40139 ( .A(n59397), .B(n59396), .Y(n39421) );
  INVX1 U40140 ( .A(n62421), .Y(n39422) );
  OR2X1 U40141 ( .A(n39424), .B(n39425), .Y(n61714) );
  INVX1 U40142 ( .A(n41974), .Y(n39424) );
  AND2X1 U40143 ( .A(n36413), .B(n61713), .Y(n39425) );
  NOR2X1 U40144 ( .A(n64353), .B(n64352), .Y(n39426) );
  AND2X1 U40145 ( .A(n40455), .B(n36565), .Y(n39427) );
  AND2X1 U40146 ( .A(n41999), .B(n39428), .Y(n41535) );
  NAND2X1 U40147 ( .A(n64681), .B(n64680), .Y(n39428) );
  AND2X1 U40148 ( .A(n61271), .B(n61276), .Y(n39429) );
  XNOR2X1 U40149 ( .A(n72686), .B(n39430), .Y(n72699) );
  XOR2X1 U40150 ( .A(n72096), .B(n72692), .Y(n39430) );
  OR2X1 U40151 ( .A(n39657), .B(n39658), .Y(n39431) );
  OR2X1 U40152 ( .A(n39432), .B(n39433), .Y(n65005) );
  OR2X1 U40153 ( .A(n64813), .B(n40947), .Y(n39432) );
  AND2X1 U40154 ( .A(n64814), .B(n38696), .Y(n39433) );
  XOR2X1 U40155 ( .A(n40191), .B(n39434), .Y(n69313) );
  XOR2X1 U40156 ( .A(n68758), .B(n39159), .Y(n39434) );
  OR2X1 U40157 ( .A(n39860), .B(n39861), .Y(n39435) );
  NOR2X1 U40158 ( .A(n39437), .B(n39438), .Y(n39436) );
  INVX1 U40159 ( .A(n39436), .Y(n67697) );
  OR2X1 U40160 ( .A(n67687), .B(n67686), .Y(n39437) );
  AND2X1 U40161 ( .A(n67692), .B(n67691), .Y(n39438) );
  OR2X1 U40162 ( .A(n39439), .B(n39440), .Y(n62515) );
  OR2X1 U40163 ( .A(n61249), .B(n61248), .Y(n39439) );
  AND2X1 U40164 ( .A(n61250), .B(n61263), .Y(n39440) );
  NOR2X1 U40165 ( .A(n39442), .B(n39443), .Y(n39441) );
  INVX1 U40166 ( .A(n38149), .Y(n60851) );
  AND2X1 U40167 ( .A(n61322), .B(n60847), .Y(n39442) );
  AND2X1 U40168 ( .A(n41921), .B(n60849), .Y(n39443) );
  OR2X1 U40169 ( .A(n66761), .B(n66764), .Y(n67118) );
  NAND2X1 U40170 ( .A(n37318), .B(n39185), .Y(n39444) );
  OR2X1 U40171 ( .A(n39445), .B(n40287), .Y(n66792) );
  AND2X1 U40172 ( .A(n41127), .B(n67339), .Y(n39445) );
  OR2X1 U40173 ( .A(n67886), .B(n39446), .Y(n67885) );
  INVX1 U40174 ( .A(n43648), .Y(n39446) );
  OR2X1 U40175 ( .A(n39448), .B(n39447), .Y(n67860) );
  INVX1 U40176 ( .A(n67863), .Y(n39447) );
  AND2X1 U40177 ( .A(n67289), .B(n67288), .Y(n39448) );
  AND2X1 U40178 ( .A(opcode_opcode_w[23]), .B(opcode_opcode_w[24]), .Y(n39449)
         );
  INVX1 U40179 ( .A(n39449), .Y(n39809) );
  OR2X1 U40180 ( .A(n40244), .B(n40245), .Y(n39450) );
  AND2X1 U40181 ( .A(n65816), .B(n65834), .Y(n39451) );
  OR2X1 U40182 ( .A(n39452), .B(n39453), .Y(n65307) );
  OR2X1 U40183 ( .A(n65137), .B(n65136), .Y(n39452) );
  AND2X1 U40184 ( .A(n65140), .B(n65139), .Y(n39453) );
  NOR2X1 U40185 ( .A(n39455), .B(n39456), .Y(n39454) );
  INVX1 U40186 ( .A(n39454), .Y(n60788) );
  AND2X1 U40187 ( .A(n60790), .B(n60487), .Y(n39455) );
  AND2X1 U40188 ( .A(n41841), .B(n60489), .Y(n39456) );
  OR2X1 U40189 ( .A(n39457), .B(n40336), .Y(n67141) );
  AND2X1 U40190 ( .A(n66079), .B(n66081), .Y(n39457) );
  NOR2X1 U40191 ( .A(n39459), .B(n39460), .Y(n39458) );
  AND2X1 U40192 ( .A(n60143), .B(n60141), .Y(n39459) );
  AND2X1 U40193 ( .A(n41847), .B(n60016), .Y(n39460) );
  OR2X1 U40194 ( .A(n67024), .B(n67025), .Y(n39461) );
  INVX1 U40195 ( .A(n39461), .Y(n39971) );
  OR2X1 U40196 ( .A(n39553), .B(n39554), .Y(n39462) );
  NOR2X1 U40197 ( .A(n39464), .B(n39465), .Y(n39463) );
  AND2X1 U40198 ( .A(n61470), .B(n38167), .Y(n39464) );
  AND2X1 U40199 ( .A(n41893), .B(n61393), .Y(n39465) );
  AND2X1 U40200 ( .A(n68340), .B(n68635), .Y(n39466) );
  OR2X1 U40201 ( .A(n41353), .B(n63740), .Y(n39467) );
  NAND2X1 U40202 ( .A(n41351), .B(n63741), .Y(n39468) );
  XOR2X1 U40203 ( .A(n67546), .B(n42810), .Y(n39469) );
  AND2X1 U40204 ( .A(n40274), .B(n41296), .Y(n39470) );
  OR2X1 U40205 ( .A(n41272), .B(n41276), .Y(n39471) );
  OR2X1 U40206 ( .A(n37887), .B(n36828), .Y(n65239) );
  NOR2X1 U40207 ( .A(n39473), .B(n39474), .Y(n39472) );
  INVX1 U40208 ( .A(n39472), .Y(n61929) );
  AND2X1 U40209 ( .A(n61926), .B(n61927), .Y(n39473) );
  AND2X1 U40210 ( .A(n42081), .B(n61928), .Y(n39474) );
  AND2X1 U40211 ( .A(n41365), .B(n64878), .Y(n39475) );
  OR2X1 U40212 ( .A(n36789), .B(n60364), .Y(n60365) );
  AND2X1 U40213 ( .A(n39476), .B(n39477), .Y(n39655) );
  NAND2X1 U40214 ( .A(n69533), .B(n38388), .Y(n39477) );
  NAND2X1 U40215 ( .A(n63039), .B(n63040), .Y(n39478) );
  NOR2X1 U40216 ( .A(n39480), .B(n39481), .Y(n39479) );
  INVX1 U40217 ( .A(n40985), .Y(n39480) );
  AND2X1 U40218 ( .A(n65013), .B(n65012), .Y(n39481) );
  OR2X1 U40219 ( .A(n40074), .B(n40075), .Y(n39482) );
  AND2X1 U40220 ( .A(n63806), .B(n63805), .Y(n39483) );
  OR2X1 U40221 ( .A(n39484), .B(n39485), .Y(n65956) );
  OR2X1 U40222 ( .A(n65587), .B(n40202), .Y(n39484) );
  AND2X1 U40223 ( .A(n65593), .B(n65592), .Y(n39485) );
  NOR2X1 U40224 ( .A(n39487), .B(n39488), .Y(n39486) );
  INVX1 U40225 ( .A(n39486), .Y(n67465) );
  INVX1 U40226 ( .A(n67479), .Y(n39487) );
  AND2X1 U40227 ( .A(n67324), .B(n41155), .Y(n39488) );
  OR2X1 U40228 ( .A(n39489), .B(n39490), .Y(n68760) );
  INVX1 U40229 ( .A(n41728), .Y(n39489) );
  AND2X1 U40230 ( .A(n68304), .B(n68303), .Y(n39490) );
  NAND2X1 U40231 ( .A(n39493), .B(n39444), .Y(n39491) );
  AND2X1 U40232 ( .A(n39491), .B(n39492), .Y(n64334) );
  OR2X1 U40233 ( .A(n64858), .B(n64023), .Y(n39492) );
  AND2X1 U40234 ( .A(n64020), .B(n64333), .Y(n39493) );
  OR2X1 U40235 ( .A(n60316), .B(n39494), .Y(n60167) );
  NAND2X1 U40236 ( .A(n43653), .B(n69538), .Y(n39495) );
  AND2X1 U40237 ( .A(n68588), .B(n39496), .Y(n68502) );
  NOR2X1 U40238 ( .A(n43562), .B(n68505), .Y(n39496) );
  OR2X1 U40239 ( .A(n39497), .B(n37376), .Y(n68273) );
  OR2X1 U40240 ( .A(n39379), .B(n40201), .Y(n39497) );
  OR2X1 U40241 ( .A(n39498), .B(n39499), .Y(n65970) );
  AND2X1 U40242 ( .A(n43664), .B(n65918), .Y(n39498) );
  AND2X1 U40243 ( .A(n65543), .B(n65919), .Y(n39499) );
  NOR2X1 U40244 ( .A(n69404), .B(n37370), .Y(n39500) );
  INVX1 U40245 ( .A(n39500), .Y(n69407) );
  NOR2X1 U40246 ( .A(n42833), .B(n39701), .Y(n39501) );
  NOR2X1 U40247 ( .A(n42833), .B(n39701), .Y(n39502) );
  AND2X1 U40248 ( .A(n37372), .B(n69493), .Y(n69494) );
  OR2X1 U40249 ( .A(n39503), .B(n39504), .Y(n65100) );
  INVX1 U40250 ( .A(n64716), .Y(n39503) );
  AND2X1 U40251 ( .A(n64467), .B(n64466), .Y(n39504) );
  AND2X1 U40252 ( .A(n61090), .B(n61089), .Y(n39505) );
  OR2X1 U40253 ( .A(n43494), .B(n40589), .Y(n61147) );
  OR2X1 U40254 ( .A(n38664), .B(n63646), .Y(n39506) );
  INVX1 U40255 ( .A(n39506), .Y(n63648) );
  OR2X1 U40256 ( .A(n39507), .B(n39508), .Y(n66570) );
  AND2X1 U40257 ( .A(n43505), .B(n66250), .Y(n39507) );
  AND2X1 U40258 ( .A(n66253), .B(n66252), .Y(n39508) );
  AND2X1 U40259 ( .A(n65714), .B(n39509), .Y(n66090) );
  INVX1 U40260 ( .A(n66088), .Y(n39509) );
  NAND2X1 U40261 ( .A(n66571), .B(n66570), .Y(n39510) );
  XOR2X1 U40262 ( .A(n69877), .B(n41017), .Y(n39511) );
  AND2X1 U40263 ( .A(n68021), .B(n68277), .Y(n39512) );
  OR2X1 U40264 ( .A(n59464), .B(n59437), .Y(n59503) );
  OR2X1 U40265 ( .A(n39513), .B(n37369), .Y(n67053) );
  AND2X1 U40266 ( .A(n67069), .B(n66787), .Y(n39513) );
  INVX1 U40267 ( .A(n39691), .Y(n39514) );
  AND2X1 U40268 ( .A(n67017), .B(n67016), .Y(n39515) );
  INVX1 U40269 ( .A(n39515), .Y(n67319) );
  OR2X1 U40270 ( .A(n40866), .B(n45168), .Y(n46007) );
  OR2X1 U40271 ( .A(n39516), .B(n39517), .Y(n69687) );
  OR2X1 U40272 ( .A(n39500), .B(n41239), .Y(n39516) );
  OR2X1 U40273 ( .A(n69402), .B(n69401), .Y(n39517) );
  NAND2X1 U40274 ( .A(n66925), .B(n39510), .Y(n39518) );
  AND2X1 U40275 ( .A(n66553), .B(n66552), .Y(n39519) );
  AND2X1 U40276 ( .A(n41239), .B(n69417), .Y(n39520) );
  NAND2X1 U40277 ( .A(n68755), .B(n68754), .Y(n39521) );
  NOR2X1 U40278 ( .A(n39523), .B(n39524), .Y(n39522) );
  INVX1 U40279 ( .A(n39393), .Y(n62371) );
  OR2X1 U40280 ( .A(n61115), .B(n61114), .Y(n39523) );
  AND2X1 U40281 ( .A(n61118), .B(n61117), .Y(n39524) );
  INVX1 U40282 ( .A(n43769), .Y(n39525) );
  AND2X1 U40283 ( .A(n39526), .B(n63460), .Y(n64000) );
  OR2X1 U40284 ( .A(n63919), .B(n63918), .Y(n39526) );
  NAND2X1 U40285 ( .A(n47701), .B(n39530), .Y(n39527) );
  AND2X1 U40286 ( .A(n39527), .B(n39528), .Y(n63222) );
  OR2X1 U40287 ( .A(n39529), .B(n42804), .Y(n39528) );
  INVX1 U40288 ( .A(n36783), .Y(n39529) );
  AND2X1 U40289 ( .A(n47702), .B(n36783), .Y(n39530) );
  OR2X1 U40290 ( .A(n38260), .B(n39531), .Y(n64061) );
  AND2X1 U40291 ( .A(n40469), .B(n36777), .Y(n39531) );
  OR2X1 U40292 ( .A(n39532), .B(n39533), .Y(n60565) );
  AND2X1 U40293 ( .A(n60431), .B(n60424), .Y(n39532) );
  AND2X1 U40294 ( .A(n60427), .B(n60426), .Y(n39533) );
  AND2X1 U40295 ( .A(n60399), .B(n39534), .Y(n60402) );
  NOR2X1 U40296 ( .A(n38183), .B(n60401), .Y(n39534) );
  AND2X1 U40297 ( .A(n67306), .B(n67305), .Y(n39535) );
  INVX1 U40298 ( .A(n39535), .Y(n67011) );
  AND2X1 U40299 ( .A(n63378), .B(n63380), .Y(n39536) );
  INVX1 U40300 ( .A(n39536), .Y(n63458) );
  AND2X1 U40301 ( .A(n61284), .B(n61283), .Y(n39538) );
  AND2X1 U40302 ( .A(n61288), .B(n61287), .Y(n39539) );
  OR2X1 U40303 ( .A(n39540), .B(n39541), .Y(n60739) );
  AND2X1 U40304 ( .A(n60416), .B(n60180), .Y(n39540) );
  AND2X1 U40305 ( .A(n41957), .B(n60182), .Y(n39541) );
  AND2X1 U40306 ( .A(n37361), .B(n39542), .Y(n59677) );
  AND2X1 U40307 ( .A(n59676), .B(n59890), .Y(n39542) );
  OR2X1 U40308 ( .A(n63702), .B(n63703), .Y(n63706) );
  NOR2X1 U40309 ( .A(n39544), .B(n39545), .Y(n39543) );
  INVX1 U40310 ( .A(n42183), .Y(n39544) );
  AND2X1 U40311 ( .A(n67312), .B(n67311), .Y(n39545) );
  OR2X1 U40312 ( .A(n36566), .B(n39546), .Y(n64929) );
  AND2X1 U40313 ( .A(n64635), .B(n64634), .Y(n39546) );
  NOR2X1 U40314 ( .A(n39548), .B(n39549), .Y(n39547) );
  AND2X1 U40315 ( .A(n61389), .B(n61390), .Y(n39548) );
  AND2X1 U40316 ( .A(n41884), .B(n61391), .Y(n39549) );
  OR2X1 U40317 ( .A(n39550), .B(n39551), .Y(n60081) );
  AND2X1 U40318 ( .A(n60053), .B(n60169), .Y(n39550) );
  AND2X1 U40319 ( .A(n41923), .B(n60056), .Y(n39551) );
  NOR2X1 U40320 ( .A(n39553), .B(n39554), .Y(n39552) );
  AND2X1 U40321 ( .A(n60283), .B(n60284), .Y(n39553) );
  AND2X1 U40322 ( .A(n60287), .B(n60288), .Y(n39554) );
  NOR2X1 U40323 ( .A(n69656), .B(n39556), .Y(n39555) );
  INVX1 U40324 ( .A(n39555), .Y(n69646) );
  INVX1 U40325 ( .A(n42998), .Y(n39556) );
  AND2X1 U40326 ( .A(n66766), .B(n67118), .Y(n39557) );
  OR2X1 U40327 ( .A(n39558), .B(n39559), .Y(n63911) );
  INVX1 U40328 ( .A(n63907), .Y(n39558) );
  AND2X1 U40329 ( .A(n63906), .B(n63905), .Y(n39559) );
  NOR2X1 U40330 ( .A(n39561), .B(n39562), .Y(n39560) );
  INVX1 U40331 ( .A(n39560), .Y(n60134) );
  AND2X1 U40332 ( .A(n37395), .B(n60007), .Y(n39561) );
  AND2X1 U40333 ( .A(n41807), .B(n60008), .Y(n39562) );
  AND2X1 U40334 ( .A(n62400), .B(n62399), .Y(n39563) );
  OR2X1 U40335 ( .A(n71151), .B(n40262), .Y(n71696) );
  OR2X1 U40336 ( .A(n39564), .B(n39565), .Y(n63640) );
  OR2X1 U40337 ( .A(n63631), .B(n63630), .Y(n39564) );
  AND2X1 U40338 ( .A(n63638), .B(n63637), .Y(n39565) );
  NOR2X1 U40339 ( .A(n37387), .B(n39567), .Y(n39566) );
  NAND2X1 U40340 ( .A(n68300), .B(n68301), .Y(n39567) );
  AND2X1 U40341 ( .A(n63133), .B(n63132), .Y(n39568) );
  AND2X1 U40342 ( .A(n60917), .B(n60916), .Y(n39569) );
  INVX1 U40343 ( .A(n39569), .Y(n60911) );
  XOR2X1 U40344 ( .A(n68753), .B(n40980), .Y(n39570) );
  AND2X1 U40345 ( .A(n60620), .B(n60623), .Y(n39571) );
  INVX1 U40346 ( .A(n40521), .Y(n39572) );
  AND2X1 U40347 ( .A(n65034), .B(n65033), .Y(n39573) );
  OR2X1 U40348 ( .A(n39574), .B(n39575), .Y(n59454) );
  AND2X1 U40349 ( .A(n59447), .B(n59460), .Y(n39574) );
  AND2X1 U40350 ( .A(n59450), .B(n59449), .Y(n39575) );
  NOR2X1 U40351 ( .A(n40144), .B(n40145), .Y(n39576) );
  NAND2X1 U40352 ( .A(n69891), .B(n39579), .Y(n39577) );
  AND2X1 U40353 ( .A(n39577), .B(n39578), .Y(n70166) );
  OR2X1 U40354 ( .A(n41274), .B(n70165), .Y(n39578) );
  AND2X1 U40355 ( .A(n39241), .B(n43529), .Y(n39579) );
  AND2X1 U40356 ( .A(n70485), .B(n70484), .Y(n39580) );
  OR2X1 U40357 ( .A(n38257), .B(n62873), .Y(n63167) );
  AND2X1 U40358 ( .A(n71226), .B(n71211), .Y(n39581) );
  INVX1 U40359 ( .A(n39581), .Y(n71214) );
  NAND2X1 U40360 ( .A(n40449), .B(n40018), .Y(n39582) );
  NAND2X1 U40361 ( .A(n40449), .B(n40018), .Y(n39583) );
  NOR2X1 U40362 ( .A(n42789), .B(n42669), .Y(n39584) );
  INVX1 U40363 ( .A(n39584), .Y(n48116) );
  AND2X1 U40364 ( .A(n40152), .B(n39585), .Y(n45450) );
  NOR2X1 U40365 ( .A(n42703), .B(n45449), .Y(n39585) );
  NOR2X1 U40366 ( .A(n39587), .B(n39588), .Y(n39586) );
  INVX1 U40367 ( .A(n39378), .Y(n67303) );
  OR2X1 U40368 ( .A(n66989), .B(n66988), .Y(n39587) );
  AND2X1 U40369 ( .A(n66995), .B(n66994), .Y(n39588) );
  OR2X1 U40370 ( .A(n39589), .B(n39590), .Y(n65828) );
  OR2X1 U40371 ( .A(n65332), .B(n65331), .Y(n39589) );
  OR2X1 U40372 ( .A(n65344), .B(n65343), .Y(n39590) );
  OR2X1 U40373 ( .A(n39233), .B(n39591), .Y(n45529) );
  OR2X1 U40374 ( .A(n46206), .B(n37048), .Y(n39591) );
  NOR2X1 U40375 ( .A(n39593), .B(n39594), .Y(n39592) );
  AND2X1 U40376 ( .A(n39638), .B(n59594), .Y(n39593) );
  AND2X1 U40377 ( .A(n59588), .B(n59589), .Y(n39594) );
  OR2X1 U40378 ( .A(n39226), .B(n39595), .Y(n69554) );
  OR2X1 U40379 ( .A(n39596), .B(n39597), .Y(n64217) );
  OR2X1 U40380 ( .A(n39380), .B(n63759), .Y(n39596) );
  AND2X1 U40381 ( .A(n63761), .B(n63760), .Y(n39597) );
  OR2X1 U40382 ( .A(n39598), .B(n39599), .Y(n47338) );
  OR2X1 U40383 ( .A(n47331), .B(n47330), .Y(n39598) );
  OR2X1 U40384 ( .A(n47337), .B(n47336), .Y(n39599) );
  AND2X1 U40385 ( .A(n39600), .B(n61263), .Y(n61248) );
  INVX1 U40386 ( .A(n42841), .Y(n39600) );
  NOR2X1 U40387 ( .A(n39602), .B(n39603), .Y(n39601) );
  INVX1 U40388 ( .A(n39601), .Y(n60485) );
  AND2X1 U40389 ( .A(n60456), .B(n60356), .Y(n39602) );
  AND2X1 U40390 ( .A(n41813), .B(n60358), .Y(n39603) );
  AND2X1 U40391 ( .A(n60950), .B(n42367), .Y(n39604) );
  INVX1 U40392 ( .A(n39604), .Y(n60959) );
  OR2X1 U40393 ( .A(n39606), .B(n39605), .Y(n66308) );
  INVX1 U40394 ( .A(n66304), .Y(n39605) );
  OR2X1 U40395 ( .A(n41645), .B(n41618), .Y(n39606) );
  OR2X1 U40396 ( .A(n40265), .B(n40266), .Y(n39607) );
  OR2X1 U40397 ( .A(n39609), .B(n39608), .Y(n66318) );
  INVX1 U40398 ( .A(n66316), .Y(n39608) );
  OR2X1 U40399 ( .A(n40978), .B(n40981), .Y(n39609) );
  OR2X1 U40400 ( .A(n39610), .B(n39611), .Y(n60960) );
  OR2X1 U40401 ( .A(n45463), .B(n45462), .Y(n39610) );
  AND2X1 U40402 ( .A(n61188), .B(n45519), .Y(n39611) );
  AND2X1 U40403 ( .A(n45307), .B(n45306), .Y(n39612) );
  NAND2X1 U40404 ( .A(n65060), .B(n65067), .Y(n39613) );
  NOR2X1 U40405 ( .A(n39615), .B(n39616), .Y(n39614) );
  OR2X1 U40406 ( .A(n60596), .B(n60595), .Y(n39615) );
  AND2X1 U40407 ( .A(n36788), .B(n60597), .Y(n39616) );
  NOR2X1 U40408 ( .A(n39618), .B(n39619), .Y(n39617) );
  AND2X1 U40409 ( .A(n59880), .B(n40121), .Y(n39618) );
  NOR2X1 U40410 ( .A(n42816), .B(n59881), .Y(n39619) );
  NOR2X1 U40411 ( .A(n42737), .B(n47965), .Y(n39620) );
  INVX1 U40412 ( .A(n39620), .Y(n47636) );
  AND2X1 U40413 ( .A(n62940), .B(n62939), .Y(n39621) );
  OR2X1 U40414 ( .A(n39622), .B(n39623), .Y(n65834) );
  INVX1 U40415 ( .A(n65323), .Y(n39622) );
  AND2X1 U40416 ( .A(n65322), .B(n65321), .Y(n39623) );
  OR2X1 U40417 ( .A(n39624), .B(n39633), .Y(n67850) );
  OR2X1 U40418 ( .A(n67539), .B(n67538), .Y(n39624) );
  OR2X1 U40419 ( .A(n39625), .B(n38395), .Y(n59474) );
  INVX1 U40420 ( .A(n40390), .Y(n39625) );
  OR2X1 U40421 ( .A(n60768), .B(n37400), .Y(n60528) );
  INVX1 U40422 ( .A(n39626), .Y(n62659) );
  INVX1 U40423 ( .A(n42063), .Y(n39627) );
  AND2X1 U40424 ( .A(n36556), .B(n61583), .Y(n39628) );
  OR2X1 U40425 ( .A(n39629), .B(n68585), .Y(n67989) );
  INVX1 U40426 ( .A(n43561), .Y(n39629) );
  NOR2X1 U40427 ( .A(n42737), .B(n39882), .Y(n39630) );
  INVX1 U40428 ( .A(n39630), .Y(n47625) );
  AND2X1 U40429 ( .A(n65878), .B(n65277), .Y(n39631) );
  AND2X1 U40430 ( .A(n60001), .B(n60000), .Y(n39632) );
  AND2X1 U40431 ( .A(n66973), .B(n66963), .Y(n39633) );
  OR2X1 U40432 ( .A(n39814), .B(n39815), .Y(n39634) );
  AND2X1 U40433 ( .A(n43577), .B(n67663), .Y(n39635) );
  INVX1 U40434 ( .A(n39635), .Y(n67999) );
  AND2X1 U40435 ( .A(n63475), .B(n63741), .Y(n39636) );
  AND2X1 U40436 ( .A(n43545), .B(n67642), .Y(n39637) );
  OR2X1 U40437 ( .A(n39763), .B(n39764), .Y(n39638) );
  INVX1 U40438 ( .A(n42814), .Y(n39639) );
  INVX1 U40439 ( .A(n39639), .Y(n39640) );
  AND2X1 U40440 ( .A(n60957), .B(n60956), .Y(n39641) );
  NOR2X1 U40441 ( .A(n39643), .B(n39644), .Y(n39642) );
  AND2X1 U40442 ( .A(n61621), .B(n61542), .Y(n39643) );
  AND2X1 U40443 ( .A(n41920), .B(n61544), .Y(n39644) );
  INVX1 U40444 ( .A(n49605), .Y(n39645) );
  NOR2X1 U40445 ( .A(n40003), .B(n40004), .Y(n39646) );
  AND2X1 U40446 ( .A(n66315), .B(n66841), .Y(n66313) );
  NAND2X1 U40447 ( .A(n44988), .B(n42724), .Y(n39647) );
  AND2X1 U40448 ( .A(n60123), .B(n60124), .Y(n39648) );
  AND2X1 U40449 ( .A(n41785), .B(n60003), .Y(n39649) );
  AND2X1 U40450 ( .A(n60952), .B(n60951), .Y(n39650) );
  OR2X1 U40451 ( .A(n39651), .B(n39652), .Y(n59147) );
  OR2X1 U40452 ( .A(n46417), .B(n46416), .Y(n39651) );
  AND2X1 U40453 ( .A(n40490), .B(n46457), .Y(n39652) );
  INVX1 U40454 ( .A(n43610), .Y(n39653) );
  OR2X1 U40455 ( .A(n45199), .B(n46927), .Y(n39654) );
  INVX1 U40456 ( .A(n39655), .Y(n69587) );
  NOR2X1 U40457 ( .A(n39657), .B(n39658), .Y(n39656) );
  OR2X1 U40458 ( .A(n63754), .B(n63753), .Y(n39657) );
  AND2X1 U40459 ( .A(n63756), .B(n63755), .Y(n39658) );
  OR2X1 U40460 ( .A(n39741), .B(n39742), .Y(n39659) );
  OR2X1 U40461 ( .A(n39660), .B(n39661), .Y(n71239) );
  OR2X1 U40462 ( .A(n70919), .B(n70918), .Y(n39660) );
  AND2X1 U40463 ( .A(n70922), .B(n70921), .Y(n39661) );
  AND2X1 U40464 ( .A(n39662), .B(n39663), .Y(n65985) );
  AND2X1 U40465 ( .A(n65976), .B(n65975), .Y(n39662) );
  AND2X1 U40466 ( .A(n65980), .B(n43560), .Y(n39663) );
  AND2X1 U40467 ( .A(n67550), .B(n39664), .Y(n67552) );
  AND2X1 U40468 ( .A(n67549), .B(n39665), .Y(n39664) );
  INVX1 U40469 ( .A(n43586), .Y(n39665) );
  NOR2X1 U40470 ( .A(n39667), .B(n39668), .Y(n39666) );
  AND2X1 U40471 ( .A(n61300), .B(n37394), .Y(n39667) );
  AND2X1 U40472 ( .A(n42039), .B(n61093), .Y(n39668) );
  AND2X1 U40473 ( .A(n42794), .B(n42666), .Y(n39669) );
  AND2X1 U40474 ( .A(n66533), .B(n43649), .Y(n39670) );
  INVX1 U40475 ( .A(n39670), .Y(n66590) );
  OR2X1 U40476 ( .A(n39671), .B(n39672), .Y(n67972) );
  AND2X1 U40477 ( .A(n67638), .B(n43550), .Y(n39671) );
  AND2X1 U40478 ( .A(n67645), .B(n67644), .Y(n39672) );
  OR2X1 U40479 ( .A(n39673), .B(n39674), .Y(n66963) );
  OR2X1 U40480 ( .A(n66639), .B(n66638), .Y(n39673) );
  AND2X1 U40481 ( .A(n66972), .B(n66964), .Y(n39674) );
  NOR2X1 U40482 ( .A(n39676), .B(n39677), .Y(n39675) );
  INVX1 U40483 ( .A(n39675), .Y(n60833) );
  AND2X1 U40484 ( .A(n60830), .B(n60831), .Y(n39676) );
  AND2X1 U40485 ( .A(n41857), .B(n60832), .Y(n39677) );
  OR2X1 U40486 ( .A(n39874), .B(n39875), .Y(n39678) );
  NAND2X1 U40487 ( .A(n67885), .B(n67884), .Y(n39679) );
  NAND2X1 U40488 ( .A(n40157), .B(n40148), .Y(n39680) );
  NAND2X1 U40489 ( .A(n38856), .B(n60617), .Y(n39681) );
  AND2X1 U40490 ( .A(n60233), .B(n60937), .Y(n39682) );
  OR2X1 U40491 ( .A(n39683), .B(n39684), .Y(n60961) );
  OR2X1 U40492 ( .A(n45542), .B(n45541), .Y(n39684) );
  NOR2X1 U40493 ( .A(n39686), .B(n39687), .Y(n39685) );
  INVX1 U40494 ( .A(n39685), .Y(n60332) );
  AND2X1 U40495 ( .A(n60361), .B(n60362), .Y(n39686) );
  AND2X1 U40496 ( .A(n41824), .B(n60132), .Y(n39687) );
  OR2X1 U40497 ( .A(n39831), .B(n39832), .Y(n39688) );
  NAND2X1 U40498 ( .A(n36703), .B(n39692), .Y(n39689) );
  AND2X1 U40499 ( .A(n39689), .B(n39690), .Y(n65619) );
  OR2X1 U40500 ( .A(n39691), .B(n64944), .Y(n39690) );
  INVX1 U40501 ( .A(n65615), .Y(n39691) );
  AND2X1 U40502 ( .A(n65615), .B(n64932), .Y(n39692) );
  OR2X1 U40503 ( .A(n39693), .B(n37359), .Y(n64874) );
  AND2X1 U40504 ( .A(n65187), .B(n64523), .Y(n39693) );
  OR2X1 U40505 ( .A(n40612), .B(n40613), .Y(n39694) );
  OR2X1 U40506 ( .A(n39770), .B(n45168), .Y(n46236) );
  NOR2X1 U40507 ( .A(n39696), .B(n39697), .Y(n39695) );
  AND2X1 U40508 ( .A(n60290), .B(n60289), .Y(n39696) );
  AND2X1 U40509 ( .A(n60296), .B(n60295), .Y(n39697) );
  OR2X1 U40510 ( .A(n59390), .B(n37378), .Y(n59429) );
  NAND2X1 U40511 ( .A(n42339), .B(n42344), .Y(n39698) );
  AND2X1 U40512 ( .A(n39698), .B(n38813), .Y(n39699) );
  OR2X1 U40513 ( .A(n39700), .B(n69198), .Y(n69259) );
  INVX1 U40514 ( .A(n41013), .Y(n39700) );
  OR2X1 U40515 ( .A(n38555), .B(n71181), .Y(n71183) );
  OR2X1 U40516 ( .A(n42834), .B(n38663), .Y(n39701) );
  OR2X1 U40517 ( .A(n39703), .B(n39702), .Y(n66215) );
  INVX1 U40518 ( .A(n66506), .Y(n39702) );
  AND2X1 U40519 ( .A(n66214), .B(n43626), .Y(n39703) );
  AND2X1 U40520 ( .A(n70588), .B(n70587), .Y(n39704) );
  INVX1 U40521 ( .A(n39704), .Y(n71043) );
  OR2X1 U40522 ( .A(n39911), .B(n39912), .Y(n39705) );
  AND2X1 U40523 ( .A(n60484), .B(n60485), .Y(n39706) );
  AND2X1 U40524 ( .A(n41825), .B(n60360), .Y(n39707) );
  AND2X1 U40525 ( .A(n65978), .B(n65994), .Y(n39708) );
  OR2X1 U40526 ( .A(n40083), .B(n40084), .Y(n39709) );
  OR2X1 U40527 ( .A(n40602), .B(n40603), .Y(n39710) );
  INVX1 U40528 ( .A(n41878), .Y(n39711) );
  AND2X1 U40529 ( .A(n60504), .B(n60503), .Y(n39712) );
  OR2X1 U40530 ( .A(n38992), .B(n38990), .Y(n59755) );
  AND2X1 U40531 ( .A(n60709), .B(n60712), .Y(n39713) );
  NAND2X1 U40532 ( .A(n59146), .B(n59678), .Y(n39714) );
  AND2X1 U40533 ( .A(n66013), .B(n66012), .Y(n39715) );
  AND2X1 U40534 ( .A(n63334), .B(n39719), .Y(n39716) );
  OR2X1 U40535 ( .A(n39716), .B(n39717), .Y(n63600) );
  AND2X1 U40536 ( .A(n39718), .B(n42844), .Y(n39717) );
  INVX1 U40537 ( .A(n63599), .Y(n39718) );
  AND2X1 U40538 ( .A(n63333), .B(n39718), .Y(n39719) );
  OR2X1 U40539 ( .A(n39720), .B(n39721), .Y(n72661) );
  OR2X1 U40540 ( .A(n72660), .B(n72709), .Y(n39720) );
  AND2X1 U40541 ( .A(n38818), .B(n40456), .Y(n39721) );
  OR2X1 U40542 ( .A(n39722), .B(n37374), .Y(n71700) );
  OR2X1 U40543 ( .A(n41047), .B(n40944), .Y(n39722) );
  OR2X1 U40544 ( .A(n61707), .B(n61706), .Y(n61708) );
  AND2X1 U40545 ( .A(n62480), .B(n62481), .Y(n39723) );
  INVX1 U40546 ( .A(n39723), .Y(n62976) );
  AND2X1 U40547 ( .A(n39423), .B(n38981), .Y(n39724) );
  NOR2X1 U40548 ( .A(n39726), .B(n39727), .Y(n39725) );
  AND2X1 U40549 ( .A(n71175), .B(n39301), .Y(n39726) );
  AND2X1 U40550 ( .A(n71177), .B(n39301), .Y(n39727) );
  NOR2X1 U40551 ( .A(n39729), .B(n39730), .Y(n39728) );
  INVX1 U40552 ( .A(n39728), .Y(n71201) );
  OR2X1 U40553 ( .A(n70864), .B(n70863), .Y(n39729) );
  AND2X1 U40554 ( .A(n70866), .B(n70865), .Y(n39730) );
  AND2X1 U40555 ( .A(n63245), .B(n63246), .Y(n62953) );
  AND2X1 U40556 ( .A(n68458), .B(n68459), .Y(n39731) );
  NAND2X1 U40557 ( .A(n36723), .B(n39735), .Y(n39732) );
  AND2X1 U40558 ( .A(n39732), .B(n39733), .Y(n60200) );
  OR2X1 U40559 ( .A(n39734), .B(n59939), .Y(n39733) );
  INVX1 U40560 ( .A(n60197), .Y(n39734) );
  AND2X1 U40561 ( .A(n60197), .B(n59938), .Y(n39735) );
  OR2X1 U40562 ( .A(n39736), .B(n39737), .Y(n63060) );
  AND2X1 U40563 ( .A(n62334), .B(n62333), .Y(n39736) );
  AND2X1 U40564 ( .A(n42112), .B(n62336), .Y(n39737) );
  OR2X1 U40565 ( .A(n39738), .B(n39739), .Y(n66257) );
  AND2X1 U40566 ( .A(n40142), .B(n66535), .Y(n39738) );
  AND2X1 U40567 ( .A(n66228), .B(n66534), .Y(n39739) );
  NOR2X1 U40568 ( .A(n39741), .B(n39742), .Y(n39740) );
  OR2X1 U40569 ( .A(n40437), .B(n65873), .Y(n39741) );
  AND2X1 U40570 ( .A(n65974), .B(n39708), .Y(n39742) );
  OR2X1 U40571 ( .A(n64448), .B(n40151), .Y(n64729) );
  OR2X1 U40572 ( .A(n39743), .B(n39744), .Y(n60617) );
  AND2X1 U40573 ( .A(n60226), .B(n38527), .Y(n39743) );
  AND2X1 U40574 ( .A(n60230), .B(n60229), .Y(n39744) );
  AND2X1 U40575 ( .A(n59752), .B(n59755), .Y(n39745) );
  NAND2X1 U40576 ( .A(n69501), .B(n69626), .Y(n39746) );
  OR2X1 U40577 ( .A(n39747), .B(n39748), .Y(n39842) );
  INVX1 U40578 ( .A(n43673), .Y(n39747) );
  OR2X1 U40579 ( .A(n63117), .B(n37382), .Y(n63672) );
  AND2X1 U40580 ( .A(n63650), .B(n63649), .Y(n39749) );
  NOR2X1 U40581 ( .A(n39751), .B(n39752), .Y(n39750) );
  AND2X1 U40582 ( .A(n60728), .B(n60727), .Y(n39751) );
  AND2X1 U40583 ( .A(n60733), .B(n60732), .Y(n39752) );
  OR2X1 U40584 ( .A(n39753), .B(n39515), .Y(n67318) );
  OR2X1 U40585 ( .A(n41178), .B(n41146), .Y(n39753) );
  NOR2X1 U40586 ( .A(n39755), .B(n39756), .Y(n39754) );
  AND2X1 U40587 ( .A(n59215), .B(n40430), .Y(n39755) );
  AND2X1 U40588 ( .A(n59217), .B(n59216), .Y(n39756) );
  AND2X1 U40589 ( .A(n63130), .B(n39926), .Y(n39757) );
  AND2X1 U40590 ( .A(n63879), .B(n63878), .Y(n39758) );
  INVX1 U40591 ( .A(n39758), .Y(n64044) );
  OR2X1 U40592 ( .A(n39759), .B(n39760), .Y(n66928) );
  INVX1 U40593 ( .A(n67584), .Y(n39759) );
  AND2X1 U40594 ( .A(n66586), .B(n66585), .Y(n39760) );
  AND2X1 U40595 ( .A(n43465), .B(n42708), .Y(n39761) );
  INVX1 U40596 ( .A(n39761), .Y(n59257) );
  NOR2X1 U40597 ( .A(n39763), .B(n39764), .Y(n39762) );
  AND2X1 U40598 ( .A(n38232), .B(n59581), .Y(n39763) );
  AND2X1 U40599 ( .A(n59584), .B(n59583), .Y(n39764) );
  NOR2X1 U40600 ( .A(n39305), .B(n39829), .Y(n39765) );
  AND2X1 U40601 ( .A(n39766), .B(n39767), .Y(n45264) );
  NOR2X1 U40602 ( .A(writeback_exec_idx_w[0]), .B(n40528), .Y(n39767) );
  NOR2X1 U40603 ( .A(n39911), .B(n39912), .Y(n39768) );
  AND2X1 U40604 ( .A(n62862), .B(n62860), .Y(n39769) );
  OR2X1 U40605 ( .A(n36608), .B(n39770), .Y(n40857) );
  INVX1 U40606 ( .A(n40512), .Y(n39770) );
  AND2X1 U40607 ( .A(n63275), .B(n62981), .Y(n39771) );
  OR2X1 U40608 ( .A(n39772), .B(n39773), .Y(n64162) );
  AND2X1 U40609 ( .A(n64161), .B(n64382), .Y(n39772) );
  NOR2X1 U40610 ( .A(n40983), .B(n64382), .Y(n39773) );
  AND2X1 U40611 ( .A(n59550), .B(n59549), .Y(n39774) );
  OR2X1 U40612 ( .A(n39775), .B(n40747), .Y(n70228) );
  NAND2X1 U40613 ( .A(n70155), .B(n70224), .Y(n39775) );
  OR2X1 U40614 ( .A(n39777), .B(n39776), .Y(n65299) );
  INVX1 U40615 ( .A(n65293), .Y(n39776) );
  OR2X1 U40616 ( .A(n41557), .B(n41608), .Y(n39777) );
  AND2X1 U40617 ( .A(n39778), .B(n37319), .Y(n65640) );
  OR2X1 U40618 ( .A(n64959), .B(n65477), .Y(n39778) );
  AND2X1 U40619 ( .A(n67324), .B(n41155), .Y(n39779) );
  AND2X1 U40620 ( .A(n59463), .B(n59503), .Y(n39780) );
  OR2X1 U40621 ( .A(n39781), .B(n39782), .Y(n63902) );
  INVX1 U40622 ( .A(n41994), .Y(n39781) );
  OR2X1 U40623 ( .A(n39783), .B(n39784), .Y(n65876) );
  OR2X1 U40624 ( .A(n39846), .B(n65269), .Y(n39783) );
  AND2X1 U40625 ( .A(n65276), .B(n65275), .Y(n39784) );
  OR2X1 U40626 ( .A(n39785), .B(n39372), .Y(n70238) );
  NOR2X1 U40627 ( .A(n70116), .B(n43584), .Y(n39785) );
  OR2X1 U40628 ( .A(n39786), .B(n39787), .Y(n59982) );
  AND2X1 U40629 ( .A(n60019), .B(n60017), .Y(n39786) );
  AND2X1 U40630 ( .A(n41843), .B(n59818), .Y(n39787) );
  NOR2X1 U40631 ( .A(n39789), .B(n39790), .Y(n39788) );
  INVX1 U40632 ( .A(n71243), .Y(n39789) );
  AND2X1 U40633 ( .A(n71234), .B(n43597), .Y(n39790) );
  OR2X1 U40634 ( .A(n39791), .B(n39792), .Y(n59597) );
  AND2X1 U40635 ( .A(n59566), .B(n59635), .Y(n39791) );
  AND2X1 U40636 ( .A(n41842), .B(n59567), .Y(n39792) );
  AND2X1 U40637 ( .A(n63619), .B(n63608), .Y(n39793) );
  INVX1 U40638 ( .A(n39793), .Y(n63883) );
  AND2X1 U40639 ( .A(n59124), .B(n40391), .Y(n39794) );
  AND2X1 U40640 ( .A(n59476), .B(n59475), .Y(n39795) );
  OR2X1 U40641 ( .A(n39796), .B(n43519), .Y(n62940) );
  OR2X1 U40642 ( .A(n43460), .B(n62466), .Y(n39796) );
  XNOR2X1 U40643 ( .A(n66883), .B(n39469), .Y(n39797) );
  XNOR2X1 U40644 ( .A(n66883), .B(n39469), .Y(n39798) );
  INVX1 U40645 ( .A(n39802), .Y(n39799) );
  INVX1 U40646 ( .A(n39806), .Y(n39800) );
  INVX1 U40647 ( .A(n48146), .Y(n39801) );
  INVX1 U40648 ( .A(n39582), .Y(n39802) );
  INVX1 U40649 ( .A(n39583), .Y(n39803) );
  INVX1 U40650 ( .A(n39583), .Y(n39804) );
  INVX1 U40651 ( .A(n39582), .Y(n39805) );
  INVX1 U40652 ( .A(n39582), .Y(n39806) );
  INVX1 U40653 ( .A(n39583), .Y(n39807) );
  INVX1 U40654 ( .A(n39582), .Y(n39808) );
  INVX1 U40655 ( .A(n38366), .Y(n39810) );
  AND2X1 U40656 ( .A(n70448), .B(n70447), .Y(n39811) );
  OR2X1 U40657 ( .A(n59284), .B(n59285), .Y(n59294) );
  OR2X1 U40658 ( .A(n40547), .B(n40548), .Y(n39812) );
  INVX1 U40659 ( .A(n39812), .Y(n40546) );
  NOR2X1 U40660 ( .A(n39814), .B(n39815), .Y(n39813) );
  AND2X1 U40661 ( .A(n61405), .B(n61406), .Y(n39814) );
  AND2X1 U40662 ( .A(n41936), .B(n61407), .Y(n39815) );
  OR2X1 U40663 ( .A(n40644), .B(n40645), .Y(n39816) );
  NAND2X1 U40664 ( .A(n64729), .B(n39820), .Y(n39817) );
  NAND2X1 U40665 ( .A(n39817), .B(n39818), .Y(n40974) );
  OR2X1 U40666 ( .A(n39819), .B(n64732), .Y(n39818) );
  INVX1 U40667 ( .A(n65026), .Y(n39819) );
  AND2X1 U40668 ( .A(n64730), .B(n65026), .Y(n39820) );
  AND2X1 U40669 ( .A(n61414), .B(n41956), .Y(n39821) );
  OR2X1 U40670 ( .A(n39821), .B(n39822), .Y(n61416) );
  OR2X1 U40671 ( .A(n39823), .B(n40012), .Y(n39822) );
  INVX1 U40672 ( .A(n61455), .Y(n39823) );
  AND2X1 U40673 ( .A(n59726), .B(n59729), .Y(n39824) );
  OR2X1 U40674 ( .A(n39825), .B(n48105), .Y(n62907) );
  INVX1 U40675 ( .A(n42377), .Y(n39825) );
  AND2X1 U40676 ( .A(n65100), .B(n65101), .Y(n39826) );
  NOR2X1 U40677 ( .A(n39828), .B(n39829), .Y(n39827) );
  OR2X1 U40678 ( .A(n62513), .B(n62512), .Y(n39828) );
  AND2X1 U40679 ( .A(n62516), .B(n62515), .Y(n39829) );
  OR2X1 U40680 ( .A(n61710), .B(n61709), .Y(n61711) );
  NOR2X1 U40681 ( .A(n39831), .B(n39832), .Y(n39830) );
  AND2X1 U40682 ( .A(n61614), .B(n61551), .Y(n39831) );
  AND2X1 U40683 ( .A(n41952), .B(n61553), .Y(n39832) );
  OR2X1 U40684 ( .A(n39833), .B(n39012), .Y(n70480) );
  AND2X1 U40685 ( .A(n41054), .B(n69573), .Y(n39833) );
  OR2X1 U40686 ( .A(n39834), .B(n39835), .Y(n62363) );
  INVX1 U40687 ( .A(n62354), .Y(n39834) );
  AND2X1 U40688 ( .A(n61099), .B(n62357), .Y(n39835) );
  AND2X1 U40689 ( .A(n64381), .B(n64380), .Y(n39836) );
  INVX1 U40690 ( .A(n39836), .Y(n64387) );
  OR2X1 U40691 ( .A(n39837), .B(n36772), .Y(n62453) );
  OR2X1 U40692 ( .A(n62896), .B(n62897), .Y(n39837) );
  OR2X1 U40693 ( .A(n65602), .B(n39838), .Y(n65606) );
  INVX1 U40694 ( .A(n43531), .Y(n39838) );
  OR2X1 U40695 ( .A(n39839), .B(n39840), .Y(n66504) );
  OR2X1 U40696 ( .A(n65983), .B(n65982), .Y(n39839) );
  NAND2X1 U40697 ( .A(n68823), .B(n68876), .Y(n39841) );
  INVX1 U40698 ( .A(n39842), .Y(n70457) );
  AND2X1 U40699 ( .A(n70510), .B(n70509), .Y(n39843) );
  INVX1 U40700 ( .A(n36706), .Y(n39844) );
  AND2X1 U40701 ( .A(n66485), .B(n66484), .Y(n39845) );
  OR2X1 U40702 ( .A(n59654), .B(n59655), .Y(n59656) );
  AND2X1 U40703 ( .A(n39147), .B(n65272), .Y(n39846) );
  INVX1 U40704 ( .A(n39846), .Y(n65268) );
  OR2X1 U40705 ( .A(n40031), .B(n40032), .Y(n39847) );
  AND2X1 U40706 ( .A(n64633), .B(n64632), .Y(n39848) );
  OR2X1 U40707 ( .A(n39849), .B(n39850), .Y(n62439) );
  AND2X1 U40708 ( .A(n61170), .B(n61169), .Y(n39849) );
  AND2X1 U40709 ( .A(n61173), .B(n61172), .Y(n39850) );
  INVX1 U40710 ( .A(n39991), .Y(n39851) );
  INVX1 U40711 ( .A(n67653), .Y(n39852) );
  NAND2X1 U40712 ( .A(n42801), .B(n62453), .Y(n39853) );
  NOR2X1 U40713 ( .A(n64175), .B(n64176), .Y(n39854) );
  INVX1 U40714 ( .A(n39854), .Y(n64456) );
  AND2X1 U40715 ( .A(n43631), .B(n36735), .Y(n39855) );
  INVX1 U40716 ( .A(n39855), .Y(n69516) );
  OR2X1 U40717 ( .A(n39856), .B(n39857), .Y(n67016) );
  OR2X1 U40718 ( .A(n66828), .B(n66827), .Y(n39856) );
  AND2X1 U40719 ( .A(n66831), .B(n66830), .Y(n39857) );
  AND2X1 U40720 ( .A(n38203), .B(n70152), .Y(n39858) );
  NOR2X1 U40721 ( .A(n39860), .B(n39861), .Y(n39859) );
  OR2X1 U40722 ( .A(n61031), .B(n61030), .Y(n39860) );
  AND2X1 U40723 ( .A(n61033), .B(n61032), .Y(n39861) );
  AND2X1 U40724 ( .A(n70248), .B(n43586), .Y(n39862) );
  INVX1 U40725 ( .A(n39862), .Y(n70561) );
  NOR2X1 U40726 ( .A(n39864), .B(n39865), .Y(n39863) );
  INVX1 U40727 ( .A(n38957), .Y(n61034) );
  AND2X1 U40728 ( .A(n36787), .B(n60584), .Y(n39864) );
  AND2X1 U40729 ( .A(n41499), .B(n60585), .Y(n39865) );
  NOR2X1 U40730 ( .A(n39867), .B(n36762), .Y(n39866) );
  INVX1 U40731 ( .A(n39866), .Y(n71414) );
  AND2X1 U40732 ( .A(n71156), .B(n71155), .Y(n39867) );
  NAND2X1 U40733 ( .A(n39650), .B(n39604), .Y(n39868) );
  NOR2X1 U40734 ( .A(n70121), .B(n39963), .Y(n39869) );
  AND2X1 U40735 ( .A(n67960), .B(n67959), .Y(n39870) );
  OR2X1 U40736 ( .A(n39871), .B(n39872), .Y(n67841) );
  OR2X1 U40737 ( .A(n67832), .B(n41403), .Y(n39871) );
  OR2X1 U40738 ( .A(n67827), .B(n37356), .Y(n39872) );
  NOR2X1 U40739 ( .A(n39874), .B(n39875), .Y(n39873) );
  AND2X1 U40740 ( .A(n60883), .B(n60882), .Y(n39874) );
  AND2X1 U40741 ( .A(n42015), .B(n60885), .Y(n39875) );
  OR2X1 U40742 ( .A(n59535), .B(n59537), .Y(n59572) );
  OR2X1 U40743 ( .A(n39876), .B(n39877), .Y(n59445) );
  AND2X1 U40744 ( .A(n59386), .B(n59388), .Y(n39876) );
  AND2X1 U40745 ( .A(n41483), .B(n59380), .Y(n39877) );
  OR2X1 U40746 ( .A(n39878), .B(n39879), .Y(n63917) );
  OR2X1 U40747 ( .A(n63454), .B(n41265), .Y(n39878) );
  AND2X1 U40748 ( .A(n63460), .B(n63918), .Y(n39879) );
  OR2X1 U40749 ( .A(n60772), .B(n39880), .Y(n60520) );
  AND2X1 U40750 ( .A(n60773), .B(n38244), .Y(n39880) );
  AND2X1 U40751 ( .A(n63134), .B(n63135), .Y(n39881) );
  NAND2X1 U40752 ( .A(n42668), .B(n42786), .Y(n39882) );
  NAND2X1 U40753 ( .A(n42667), .B(n42786), .Y(n39883) );
  OR2X1 U40754 ( .A(n39884), .B(n39885), .Y(n66198) );
  AND2X1 U40755 ( .A(n65843), .B(n66192), .Y(n39884) );
  AND2X1 U40756 ( .A(n65851), .B(n65850), .Y(n39885) );
  NOR2X1 U40757 ( .A(n41767), .B(n41768), .Y(n39886) );
  AND2X1 U40758 ( .A(n43677), .B(n70504), .Y(n39887) );
  INVX1 U40759 ( .A(n39887), .Y(n70501) );
  AND2X1 U40760 ( .A(n67945), .B(n67946), .Y(n39888) );
  OR2X1 U40761 ( .A(n39889), .B(n39890), .Y(n71153) );
  OR2X1 U40762 ( .A(n41307), .B(n71110), .Y(n39889) );
  OR2X1 U40763 ( .A(n41301), .B(n71113), .Y(n39890) );
  AND2X1 U40764 ( .A(n65458), .B(n65457), .Y(n39891) );
  NOR2X1 U40765 ( .A(n39893), .B(n39894), .Y(n39892) );
  AND2X1 U40766 ( .A(n39710), .B(n59867), .Y(n39893) );
  AND2X1 U40767 ( .A(n59871), .B(n59870), .Y(n39894) );
  AND2X1 U40768 ( .A(n65910), .B(n66514), .Y(n39895) );
  OR2X1 U40769 ( .A(n39896), .B(n39897), .Y(n66506) );
  AND2X1 U40770 ( .A(n43620), .B(n65611), .Y(n39896) );
  AND2X1 U40771 ( .A(n65613), .B(n65614), .Y(n39897) );
  AND2X1 U40772 ( .A(n59343), .B(n59342), .Y(n39898) );
  AND2X1 U40773 ( .A(n61204), .B(n39061), .Y(n39899) );
  NOR2X1 U40774 ( .A(n39901), .B(n39902), .Y(n39900) );
  AND2X1 U40775 ( .A(n59930), .B(n40242), .Y(n39901) );
  AND2X1 U40776 ( .A(n59934), .B(n59933), .Y(n39902) );
  OR2X1 U40777 ( .A(n65521), .B(n65520), .Y(n39903) );
  OR2X1 U40778 ( .A(n60263), .B(n37377), .Y(n60665) );
  OR2X1 U40779 ( .A(n39904), .B(n39905), .Y(n66176) );
  AND2X1 U40780 ( .A(n65835), .B(n65823), .Y(n39904) );
  AND2X1 U40781 ( .A(n65826), .B(n65825), .Y(n39905) );
  OR2X1 U40782 ( .A(n46394), .B(n46231), .Y(n46903) );
  AND2X1 U40783 ( .A(n41054), .B(n69573), .Y(n39906) );
  INVX1 U40784 ( .A(n39906), .Y(n70174) );
  OR2X1 U40785 ( .A(n39907), .B(n39908), .Y(n60584) );
  OR2X1 U40786 ( .A(n60220), .B(n60219), .Y(n39907) );
  AND2X1 U40787 ( .A(n60222), .B(n60221), .Y(n39908) );
  AND2X1 U40788 ( .A(n39714), .B(n59231), .Y(n39909) );
  NOR2X1 U40789 ( .A(n39911), .B(n39912), .Y(n39910) );
  INVX1 U40790 ( .A(n63308), .Y(n39911) );
  AND2X1 U40791 ( .A(n63307), .B(n62882), .Y(n39912) );
  AND2X1 U40792 ( .A(n64022), .B(n64023), .Y(n39913) );
  NOR2X1 U40793 ( .A(n39915), .B(n39916), .Y(n39914) );
  AND2X1 U40794 ( .A(n60207), .B(n40435), .Y(n39915) );
  AND2X1 U40795 ( .A(n60211), .B(n60210), .Y(n39916) );
  OR2X1 U40796 ( .A(n39917), .B(n39918), .Y(n66205) );
  OR2X1 U40797 ( .A(n65654), .B(n65653), .Y(n39917) );
  AND2X1 U40798 ( .A(n65662), .B(n65661), .Y(n39918) );
  AND2X1 U40799 ( .A(n69515), .B(n69516), .Y(n39919) );
  OR2X1 U40800 ( .A(n39920), .B(n39921), .Y(n63132) );
  OR2X1 U40801 ( .A(n62845), .B(n62844), .Y(n39920) );
  AND2X1 U40802 ( .A(n62848), .B(n62847), .Y(n39921) );
  OR2X1 U40803 ( .A(n43697), .B(n72699), .Y(n72697) );
  AND2X1 U40804 ( .A(n71137), .B(n43696), .Y(n39922) );
  AND2X1 U40805 ( .A(n66079), .B(n39343), .Y(n39923) );
  NOR2X1 U40806 ( .A(n39995), .B(n39996), .Y(n39924) );
  OR2X1 U40807 ( .A(n43585), .B(n70248), .Y(n70562) );
  AND2X1 U40808 ( .A(n70788), .B(n36564), .Y(n39925) );
  INVX1 U40809 ( .A(n39925), .Y(n70814) );
  NAND2X1 U40810 ( .A(n62841), .B(n62840), .Y(n39926) );
  OR2X1 U40811 ( .A(n70136), .B(n39927), .Y(n70128) );
  INVX1 U40812 ( .A(n43538), .Y(n39927) );
  OR2X1 U40813 ( .A(n66224), .B(n39928), .Y(n66523) );
  INVX1 U40814 ( .A(n43552), .Y(n39928) );
  AND2X1 U40815 ( .A(n66483), .B(n66479), .Y(n39929) );
  AND2X1 U40816 ( .A(n68761), .B(n68760), .Y(n39930) );
  NAND2X1 U40817 ( .A(n38193), .B(n65875), .Y(n39931) );
  OR2X1 U40818 ( .A(n39932), .B(n39933), .Y(n64328) );
  AND2X1 U40819 ( .A(n63896), .B(n64010), .Y(n39932) );
  NOR2X1 U40820 ( .A(n41603), .B(n41604), .Y(n39933) );
  INVX1 U40821 ( .A(n64459), .Y(n39934) );
  AND2X1 U40822 ( .A(n64458), .B(n64457), .Y(n39935) );
  OR2X1 U40823 ( .A(n38484), .B(n65987), .Y(n39936) );
  INVX1 U40824 ( .A(n42226), .Y(n39937) );
  INVX1 U40825 ( .A(n38459), .Y(n39938) );
  INVX1 U40826 ( .A(n38459), .Y(n39939) );
  INVX1 U40827 ( .A(n38459), .Y(n39940) );
  INVX1 U40828 ( .A(n38459), .Y(n39941) );
  INVX1 U40829 ( .A(n38459), .Y(n39942) );
  INVX1 U40830 ( .A(n38459), .Y(n39943) );
  INVX1 U40831 ( .A(n63551), .Y(n39944) );
  INVX1 U40832 ( .A(n63551), .Y(n39945) );
  INVX1 U40833 ( .A(n63551), .Y(n39946) );
  AND2X1 U40834 ( .A(n41440), .B(n37416), .Y(n67679) );
  INVX1 U40835 ( .A(n39259), .Y(n39947) );
  AND2X1 U40836 ( .A(n66865), .B(n66011), .Y(n39948) );
  OR2X1 U40837 ( .A(n39949), .B(n39950), .Y(n69601) );
  OR2X1 U40838 ( .A(n69521), .B(n69520), .Y(n39949) );
  AND2X1 U40839 ( .A(n69525), .B(n69524), .Y(n39950) );
  AND2X1 U40840 ( .A(n72721), .B(n39951), .Y(n72718) );
  AND2X1 U40841 ( .A(n72717), .B(n72719), .Y(n39951) );
  AND2X1 U40842 ( .A(n43697), .B(n71422), .Y(n71421) );
  NAND2X1 U40843 ( .A(n43619), .B(n67861), .Y(n39952) );
  OR2X1 U40844 ( .A(n39953), .B(n39954), .Y(n69840) );
  AND2X1 U40845 ( .A(n69295), .B(n43586), .Y(n39953) );
  AND2X1 U40846 ( .A(n38617), .B(n69298), .Y(n39954) );
  NOR2X1 U40847 ( .A(n39956), .B(n39957), .Y(n39955) );
  AND2X1 U40848 ( .A(n59873), .B(n59872), .Y(n39956) );
  AND2X1 U40849 ( .A(n59877), .B(n59876), .Y(n39957) );
  OR2X1 U40850 ( .A(n39958), .B(n70240), .Y(n70901) );
  INVX1 U40851 ( .A(n43577), .Y(n39958) );
  INVX1 U40852 ( .A(n60942), .Y(n39959) );
  INVX1 U40853 ( .A(n43519), .Y(n39960) );
  INVX1 U40854 ( .A(n43519), .Y(n39961) );
  NOR2X1 U40855 ( .A(n70121), .B(n39963), .Y(n39962) );
  INVX1 U40856 ( .A(n39869), .Y(n70566) );
  AND2X1 U40857 ( .A(n70240), .B(n43573), .Y(n39963) );
  AND2X1 U40858 ( .A(n60248), .B(n39966), .Y(n39964) );
  OR2X1 U40859 ( .A(n39964), .B(n39965), .Y(n60596) );
  AND2X1 U40860 ( .A(n36788), .B(n40615), .Y(n39965) );
  AND2X1 U40861 ( .A(n60249), .B(n36788), .Y(n39966) );
  AND2X1 U40862 ( .A(n64668), .B(n64667), .Y(n39967) );
  INVX1 U40863 ( .A(n39967), .Y(n65522) );
  OR2X1 U40864 ( .A(n39753), .B(n39515), .Y(n67814) );
  AND2X1 U40865 ( .A(n66349), .B(n66348), .Y(n39968) );
  OR2X1 U40866 ( .A(n39970), .B(n39969), .Y(n68063) );
  INVX1 U40867 ( .A(n68062), .Y(n39969) );
  OR2X1 U40868 ( .A(n41187), .B(n41441), .Y(n39970) );
  OR2X1 U40869 ( .A(n40135), .B(n40136), .Y(n39972) );
  AND2X1 U40870 ( .A(n36428), .B(n68232), .Y(n39973) );
  OR2X1 U40871 ( .A(n39974), .B(n39975), .Y(n67556) );
  OR2X1 U40872 ( .A(n67190), .B(n67189), .Y(n39974) );
  AND2X1 U40873 ( .A(n43576), .B(n67191), .Y(n39975) );
  AND2X1 U40874 ( .A(n68812), .B(n68811), .Y(n39976) );
  OR2X1 U40875 ( .A(n39977), .B(n39978), .Y(n64687) );
  OR2X1 U40876 ( .A(n41552), .B(n64684), .Y(n39977) );
  AND2X1 U40877 ( .A(n64686), .B(n64685), .Y(n39978) );
  AND2X1 U40878 ( .A(n67358), .B(n67139), .Y(n39979) );
  INVX1 U40879 ( .A(n39979), .Y(n67352) );
  NOR2X1 U40880 ( .A(n43659), .B(n65965), .Y(n39980) );
  INVX1 U40881 ( .A(n39980), .Y(n66259) );
  NAND2X1 U40882 ( .A(n69840), .B(n39984), .Y(n39981) );
  OR2X1 U40883 ( .A(n39983), .B(n69839), .Y(n39982) );
  INVX1 U40884 ( .A(n69847), .Y(n39983) );
  AND2X1 U40885 ( .A(n69299), .B(n69847), .Y(n39984) );
  NOR2X1 U40886 ( .A(n63113), .B(n39987), .Y(n39986) );
  INVX1 U40887 ( .A(n39986), .Y(n63443) );
  AND2X1 U40888 ( .A(n63445), .B(n63444), .Y(n39987) );
  AND2X1 U40889 ( .A(n43471), .B(n72811), .Y(n40619) );
  NOR2X1 U40890 ( .A(n40079), .B(n37358), .Y(n39988) );
  NAND2X1 U40891 ( .A(n66521), .B(n39992), .Y(n39989) );
  AND2X1 U40892 ( .A(n39989), .B(n39990), .Y(n66890) );
  OR2X1 U40893 ( .A(n39991), .B(n66523), .Y(n39990) );
  INVX1 U40894 ( .A(n66525), .Y(n39991) );
  AND2X1 U40895 ( .A(n66522), .B(n66525), .Y(n39992) );
  NAND2X1 U40896 ( .A(n61012), .B(n61013), .Y(n39993) );
  OR2X1 U40897 ( .A(n43639), .B(n65245), .Y(n65900) );
  NOR2X1 U40898 ( .A(n39995), .B(n39996), .Y(n39994) );
  INVX1 U40899 ( .A(n39924), .Y(n66951) );
  INVX1 U40900 ( .A(n66977), .Y(n39995) );
  AND2X1 U40901 ( .A(n66034), .B(n66033), .Y(n39996) );
  OR2X1 U40902 ( .A(n39997), .B(n39998), .Y(n59626) );
  AND2X1 U40903 ( .A(n59601), .B(n59556), .Y(n39997) );
  AND2X1 U40904 ( .A(n41797), .B(n59557), .Y(n39998) );
  NOR2X1 U40905 ( .A(n40000), .B(n40001), .Y(n39999) );
  INVX1 U40906 ( .A(n39999), .Y(n60877) );
  AND2X1 U40907 ( .A(n60875), .B(n38612), .Y(n40000) );
  AND2X1 U40908 ( .A(n42007), .B(n60876), .Y(n40001) );
  NOR2X1 U40909 ( .A(n40003), .B(n40004), .Y(n40002) );
  INVX1 U40910 ( .A(n39646), .Y(n69176) );
  AND2X1 U40911 ( .A(n68001), .B(n39958), .Y(n40003) );
  AND2X1 U40912 ( .A(n67998), .B(n39958), .Y(n40004) );
  OR2X1 U40913 ( .A(n61722), .B(n61721), .Y(n61723) );
  AND2X1 U40914 ( .A(n65763), .B(n65762), .Y(n40005) );
  OR2X1 U40915 ( .A(n67659), .B(n40006), .Y(n67558) );
  AND2X1 U40916 ( .A(n43580), .B(n39852), .Y(n40006) );
  OR2X1 U40917 ( .A(n40007), .B(n40008), .Y(n63048) );
  INVX1 U40918 ( .A(n42052), .Y(n40007) );
  AND2X1 U40919 ( .A(n39666), .B(n62559), .Y(n40008) );
  NOR2X1 U40920 ( .A(n38240), .B(n39993), .Y(n40009) );
  OR2X1 U40921 ( .A(n61148), .B(n40010), .Y(n61149) );
  INVX1 U40922 ( .A(n60971), .Y(n40010) );
  NOR2X1 U40923 ( .A(n40012), .B(n40013), .Y(n40011) );
  INVX1 U40924 ( .A(n40011), .Y(n61415) );
  AND2X1 U40925 ( .A(n61412), .B(n61413), .Y(n40012) );
  AND2X1 U40926 ( .A(n41956), .B(n61414), .Y(n40013) );
  AND2X1 U40927 ( .A(n62430), .B(n62428), .Y(n40014) );
  NOR2X1 U40928 ( .A(n39723), .B(n62483), .Y(n40015) );
  OR2X1 U40929 ( .A(n40016), .B(n40017), .Y(n63432) );
  INVX1 U40930 ( .A(n42073), .Y(n40016) );
  AND2X1 U40931 ( .A(n40195), .B(n63111), .Y(n40017) );
  AND2X1 U40932 ( .A(n44963), .B(n42725), .Y(n40018) );
  AND2X1 U40933 ( .A(n40835), .B(n40836), .Y(n40019) );
  NOR2X1 U40934 ( .A(n40021), .B(n40022), .Y(n40020) );
  OR2X1 U40935 ( .A(n40770), .B(n41197), .Y(n40021) );
  AND2X1 U40936 ( .A(n69911), .B(n69572), .Y(n40022) );
  AND2X1 U40937 ( .A(n62889), .B(n63292), .Y(n62888) );
  AND2X1 U40938 ( .A(n43019), .B(n40018), .Y(n40023) );
  INVX1 U40939 ( .A(n40023), .Y(n47685) );
  AND2X1 U40940 ( .A(n62428), .B(n62429), .Y(n40024) );
  INVX1 U40941 ( .A(n40024), .Y(n62982) );
  AND2X1 U40942 ( .A(n64520), .B(n64521), .Y(n40025) );
  INVX1 U40943 ( .A(n48380), .Y(n40026) );
  AND2X1 U40944 ( .A(n39297), .B(n67675), .Y(n40027) );
  AND2X1 U40945 ( .A(n62366), .B(n62365), .Y(n40028) );
  OR2X1 U40946 ( .A(n40029), .B(n69872), .Y(n69585) );
  AND2X1 U40947 ( .A(n43642), .B(n69257), .Y(n40029) );
  NOR2X1 U40948 ( .A(n40031), .B(n40032), .Y(n40030) );
  AND2X1 U40949 ( .A(n61609), .B(n61556), .Y(n40031) );
  AND2X1 U40950 ( .A(n41971), .B(n61558), .Y(n40032) );
  OR2X1 U40951 ( .A(n40033), .B(n40034), .Y(u_muldiv_result_r[31]) );
  NOR2X1 U40952 ( .A(n40541), .B(n40542), .Y(n40034) );
  NOR2X1 U40953 ( .A(n40870), .B(n58469), .Y(n40035) );
  INVX1 U40954 ( .A(n40035), .Y(n57605) );
  OR2X1 U40955 ( .A(n40036), .B(n40037), .Y(n59648) );
  AND2X1 U40956 ( .A(n59642), .B(n59641), .Y(n40036) );
  AND2X1 U40957 ( .A(n59644), .B(n59643), .Y(n40037) );
  OR2X1 U40958 ( .A(n40109), .B(n40110), .Y(n40038) );
  OR2X1 U40959 ( .A(n40039), .B(n40040), .Y(n60444) );
  AND2X1 U40960 ( .A(n60512), .B(n60511), .Y(n40039) );
  AND2X1 U40961 ( .A(n60387), .B(n60386), .Y(n40040) );
  NAND2X1 U40962 ( .A(n42149), .B(n47422), .Y(n40041) );
  NAND2X1 U40963 ( .A(n42149), .B(n47422), .Y(n40042) );
  OR2X1 U40964 ( .A(n40044), .B(n40043), .Y(n66569) );
  AND2X1 U40965 ( .A(n66566), .B(n43699), .Y(n40044) );
  OR2X1 U40966 ( .A(n65037), .B(n37397), .Y(n65429) );
  OR2X1 U40967 ( .A(n40045), .B(n40046), .Y(n62397) );
  AND2X1 U40968 ( .A(n61120), .B(n61119), .Y(n40045) );
  AND2X1 U40969 ( .A(n61125), .B(n61124), .Y(n40046) );
  NOR2X1 U40970 ( .A(n40048), .B(n40049), .Y(n40047) );
  INVX1 U40971 ( .A(n40047), .Y(n59635) );
  AND2X1 U40972 ( .A(n38796), .B(n59600), .Y(n40048) );
  AND2X1 U40973 ( .A(n41827), .B(n59565), .Y(n40049) );
  OR2X1 U40974 ( .A(n43698), .B(n66918), .Y(n67607) );
  OR2X1 U40975 ( .A(n40050), .B(n40051), .Y(n61192) );
  OR2X1 U40976 ( .A(n60947), .B(n60946), .Y(n40050) );
  OR2X1 U40977 ( .A(n60949), .B(n60948), .Y(n40051) );
  AND2X1 U40978 ( .A(n64687), .B(n38377), .Y(n40052) );
  NOR2X1 U40979 ( .A(n40054), .B(n40055), .Y(n40053) );
  INVX1 U40980 ( .A(n40053), .Y(n60141) );
  AND2X1 U40981 ( .A(n60102), .B(n60013), .Y(n40054) );
  AND2X1 U40982 ( .A(n41835), .B(n60014), .Y(n40055) );
  OR2X1 U40983 ( .A(n40056), .B(n40057), .Y(n68200) );
  INVX1 U40984 ( .A(n67652), .Y(n40056) );
  AND2X1 U40985 ( .A(n67651), .B(n68263), .Y(n40057) );
  OR2X1 U40986 ( .A(n40058), .B(n40059), .Y(n66937) );
  AND2X1 U40987 ( .A(n43565), .B(n66616), .Y(n40058) );
  AND2X1 U40988 ( .A(n66618), .B(n66617), .Y(n40059) );
  OR2X1 U40989 ( .A(n60587), .B(n60661), .Y(n61019) );
  OR2X1 U40990 ( .A(n40060), .B(n40061), .Y(n67640) );
  OR2X1 U40991 ( .A(n37385), .B(n67207), .Y(n40060) );
  AND2X1 U40992 ( .A(n67215), .B(n67214), .Y(n40061) );
  OR2X1 U40993 ( .A(n40062), .B(n40063), .Y(n61324) );
  AND2X1 U40994 ( .A(n60840), .B(n36417), .Y(n40062) );
  AND2X1 U40995 ( .A(n41902), .B(n60841), .Y(n40063) );
  AND2X1 U40996 ( .A(n63165), .B(n63164), .Y(n40064) );
  OR2X1 U40997 ( .A(n40065), .B(n40066), .Y(n60440) );
  AND2X1 U40998 ( .A(n60161), .B(n60162), .Y(n40065) );
  AND2X1 U40999 ( .A(n41910), .B(n60163), .Y(n40066) );
  NOR2X1 U41000 ( .A(n40068), .B(n40069), .Y(n40067) );
  AND2X1 U41001 ( .A(n60779), .B(n60506), .Y(n40068) );
  AND2X1 U41002 ( .A(n41889), .B(n60508), .Y(n40069) );
  OR2X1 U41003 ( .A(n40070), .B(n40071), .Y(n64356) );
  OR2X1 U41004 ( .A(n64049), .B(n64048), .Y(n40070) );
  AND2X1 U41005 ( .A(n64050), .B(n39431), .Y(n40071) );
  AND2X1 U41006 ( .A(n42044), .B(n64666), .Y(n40072) );
  NOR2X1 U41007 ( .A(n40074), .B(n40075), .Y(n40073) );
  AND2X1 U41008 ( .A(n61428), .B(n61429), .Y(n40074) );
  AND2X1 U41009 ( .A(n42031), .B(n61430), .Y(n40075) );
  INVX1 U41010 ( .A(n42855), .Y(n40076) );
  AND2X1 U41011 ( .A(n65866), .B(n65865), .Y(n40077) );
  NOR2X1 U41012 ( .A(n40079), .B(n37358), .Y(n40078) );
  OR2X1 U41013 ( .A(n41258), .B(n41290), .Y(n40079) );
  OR2X1 U41014 ( .A(n40080), .B(n40081), .Y(n62494) );
  AND2X1 U41015 ( .A(n61130), .B(n61129), .Y(n40080) );
  AND2X1 U41016 ( .A(n61133), .B(n61134), .Y(n40081) );
  NOR2X1 U41017 ( .A(n40083), .B(n40084), .Y(n40082) );
  AND2X1 U41018 ( .A(n61220), .B(n61219), .Y(n40083) );
  AND2X1 U41019 ( .A(n61224), .B(n61223), .Y(n40084) );
  AND2X1 U41020 ( .A(n67283), .B(n41066), .Y(n40085) );
  AND2X1 U41021 ( .A(n61168), .B(n61167), .Y(n40086) );
  AND2X1 U41022 ( .A(n40772), .B(n40771), .Y(n40087) );
  AND2X1 U41023 ( .A(n70534), .B(n70535), .Y(n40088) );
  INVX1 U41024 ( .A(n67249), .Y(n40089) );
  NOR2X1 U41025 ( .A(n40089), .B(n67250), .Y(n40090) );
  OR2X1 U41026 ( .A(n40091), .B(n40092), .Y(n62344) );
  AND2X1 U41027 ( .A(n61094), .B(n39678), .Y(n40091) );
  AND2X1 U41028 ( .A(n42025), .B(n61096), .Y(n40092) );
  OR2X1 U41029 ( .A(n43657), .B(n70475), .Y(n70513) );
  XNOR2X1 U41030 ( .A(n68195), .B(n68796), .Y(n40093) );
  AND2X1 U41031 ( .A(n62437), .B(n62436), .Y(n40094) );
  OR2X1 U41032 ( .A(n40095), .B(n40096), .Y(n70829) );
  OR2X1 U41033 ( .A(n39331), .B(n70474), .Y(n40095) );
  AND2X1 U41034 ( .A(n70475), .B(n43658), .Y(n40096) );
  NAND2X1 U41035 ( .A(n40386), .B(n40100), .Y(n40097) );
  AND2X1 U41036 ( .A(n40097), .B(n40098), .Y(n64541) );
  OR2X1 U41037 ( .A(n40099), .B(n63976), .Y(n40098) );
  INVX1 U41038 ( .A(n63977), .Y(n40099) );
  AND2X1 U41039 ( .A(n40387), .B(n63977), .Y(n40100) );
  OR2X1 U41040 ( .A(n40101), .B(n40102), .Y(n61732) );
  INVX1 U41041 ( .A(n42030), .Y(n40101) );
  OR2X1 U41042 ( .A(n40103), .B(n40104), .Y(n68078) );
  OR2X1 U41043 ( .A(n67695), .B(n67694), .Y(n40103) );
  AND2X1 U41044 ( .A(n67697), .B(n67696), .Y(n40104) );
  NOR2X1 U41045 ( .A(n43688), .B(n64582), .Y(n40105) );
  OR2X1 U41046 ( .A(n40494), .B(n40495), .Y(n40106) );
  NAND2X1 U41047 ( .A(n40523), .B(n42772), .Y(n40107) );
  NOR2X1 U41048 ( .A(n40109), .B(n40110), .Y(n40108) );
  AND2X1 U41049 ( .A(n61605), .B(n61563), .Y(n40109) );
  AND2X1 U41050 ( .A(n41990), .B(n61564), .Y(n40110) );
  NOR2X1 U41051 ( .A(n40112), .B(n40113), .Y(n40111) );
  AND2X1 U41052 ( .A(n38280), .B(n59863), .Y(n40112) );
  NOR2X1 U41053 ( .A(n59864), .B(n40646), .Y(n40113) );
  NAND2X1 U41054 ( .A(n65237), .B(n40117), .Y(n40114) );
  AND2X1 U41055 ( .A(n40114), .B(n40115), .Y(n65961) );
  OR2X1 U41056 ( .A(n40116), .B(n65604), .Y(n40115) );
  INVX1 U41057 ( .A(n65606), .Y(n40116) );
  AND2X1 U41058 ( .A(n65238), .B(n65606), .Y(n40117) );
  NAND2X1 U41059 ( .A(n66569), .B(n40120), .Y(n40118) );
  AND2X1 U41060 ( .A(n40118), .B(n40119), .Y(n67609) );
  OR2X1 U41061 ( .A(n36410), .B(n66920), .Y(n40119) );
  AND2X1 U41062 ( .A(n67607), .B(n66568), .Y(n40120) );
  NAND2X1 U41063 ( .A(n59675), .B(n59674), .Y(n40121) );
  AND2X1 U41064 ( .A(n66075), .B(n66076), .Y(n40122) );
  AND2X1 U41065 ( .A(n70211), .B(n70210), .Y(n40123) );
  OR2X1 U41066 ( .A(n40124), .B(n40125), .Y(n67914) );
  AND2X1 U41067 ( .A(n43706), .B(n67244), .Y(n40124) );
  AND2X1 U41068 ( .A(n37907), .B(n67245), .Y(n40125) );
  OR2X1 U41069 ( .A(n40126), .B(n40127), .Y(n71179) );
  OR2X1 U41070 ( .A(n40088), .B(n37402), .Y(n40126) );
  AND2X1 U41071 ( .A(n43631), .B(n70854), .Y(n40127) );
  NOR2X1 U41072 ( .A(n40129), .B(n67005), .Y(n40128) );
  INVX1 U41073 ( .A(n40128), .Y(n67506) );
  OR2X1 U41074 ( .A(n38139), .B(n67167), .Y(n40129) );
  AND2X1 U41075 ( .A(n67708), .B(n40130), .Y(n67711) );
  AND2X1 U41076 ( .A(n67707), .B(n40131), .Y(n40130) );
  INVX1 U41077 ( .A(n67709), .Y(n40131) );
  OR2X1 U41078 ( .A(n40132), .B(n40133), .Y(n65017) );
  INVX1 U41079 ( .A(n64393), .Y(n40132) );
  NOR2X1 U41080 ( .A(n40135), .B(n40136), .Y(n40134) );
  AND2X1 U41081 ( .A(n67501), .B(n67500), .Y(n40135) );
  AND2X1 U41082 ( .A(n67504), .B(n67503), .Y(n40136) );
  AND2X1 U41083 ( .A(n65606), .B(n65605), .Y(n40137) );
  OR2X1 U41084 ( .A(n40138), .B(n40139), .Y(n71733) );
  OR2X1 U41085 ( .A(n71694), .B(n71693), .Y(n40138) );
  NOR2X1 U41086 ( .A(n40141), .B(n67146), .Y(n40140) );
  INVX1 U41087 ( .A(n40140), .Y(n67360) );
  INVX1 U41088 ( .A(n67359), .Y(n40141) );
  OR2X1 U41089 ( .A(n70846), .B(n40142), .Y(n71174) );
  INVX1 U41090 ( .A(n43647), .Y(n40142) );
  NOR2X1 U41091 ( .A(n40144), .B(n40145), .Y(n40143) );
  INVX1 U41092 ( .A(n39576), .Y(n72678) );
  OR2X1 U41093 ( .A(n71432), .B(n71431), .Y(n40144) );
  AND2X1 U41094 ( .A(n38860), .B(n71437), .Y(n40145) );
  OR2X1 U41095 ( .A(n63302), .B(n37407), .Y(n63774) );
  OR2X1 U41096 ( .A(n40146), .B(n40147), .Y(n71212) );
  AND2X1 U41097 ( .A(n70885), .B(n70884), .Y(n40146) );
  AND2X1 U41098 ( .A(n70887), .B(n39629), .Y(n40147) );
  NOR2X1 U41099 ( .A(n40149), .B(n40150), .Y(n40148) );
  OR2X1 U41100 ( .A(n45782), .B(n45781), .Y(n40149) );
  OR2X1 U41101 ( .A(n45793), .B(n45792), .Y(n40150) );
  AND2X1 U41102 ( .A(n64150), .B(n64061), .Y(n40151) );
  INVX1 U41103 ( .A(n40151), .Y(n64447) );
  INVX1 U41104 ( .A(n40525), .Y(n40152) );
  AND2X1 U41105 ( .A(n70164), .B(n70165), .Y(n40153) );
  INVX1 U41106 ( .A(n40153), .Y(n70212) );
  OR2X1 U41107 ( .A(n65366), .B(n65365), .Y(n65739) );
  INVX1 U41108 ( .A(n47621), .Y(n40154) );
  OR2X1 U41109 ( .A(n40615), .B(n40616), .Y(n40155) );
  OR2X1 U41110 ( .A(n40239), .B(n40240), .Y(n40156) );
  AND2X1 U41111 ( .A(n45773), .B(n45772), .Y(n40157) );
  INVX1 U41112 ( .A(n47664), .Y(n40158) );
  OR2X1 U41113 ( .A(n40333), .B(n40161), .Y(n40159) );
  AND2X1 U41114 ( .A(n40159), .B(n40160), .Y(n64585) );
  OR2X1 U41115 ( .A(n40105), .B(n64584), .Y(n40160) );
  OR2X1 U41116 ( .A(n40332), .B(n40105), .Y(n40161) );
  AND2X1 U41117 ( .A(n70513), .B(n70829), .Y(n40162) );
  OR2X1 U41118 ( .A(n41295), .B(n40165), .Y(n40163) );
  AND2X1 U41119 ( .A(n40163), .B(n40164), .Y(n69522) );
  OR2X1 U41120 ( .A(n39855), .B(n68561), .Y(n40164) );
  OR2X1 U41121 ( .A(n41294), .B(n39855), .Y(n40165) );
  NAND2X1 U41122 ( .A(n68445), .B(n68743), .Y(n40166) );
  INVX1 U41123 ( .A(n40167), .Y(n69863) );
  AND2X1 U41124 ( .A(n68236), .B(n68235), .Y(n40168) );
  INVX1 U41125 ( .A(n47685), .Y(n40169) );
  OR2X1 U41126 ( .A(n40170), .B(n40171), .Y(n59976) );
  AND2X1 U41127 ( .A(n60044), .B(n38845), .Y(n40170) );
  AND2X1 U41128 ( .A(n59839), .B(n59838), .Y(n40171) );
  AND2X1 U41129 ( .A(n64661), .B(n64660), .Y(n40172) );
  AND2X1 U41130 ( .A(n70482), .B(n36548), .Y(n40173) );
  AND2X1 U41131 ( .A(n40174), .B(n40175), .Y(n68528) );
  OR2X1 U41132 ( .A(n40176), .B(n68541), .Y(n40175) );
  INVX1 U41133 ( .A(n68544), .Y(n40176) );
  OR2X1 U41134 ( .A(n40177), .B(n40178), .Y(n59553) );
  AND2X1 U41135 ( .A(n59540), .B(n39795), .Y(n40177) );
  AND2X1 U41136 ( .A(n59479), .B(n59478), .Y(n40178) );
  OR2X1 U41137 ( .A(n40231), .B(n40232), .Y(n40179) );
  INVX1 U41138 ( .A(n40179), .Y(n40230) );
  NAND2X1 U41139 ( .A(n68748), .B(n40182), .Y(n40180) );
  NAND2X1 U41140 ( .A(n40180), .B(n40181), .Y(n41383) );
  AND2X1 U41141 ( .A(n68749), .B(n41729), .Y(n40182) );
  OR2X1 U41142 ( .A(n40183), .B(n40184), .Y(n72701) );
  AND2X1 U41143 ( .A(n41454), .B(n72665), .Y(n40183) );
  AND2X1 U41144 ( .A(n41014), .B(n72667), .Y(n40184) );
  INVX1 U41145 ( .A(n62393), .Y(n40185) );
  NOR2X1 U41146 ( .A(n40187), .B(n40188), .Y(n40186) );
  OR2X1 U41147 ( .A(n68919), .B(n68918), .Y(n40187) );
  AND2X1 U41148 ( .A(n68922), .B(n68921), .Y(n40188) );
  OR2X1 U41149 ( .A(n40189), .B(n40190), .Y(n72098) );
  AND2X1 U41150 ( .A(n71418), .B(n43696), .Y(n40189) );
  AND2X1 U41151 ( .A(n41018), .B(n71711), .Y(n40190) );
  INVX1 U41152 ( .A(n40191), .Y(n68759) );
  OR2X1 U41153 ( .A(n38190), .B(n69276), .Y(n69260) );
  AND2X1 U41154 ( .A(n72644), .B(n72645), .Y(n40192) );
  INVX1 U41155 ( .A(n40192), .Y(n72722) );
  OR2X1 U41156 ( .A(n65465), .B(n65466), .Y(n66185) );
  AND2X1 U41157 ( .A(n40193), .B(n40194), .Y(n68052) );
  OR2X1 U41158 ( .A(n67839), .B(n67838), .Y(n40193) );
  AND2X1 U41159 ( .A(n67843), .B(n67842), .Y(n40194) );
  NOR2X1 U41160 ( .A(n40196), .B(n40197), .Y(n40195) );
  INVX1 U41161 ( .A(n40195), .Y(n63110) );
  AND2X1 U41162 ( .A(n36782), .B(n63046), .Y(n40196) );
  AND2X1 U41163 ( .A(n42062), .B(n63050), .Y(n40197) );
  NAND2X1 U41164 ( .A(n63923), .B(n63922), .Y(n40198) );
  AND2X1 U41165 ( .A(n65482), .B(n65641), .Y(n40199) );
  NAND2X1 U41166 ( .A(n64312), .B(n64311), .Y(n40200) );
  AND2X1 U41167 ( .A(n43581), .B(n67855), .Y(n40201) );
  INVX1 U41168 ( .A(n40201), .Y(n68005) );
  NOR2X1 U41169 ( .A(n40203), .B(n65226), .Y(n40202) );
  INVX1 U41170 ( .A(n40202), .Y(n65586) );
  INVX1 U41171 ( .A(n43505), .Y(n40203) );
  NAND2X1 U41172 ( .A(n62348), .B(n62349), .Y(n40204) );
  AND2X1 U41173 ( .A(n40204), .B(n40205), .Y(n62830) );
  AND2X1 U41174 ( .A(n62351), .B(n40206), .Y(n40205) );
  INVX1 U41175 ( .A(n62828), .Y(n40206) );
  OR2X1 U41176 ( .A(n40207), .B(n40208), .Y(n68012) );
  OR2X1 U41177 ( .A(n67301), .B(n67300), .Y(n40207) );
  AND2X1 U41178 ( .A(n67304), .B(n67303), .Y(n40208) );
  OR2X1 U41179 ( .A(n40209), .B(n68751), .Y(n68452) );
  INVX1 U41180 ( .A(n68749), .Y(n40209) );
  OR2X1 U41181 ( .A(n67677), .B(n37356), .Y(n68283) );
  NAND2X1 U41182 ( .A(n67652), .B(n40421), .Y(n40210) );
  OR2X1 U41183 ( .A(n64583), .B(n40211), .Y(n64547) );
  OR2X1 U41184 ( .A(n40105), .B(n43687), .Y(n40211) );
  OR2X1 U41185 ( .A(n40212), .B(n37404), .Y(n65227) );
  AND2X1 U41186 ( .A(n41222), .B(n65588), .Y(n40212) );
  AND2X1 U41187 ( .A(n43506), .B(n38558), .Y(n40213) );
  INVX1 U41188 ( .A(n68835), .Y(n40214) );
  OR2X1 U41189 ( .A(n40422), .B(n69543), .Y(n40215) );
  AND2X1 U41190 ( .A(n67662), .B(n67663), .Y(n40216) );
  AND2X1 U41191 ( .A(n63640), .B(n63639), .Y(n40217) );
  NAND2X1 U41192 ( .A(n63484), .B(n63483), .Y(n40218) );
  OR2X1 U41193 ( .A(n40219), .B(n40220), .Y(n61300) );
  AND2X1 U41194 ( .A(n61431), .B(n36517), .Y(n40219) );
  AND2X1 U41195 ( .A(n42027), .B(n60881), .Y(n40220) );
  OR2X1 U41196 ( .A(n40221), .B(n40222), .Y(n61680) );
  INVX1 U41197 ( .A(n41882), .Y(n40221) );
  AND2X1 U41198 ( .A(n61803), .B(n61679), .Y(n40222) );
  OR2X1 U41199 ( .A(n40223), .B(n40224), .Y(n61684) );
  INVX1 U41200 ( .A(n41891), .Y(n40223) );
  AND2X1 U41201 ( .A(n61800), .B(n61801), .Y(n40224) );
  AND2X1 U41202 ( .A(n41291), .B(n65863), .Y(n40225) );
  INVX1 U41203 ( .A(n40225), .Y(n66862) );
  AND2X1 U41204 ( .A(n64637), .B(n64929), .Y(n40226) );
  AND2X1 U41205 ( .A(n39187), .B(n43559), .Y(n40227) );
  NAND2X1 U41206 ( .A(n38493), .B(n38636), .Y(n40229) );
  AND2X1 U41207 ( .A(n61451), .B(n40289), .Y(n40231) );
  AND2X1 U41208 ( .A(n41986), .B(n61421), .Y(n40232) );
  OR2X1 U41209 ( .A(n40233), .B(n40234), .Y(n61434) );
  INVX1 U41210 ( .A(n42043), .Y(n40233) );
  AND2X1 U41211 ( .A(n40073), .B(n61441), .Y(n40234) );
  OR2X1 U41212 ( .A(n72677), .B(n38047), .Y(n71741) );
  AND2X1 U41213 ( .A(n68596), .B(n68595), .Y(n40235) );
  NOR2X1 U41214 ( .A(n38555), .B(n70527), .Y(n40236) );
  INVX1 U41215 ( .A(n40236), .Y(n70849) );
  AND2X1 U41216 ( .A(n62951), .B(n37373), .Y(n40237) );
  INVX1 U41217 ( .A(n40237), .Y(n63247) );
  NOR2X1 U41218 ( .A(n40239), .B(n40240), .Y(n40238) );
  AND2X1 U41219 ( .A(n61601), .B(n61569), .Y(n40239) );
  AND2X1 U41220 ( .A(n42014), .B(n61571), .Y(n40240) );
  OR2X1 U41221 ( .A(n40419), .B(n40420), .Y(n40241) );
  OR2X1 U41222 ( .A(n40657), .B(n40658), .Y(n40242) );
  NOR2X1 U41223 ( .A(n40244), .B(n40245), .Y(n40243) );
  AND2X1 U41224 ( .A(n60835), .B(n60836), .Y(n40244) );
  AND2X1 U41225 ( .A(n41881), .B(n60837), .Y(n40245) );
  OR2X1 U41226 ( .A(n66056), .B(n40246), .Y(n66091) );
  OR2X1 U41227 ( .A(n66323), .B(n66438), .Y(n40247) );
  INVX1 U41228 ( .A(n40247), .Y(n40287) );
  AND2X1 U41229 ( .A(n42696), .B(n39449), .Y(n40248) );
  AND2X1 U41230 ( .A(n42696), .B(n39449), .Y(n40249) );
  OR2X1 U41231 ( .A(n40250), .B(n40251), .Y(n64530) );
  OR2X1 U41232 ( .A(n64256), .B(n64255), .Y(n40250) );
  AND2X1 U41233 ( .A(n64259), .B(n64258), .Y(n40251) );
  AND2X1 U41234 ( .A(n70160), .B(n70159), .Y(n40252) );
  NOR2X1 U41235 ( .A(n40254), .B(n40255), .Y(n40253) );
  OR2X1 U41236 ( .A(n46082), .B(n46081), .Y(n40254) );
  OR2X1 U41237 ( .A(n46092), .B(n46091), .Y(n40255) );
  OR2X1 U41238 ( .A(n40256), .B(n40257), .Y(n60768) );
  AND2X1 U41239 ( .A(n60525), .B(n37403), .Y(n40256) );
  AND2X1 U41240 ( .A(n60527), .B(n60526), .Y(n40257) );
  INVX1 U41241 ( .A(n43772), .Y(n40258) );
  INVX1 U41242 ( .A(n40258), .Y(n40259) );
  INVX1 U41243 ( .A(n40258), .Y(n40260) );
  OR2X1 U41244 ( .A(n63609), .B(n37412), .Y(n63619) );
  NAND2X1 U41245 ( .A(n65008), .B(n65007), .Y(n40261) );
  AND2X1 U41246 ( .A(n43521), .B(n40955), .Y(n40262) );
  OR2X1 U41247 ( .A(n43656), .B(n70508), .Y(n71105) );
  NOR2X1 U41248 ( .A(n43699), .B(n65585), .Y(n40263) );
  NOR2X1 U41249 ( .A(n40265), .B(n40266), .Y(n40264) );
  AND2X1 U41250 ( .A(n59788), .B(n59610), .Y(n40265) );
  AND2X1 U41251 ( .A(n41759), .B(n59611), .Y(n40266) );
  AND2X1 U41252 ( .A(n67051), .B(n67050), .Y(n40267) );
  OR2X1 U41253 ( .A(n40268), .B(n40269), .Y(n60573) );
  AND2X1 U41254 ( .A(n60186), .B(n60185), .Y(n40268) );
  AND2X1 U41255 ( .A(n60191), .B(n60190), .Y(n40269) );
  AND2X1 U41256 ( .A(n65346), .B(n65347), .Y(n65112) );
  OR2X1 U41257 ( .A(n40270), .B(n40271), .Y(n66585) );
  AND2X1 U41258 ( .A(n41076), .B(n43658), .Y(n40270) );
  AND2X1 U41259 ( .A(n65968), .B(n66262), .Y(n40271) );
  NAND2X1 U41260 ( .A(n65016), .B(n65017), .Y(n40272) );
  INVX1 U41261 ( .A(n48390), .Y(n40273) );
  OR2X1 U41262 ( .A(n67968), .B(n67967), .Y(n40274) );
  AND2X1 U41263 ( .A(n40274), .B(n40275), .Y(n68253) );
  AND2X1 U41264 ( .A(n40276), .B(n41296), .Y(n40275) );
  INVX1 U41265 ( .A(n43635), .Y(n40276) );
  OR2X1 U41266 ( .A(n42832), .B(n42831), .Y(n40277) );
  NAND2X1 U41267 ( .A(n42813), .B(n59135), .Y(n40278) );
  NAND2X1 U41268 ( .A(n63033), .B(n63035), .Y(n40279) );
  NAND2X1 U41269 ( .A(n63033), .B(n63035), .Y(n40280) );
  OR2X1 U41270 ( .A(n40281), .B(n40282), .Y(n59390) );
  AND2X1 U41271 ( .A(n59346), .B(n59347), .Y(n40281) );
  AND2X1 U41272 ( .A(n59349), .B(n59348), .Y(n40282) );
  OR2X1 U41273 ( .A(n40283), .B(n40284), .Y(n64487) );
  OR2X1 U41274 ( .A(n64043), .B(n64042), .Y(n40283) );
  AND2X1 U41275 ( .A(n64225), .B(n64044), .Y(n40284) );
  OR2X1 U41276 ( .A(n40285), .B(n40286), .Y(n64577) );
  OR2X1 U41277 ( .A(n64550), .B(n64549), .Y(n40285) );
  AND2X1 U41278 ( .A(n64552), .B(n64580), .Y(n40286) );
  OR2X1 U41279 ( .A(n38807), .B(n38662), .Y(n46014) );
  OR2X1 U41280 ( .A(n40639), .B(n40640), .Y(n40288) );
  OR2X1 U41281 ( .A(n40609), .B(n40610), .Y(n40289) );
  OR2X1 U41282 ( .A(n40290), .B(n40291), .Y(n59149) );
  AND2X1 U41283 ( .A(n46572), .B(n2468), .Y(n40291) );
  OR2X1 U41284 ( .A(n40292), .B(n40293), .Y(n60776) );
  AND2X1 U41285 ( .A(n60843), .B(n38618), .Y(n40292) );
  AND2X1 U41286 ( .A(n41901), .B(n60510), .Y(n40293) );
  OR2X1 U41287 ( .A(n40294), .B(n39749), .Y(n40533) );
  OR2X1 U41288 ( .A(n63648), .B(n63647), .Y(n40294) );
  INVX1 U41289 ( .A(n40325), .Y(n40295) );
  OR2X1 U41290 ( .A(n40296), .B(n40326), .Y(n66577) );
  NAND2X1 U41291 ( .A(n40295), .B(n66234), .Y(n40296) );
  OR2X1 U41292 ( .A(n40297), .B(n40298), .Y(n59782) );
  AND2X1 U41293 ( .A(n59812), .B(n59810), .Y(n40297) );
  AND2X1 U41294 ( .A(n41809), .B(n59625), .Y(n40298) );
  AND2X1 U41295 ( .A(n40299), .B(n40300), .Y(n72104) );
  OR2X1 U41296 ( .A(n72665), .B(n72100), .Y(n40299) );
  OR2X1 U41297 ( .A(n72666), .B(n72103), .Y(n40300) );
  AND2X1 U41298 ( .A(n70528), .B(n70529), .Y(n40301) );
  OR2X1 U41299 ( .A(n43620), .B(n67961), .Y(n40302) );
  AND2X1 U41300 ( .A(n67981), .B(n40951), .Y(n40303) );
  INVX1 U41301 ( .A(n40303), .Y(n68573) );
  AND2X1 U41302 ( .A(n43676), .B(n72677), .Y(n40304) );
  OR2X1 U41303 ( .A(n40305), .B(n40306), .Y(n63711) );
  AND2X1 U41304 ( .A(n37926), .B(n63427), .Y(n40305) );
  AND2X1 U41305 ( .A(n42094), .B(n63429), .Y(n40306) );
  NAND2X1 U41306 ( .A(n67170), .B(n67510), .Y(n40307) );
  AND2X1 U41307 ( .A(n68740), .B(n68073), .Y(n40308) );
  NAND2X1 U41308 ( .A(n66055), .B(n66091), .Y(n40309) );
  OR2X1 U41309 ( .A(n40310), .B(n40311), .Y(n71171) );
  OR2X1 U41310 ( .A(n40301), .B(n40236), .Y(n40310) );
  AND2X1 U41311 ( .A(n43665), .B(n70852), .Y(n40311) );
  AND2X1 U41312 ( .A(n41266), .B(n39511), .Y(n40312) );
  NAND2X1 U41313 ( .A(n65429), .B(n65086), .Y(n40313) );
  AND2X1 U41314 ( .A(n61584), .B(n61585), .Y(n40315) );
  AND2X1 U41315 ( .A(n42074), .B(n61586), .Y(n40316) );
  NAND2X1 U41316 ( .A(n68005), .B(n41075), .Y(n40317) );
  OR2X1 U41317 ( .A(n68262), .B(n68261), .Y(n40318) );
  OR2X1 U41318 ( .A(n40318), .B(n40319), .Y(n68267) );
  OR2X1 U41319 ( .A(n43539), .B(n40495), .Y(n40319) );
  NAND2X1 U41320 ( .A(n70841), .B(n70840), .Y(n40320) );
  OR2X1 U41321 ( .A(n39797), .B(n43579), .Y(n67193) );
  OR2X1 U41322 ( .A(n40321), .B(n40322), .Y(n64192) );
  OR2X1 U41323 ( .A(n63592), .B(n63591), .Y(n40321) );
  AND2X1 U41324 ( .A(n63595), .B(n63594), .Y(n40322) );
  OR2X1 U41325 ( .A(n38135), .B(n40252), .Y(n70209) );
  OR2X1 U41326 ( .A(n40323), .B(n37367), .Y(n68871) );
  AND2X1 U41327 ( .A(n68883), .B(n68825), .Y(n40323) );
  NOR2X1 U41328 ( .A(n40325), .B(n40326), .Y(n40324) );
  AND2X1 U41329 ( .A(n43676), .B(n65596), .Y(n40325) );
  AND2X1 U41330 ( .A(n65600), .B(n65601), .Y(n40326) );
  NAND2X1 U41331 ( .A(n66438), .B(n66323), .Y(n40327) );
  OR2X1 U41332 ( .A(n40870), .B(n36816), .Y(n40328) );
  OR2X1 U41333 ( .A(n42866), .B(n42694), .Y(n45244) );
  OR2X1 U41334 ( .A(n40329), .B(n40330), .Y(n63685) );
  INVX1 U41335 ( .A(n42113), .Y(n40329) );
  NAND2X1 U41336 ( .A(n66299), .B(n66954), .Y(n40331) );
  OR2X1 U41337 ( .A(n40332), .B(n40333), .Y(n64583) );
  AND2X1 U41338 ( .A(n43676), .B(n63969), .Y(n40332) );
  AND2X1 U41339 ( .A(n63972), .B(n63971), .Y(n40333) );
  NAND2X1 U41340 ( .A(n41122), .B(n40337), .Y(n40334) );
  AND2X1 U41341 ( .A(n40334), .B(n40335), .Y(n66673) );
  OR2X1 U41342 ( .A(n40336), .B(n66079), .Y(n40335) );
  INVX1 U41343 ( .A(n38922), .Y(n40336) );
  AND2X1 U41344 ( .A(n66078), .B(n38922), .Y(n40337) );
  OR2X1 U41345 ( .A(n43528), .B(n40338), .Y(n70210) );
  AND2X1 U41346 ( .A(n41033), .B(n38174), .Y(n40338) );
  OR2X1 U41347 ( .A(n40339), .B(n40340), .Y(n66617) );
  AND2X1 U41348 ( .A(n43561), .B(n66282), .Y(n40339) );
  AND2X1 U41349 ( .A(n66283), .B(n66504), .Y(n40340) );
  OR2X1 U41350 ( .A(n40341), .B(n40342), .Y(n67026) );
  AND2X1 U41351 ( .A(n66441), .B(n66440), .Y(n40341) );
  AND2X1 U41352 ( .A(n66444), .B(n66443), .Y(n40342) );
  OR2X1 U41353 ( .A(n43688), .B(n69551), .Y(n69573) );
  AND2X1 U41354 ( .A(n59402), .B(n59401), .Y(n40343) );
  NOR2X1 U41355 ( .A(n64908), .B(n40345), .Y(n40344) );
  INVX1 U41356 ( .A(n40344), .Y(n65233) );
  INVX1 U41357 ( .A(n43531), .Y(n40345) );
  OR2X1 U41358 ( .A(n40346), .B(n40347), .Y(n59464) );
  AND2X1 U41359 ( .A(n59421), .B(n36524), .Y(n40346) );
  AND2X1 U41360 ( .A(n42160), .B(n59422), .Y(n40347) );
  OR2X1 U41361 ( .A(n40348), .B(n40349), .Y(n68231) );
  OR2X1 U41362 ( .A(n67929), .B(n67928), .Y(n40348) );
  AND2X1 U41363 ( .A(n67932), .B(n43530), .Y(n40349) );
  OR2X1 U41364 ( .A(n39343), .B(n66079), .Y(n67140) );
  OR2X1 U41365 ( .A(n40350), .B(n40351), .Y(n69928) );
  AND2X1 U41366 ( .A(n69866), .B(n69865), .Y(n40350) );
  AND2X1 U41367 ( .A(n43665), .B(n69867), .Y(n40351) );
  OR2X1 U41368 ( .A(n40352), .B(n40353), .Y(n63105) );
  AND2X1 U41369 ( .A(n62824), .B(n62823), .Y(n40352) );
  AND2X1 U41370 ( .A(n42075), .B(n62826), .Y(n40353) );
  AND2X1 U41371 ( .A(n61355), .B(n61354), .Y(n40354) );
  OR2X1 U41372 ( .A(n40355), .B(n40356), .Y(n67285) );
  OR2X1 U41373 ( .A(n36763), .B(n66610), .Y(n40355) );
  AND2X1 U41374 ( .A(n66614), .B(n43624), .Y(n40356) );
  NOR2X1 U41375 ( .A(n40358), .B(n40359), .Y(n40357) );
  AND2X1 U41376 ( .A(n60867), .B(n60868), .Y(n40358) );
  AND2X1 U41377 ( .A(n41972), .B(n60869), .Y(n40359) );
  INVX1 U41378 ( .A(n42897), .Y(n40360) );
  XNOR2X1 U41379 ( .A(n64494), .B(n39014), .Y(n40361) );
  NOR2X1 U41380 ( .A(n40363), .B(n40364), .Y(n40362) );
  AND2X1 U41381 ( .A(n59628), .B(n59626), .Y(n40363) );
  AND2X1 U41382 ( .A(n41812), .B(n59560), .Y(n40364) );
  OR2X1 U41383 ( .A(n43749), .B(n38518), .Y(n59791) );
  OR2X1 U41384 ( .A(n40365), .B(n40366), .Y(n60779) );
  AND2X1 U41385 ( .A(n60781), .B(n39694), .Y(n40365) );
  AND2X1 U41386 ( .A(n41879), .B(n60502), .Y(n40366) );
  OR2X1 U41387 ( .A(n40367), .B(n40368), .Y(n72097) );
  AND2X1 U41388 ( .A(n71708), .B(n71707), .Y(n40368) );
  OR2X1 U41389 ( .A(n40369), .B(n40370), .Y(n67259) );
  OR2X1 U41390 ( .A(n66898), .B(n66897), .Y(n40369) );
  OR2X1 U41391 ( .A(n41413), .B(n66900), .Y(n40370) );
  AND2X1 U41392 ( .A(n61185), .B(n59226), .Y(n40371) );
  INVX1 U41393 ( .A(n40371), .Y(n59227) );
  OR2X1 U41394 ( .A(n40532), .B(n40372), .Y(n46383) );
  NAND2X1 U41395 ( .A(n47422), .B(n40374), .Y(n40372) );
  INVX1 U41396 ( .A(n40373), .Y(n40374) );
  OR2X1 U41397 ( .A(n58820), .B(n40870), .Y(n46570) );
  AND2X1 U41398 ( .A(n59922), .B(n59921), .Y(n40375) );
  OR2X1 U41399 ( .A(n40376), .B(n40377), .Y(n63341) );
  INVX1 U41400 ( .A(n63348), .Y(n40376) );
  AND2X1 U41401 ( .A(n39563), .B(n62869), .Y(n40377) );
  INVX1 U41402 ( .A(n36617), .Y(n40378) );
  OR2X1 U41403 ( .A(n42813), .B(n59135), .Y(n40379) );
  OR2X1 U41404 ( .A(n40380), .B(n40381), .Y(n62824) );
  AND2X1 U41405 ( .A(n62340), .B(n36582), .Y(n40380) );
  AND2X1 U41406 ( .A(n42064), .B(n62341), .Y(n40381) );
  NAND2X1 U41407 ( .A(n39426), .B(n64357), .Y(n40382) );
  NAND2X1 U41408 ( .A(n38493), .B(n38827), .Y(n40383) );
  OR2X1 U41409 ( .A(n40384), .B(n40385), .Y(n66531) );
  OR2X1 U41410 ( .A(n65922), .B(n65921), .Y(n40384) );
  NOR2X1 U41411 ( .A(n65927), .B(n65926), .Y(n40385) );
  NAND2X1 U41412 ( .A(n63685), .B(n40389), .Y(n40386) );
  OR2X1 U41413 ( .A(n40388), .B(n63933), .Y(n40387) );
  INVX1 U41414 ( .A(n63935), .Y(n40388) );
  AND2X1 U41415 ( .A(n63686), .B(n63935), .Y(n40389) );
  NAND2X1 U41416 ( .A(n42376), .B(n36714), .Y(n40390) );
  NAND2X1 U41417 ( .A(n42376), .B(n36714), .Y(n40391) );
  OR2X1 U41418 ( .A(n42784), .B(n45168), .Y(n46231) );
  INVX1 U41419 ( .A(n43473), .Y(n40392) );
  INVX1 U41420 ( .A(n43473), .Y(n40393) );
  NAND2X1 U41421 ( .A(n42221), .B(n40253), .Y(n40394) );
  NOR2X1 U41422 ( .A(n40396), .B(n40397), .Y(n40395) );
  OR2X1 U41423 ( .A(n36790), .B(n70804), .Y(n40396) );
  AND2X1 U41424 ( .A(n70813), .B(n70812), .Y(n40397) );
  INVX1 U41425 ( .A(n40401), .Y(n40398) );
  AND2X1 U41426 ( .A(n59909), .B(n59908), .Y(n40399) );
  OR2X1 U41427 ( .A(n40400), .B(n38062), .Y(n69911) );
  AND2X1 U41428 ( .A(n69571), .B(n69240), .Y(n40400) );
  AND2X1 U41429 ( .A(n39502), .B(n45520), .Y(n40401) );
  INVX1 U41430 ( .A(n40401), .Y(n42671) );
  OR2X1 U41431 ( .A(n40402), .B(n40403), .Y(n63054) );
  AND2X1 U41432 ( .A(n62337), .B(n38499), .Y(n40402) );
  AND2X1 U41433 ( .A(n62339), .B(n42082), .Y(n40403) );
  AND2X1 U41434 ( .A(n40513), .B(n58254), .Y(n40404) );
  NAND2X1 U41435 ( .A(n40123), .B(n70766), .Y(n40405) );
  OR2X1 U41436 ( .A(n40527), .B(n40526), .Y(n40406) );
  OR2X1 U41437 ( .A(n40527), .B(n40526), .Y(n40407) );
  OR2X1 U41438 ( .A(n40408), .B(n40409), .Y(n59535) );
  AND2X1 U41439 ( .A(n59491), .B(n59561), .Y(n40408) );
  AND2X1 U41440 ( .A(n41808), .B(n59492), .Y(n40409) );
  OR2X1 U41441 ( .A(n40410), .B(n40411), .Y(n59538) );
  AND2X1 U41442 ( .A(n59555), .B(n59553), .Y(n40410) );
  AND2X1 U41443 ( .A(n41773), .B(n59482), .Y(n40411) );
  OR2X1 U41444 ( .A(n40412), .B(n40413), .Y(n63424) );
  AND2X1 U41445 ( .A(n63100), .B(n63099), .Y(n40412) );
  AND2X1 U41446 ( .A(n42100), .B(n63103), .Y(n40413) );
  AND2X1 U41447 ( .A(n66607), .B(n66606), .Y(n40414) );
  OR2X1 U41448 ( .A(n68903), .B(n38842), .Y(n69517) );
  NOR2X1 U41449 ( .A(n40416), .B(n40417), .Y(n40415) );
  INVX1 U41450 ( .A(n40415), .Y(n67548) );
  AND2X1 U41451 ( .A(n66877), .B(n66876), .Y(n40416) );
  AND2X1 U41452 ( .A(n66881), .B(n66880), .Y(n40417) );
  INVX1 U41453 ( .A(n69193), .Y(n40418) );
  OR2X1 U41454 ( .A(n38571), .B(n37373), .Y(n63245) );
  OR2X1 U41455 ( .A(n36751), .B(n67650), .Y(n68263) );
  OR2X1 U41456 ( .A(n62961), .B(n62960), .Y(n40419) );
  AND2X1 U41457 ( .A(n62963), .B(n62962), .Y(n40420) );
  NAND2X1 U41458 ( .A(n67651), .B(n68263), .Y(n40421) );
  AND2X1 U41459 ( .A(n41095), .B(n68230), .Y(n40422) );
  INVX1 U41460 ( .A(n49582), .Y(n40423) );
  INVX1 U41461 ( .A(n49582), .Y(n40424) );
  INVX1 U41462 ( .A(n49582), .Y(n40425) );
  INVX1 U41463 ( .A(n49582), .Y(n40426) );
  INVX1 U41464 ( .A(n40423), .Y(n40427) );
  INVX1 U41465 ( .A(n40423), .Y(n40428) );
  OR2X1 U41466 ( .A(n43627), .B(n66507), .Y(n66609) );
  INVX1 U41467 ( .A(n38994), .Y(n40429) );
  OR2X1 U41468 ( .A(n40629), .B(n40630), .Y(n40430) );
  OR2X1 U41469 ( .A(n40431), .B(n37358), .Y(n64686) );
  OR2X1 U41470 ( .A(n41258), .B(n41290), .Y(n40431) );
  INVX1 U41471 ( .A(n49573), .Y(n40432) );
  OR2X1 U41472 ( .A(n40433), .B(n40434), .Y(n61531) );
  AND2X1 U41473 ( .A(n61631), .B(n61527), .Y(n40433) );
  AND2X1 U41474 ( .A(n41877), .B(n61529), .Y(n40434) );
  OR2X1 U41475 ( .A(n40664), .B(n40665), .Y(n40435) );
  AND2X1 U41476 ( .A(n66274), .B(n66275), .Y(n40436) );
  AND2X1 U41477 ( .A(n38781), .B(n65872), .Y(n40437) );
  INVX1 U41478 ( .A(n40437), .Y(n65975) );
  AND2X1 U41479 ( .A(n63917), .B(n63916), .Y(n40438) );
  NAND2X1 U41480 ( .A(n64854), .B(n64853), .Y(n40439) );
  OR2X1 U41481 ( .A(n40441), .B(n40440), .Y(n63649) );
  INVX1 U41482 ( .A(n63145), .Y(n40440) );
  AND2X1 U41483 ( .A(n63143), .B(n63142), .Y(n40441) );
  OR2X1 U41484 ( .A(n40442), .B(n40443), .Y(n66275) );
  AND2X1 U41485 ( .A(n65914), .B(n65913), .Y(n40442) );
  AND2X1 U41486 ( .A(n65915), .B(n43632), .Y(n40443) );
  NOR2X1 U41487 ( .A(n40445), .B(n36757), .Y(n40444) );
  OR2X1 U41488 ( .A(n59127), .B(n59126), .Y(n40445) );
  AND2X1 U41489 ( .A(n42825), .B(n39794), .Y(n40446) );
  AND2X1 U41490 ( .A(n46216), .B(n58254), .Y(n40447) );
  AND2X1 U41491 ( .A(n44988), .B(n42723), .Y(n40448) );
  AND2X1 U41492 ( .A(opcode_opcode_w[18]), .B(n42792), .Y(n40449) );
  OR2X1 U41493 ( .A(n40450), .B(n40451), .Y(n59724) );
  AND2X1 U41494 ( .A(n36442), .B(n39114), .Y(n40450) );
  AND2X1 U41495 ( .A(n59327), .B(n59218), .Y(n40451) );
  INVX1 U41496 ( .A(n42763), .Y(n40453) );
  INVX1 U41497 ( .A(n42761), .Y(n40454) );
  AND2X1 U41498 ( .A(n71715), .B(n72107), .Y(n40455) );
  INVX1 U41499 ( .A(n40455), .Y(n72716) );
  OR2X1 U41500 ( .A(n40456), .B(n72646), .Y(n72719) );
  INVX1 U41501 ( .A(n43707), .Y(n40456) );
  XNOR2X1 U41502 ( .A(n36631), .B(n72104), .Y(n40457) );
  OR2X1 U41503 ( .A(n40458), .B(n40459), .Y(n63629) );
  OR2X1 U41504 ( .A(n62866), .B(n62865), .Y(n40458) );
  AND2X1 U41505 ( .A(n62867), .B(n37379), .Y(n40459) );
  INVX1 U41506 ( .A(n40462), .Y(n40460) );
  INVX1 U41507 ( .A(n43770), .Y(n40461) );
  INVX1 U41508 ( .A(n43770), .Y(n40462) );
  INVX1 U41509 ( .A(n43771), .Y(n40463) );
  INVX1 U41510 ( .A(n43771), .Y(n40464) );
  INVX1 U41511 ( .A(n43771), .Y(n40465) );
  INVX1 U41512 ( .A(n43770), .Y(n40466) );
  INVX1 U41513 ( .A(n43770), .Y(n40467) );
  INVX1 U41514 ( .A(n43770), .Y(n40468) );
  AND2X1 U41515 ( .A(n63527), .B(n63526), .Y(n40469) );
  INVX1 U41516 ( .A(n43748), .Y(n40470) );
  INVX1 U41517 ( .A(n43748), .Y(n40471) );
  INVX1 U41518 ( .A(n43749), .Y(n40472) );
  INVX1 U41519 ( .A(n43749), .Y(n40473) );
  INVX1 U41520 ( .A(n43748), .Y(n40474) );
  INVX1 U41521 ( .A(n43748), .Y(n40475) );
  INVX1 U41522 ( .A(n43748), .Y(n40476) );
  INVX1 U41523 ( .A(n40470), .Y(n40477) );
  AND2X1 U41524 ( .A(n39573), .B(n65364), .Y(n40478) );
  OR2X1 U41525 ( .A(n42881), .B(n40479), .Y(n45507) );
  INVX1 U41526 ( .A(n36707), .Y(n40479) );
  OR2X1 U41527 ( .A(n43636), .B(n67219), .Y(n67872) );
  AND2X1 U41528 ( .A(n38902), .B(n63322), .Y(n40480) );
  AND2X1 U41529 ( .A(n69586), .B(n69585), .Y(n40481) );
  INVX1 U41530 ( .A(n40481), .Y(n69880) );
  INVX1 U41531 ( .A(n43723), .Y(n40482) );
  INVX1 U41532 ( .A(n43722), .Y(n40483) );
  INVX1 U41533 ( .A(n43723), .Y(n40484) );
  INVX1 U41534 ( .A(n43723), .Y(n40485) );
  INVX1 U41535 ( .A(n43723), .Y(n40486) );
  INVX1 U41536 ( .A(n43722), .Y(n40487) );
  INVX1 U41537 ( .A(n43722), .Y(n40488) );
  INVX1 U41538 ( .A(n43722), .Y(n40489) );
  INVX1 U41539 ( .A(n42885), .Y(n40490) );
  NAND2X1 U41540 ( .A(n68963), .B(n69655), .Y(n40491) );
  NOR2X1 U41541 ( .A(n66890), .B(n37362), .Y(n40492) );
  INVX1 U41542 ( .A(n40492), .Y(n67209) );
  NOR2X1 U41543 ( .A(n40494), .B(n40495), .Y(n40493) );
  OR2X1 U41544 ( .A(n68262), .B(n68261), .Y(n40494) );
  AND2X1 U41545 ( .A(n68266), .B(n68265), .Y(n40495) );
  AND2X1 U41546 ( .A(n39614), .B(n60974), .Y(n40496) );
  INVX1 U41547 ( .A(n42222), .Y(n40497) );
  OR2X1 U41548 ( .A(n61531), .B(n61530), .Y(n61532) );
  AND2X1 U41549 ( .A(n45710), .B(n45176), .Y(n40499) );
  AND2X1 U41550 ( .A(n40157), .B(n40148), .Y(n40500) );
  INVX1 U41551 ( .A(n40500), .Y(n71297) );
  OR2X1 U41552 ( .A(n40502), .B(n40501), .Y(n64496) );
  INVX1 U41553 ( .A(n64040), .Y(n40501) );
  OR2X1 U41554 ( .A(n64037), .B(n64036), .Y(n40502) );
  AND2X1 U41555 ( .A(n38128), .B(n71184), .Y(n40503) );
  AND2X1 U41556 ( .A(n67872), .B(n67220), .Y(n40504) );
  AND2X1 U41557 ( .A(n45176), .B(n46014), .Y(n40505) );
  INVX1 U41558 ( .A(n40505), .Y(n49699) );
  OR2X1 U41559 ( .A(n37380), .B(n40506), .Y(n63612) );
  NOR2X1 U41560 ( .A(n63355), .B(n41287), .Y(n40506) );
  INVX1 U41561 ( .A(n36708), .Y(n40507) );
  INVX1 U41562 ( .A(n42486), .Y(n40508) );
  INVX1 U41563 ( .A(n36707), .Y(n40509) );
  INVX1 U41564 ( .A(n42486), .Y(n40510) );
  INVX1 U41565 ( .A(n36708), .Y(n40511) );
  INVX1 U41566 ( .A(n36776), .Y(n40512) );
  INVX1 U41567 ( .A(n36776), .Y(n40513) );
  INVX1 U41568 ( .A(n49599), .Y(n40514) );
  INVX1 U41569 ( .A(n49599), .Y(n40515) );
  OR2X1 U41570 ( .A(n40516), .B(n42814), .Y(n49588) );
  OR2X1 U41571 ( .A(opcode_opcode_w[21]), .B(opcode_opcode_w[20]), .Y(n40516)
         );
  OR2X1 U41572 ( .A(n40532), .B(n46007), .Y(n40517) );
  AND2X1 U41573 ( .A(n68931), .B(n68930), .Y(n40518) );
  OR2X1 U41574 ( .A(n38807), .B(n45181), .Y(n45710) );
  INVX1 U41575 ( .A(n49594), .Y(n40519) );
  INVX1 U41576 ( .A(n49594), .Y(n40520) );
  AND2X1 U41577 ( .A(n40590), .B(n46309), .Y(n40521) );
  NAND2X1 U41578 ( .A(n38652), .B(n62460), .Y(n40522) );
  AND2X1 U41579 ( .A(n44982), .B(opcode_opcode_w[22]), .Y(n40523) );
  OR2X1 U41580 ( .A(n58820), .B(n40479), .Y(n57608) );
  NAND2X1 U41581 ( .A(n38493), .B(n39853), .Y(n40524) );
  AND2X1 U41582 ( .A(n45520), .B(n39501), .Y(n40525) );
  INVX1 U41583 ( .A(n40525), .Y(n45188) );
  OR2X1 U41584 ( .A(n40527), .B(n40526), .Y(n49630) );
  INVX1 U41585 ( .A(n46404), .Y(n40526) );
  OR2X1 U41586 ( .A(n40525), .B(n46235), .Y(n40527) );
  INVX1 U41587 ( .A(n42750), .Y(n40528) );
  OR2X1 U41588 ( .A(n36600), .B(n45200), .Y(n49610) );
  OR2X1 U41589 ( .A(n40529), .B(n42866), .Y(n49582) );
  INVX1 U41590 ( .A(n40523), .Y(n40529) );
  NOR2X1 U41591 ( .A(n40532), .B(n46007), .Y(n40531) );
  OR2X1 U41592 ( .A(n42703), .B(n46024), .Y(n40532) );
  OR2X1 U41593 ( .A(n42807), .B(n42740), .Y(n40534) );
  INVX1 U41594 ( .A(n45871), .Y(n40535) );
  INVX1 U41595 ( .A(n45871), .Y(n40536) );
  AND2X1 U41596 ( .A(n38947), .B(n42770), .Y(n40537) );
  INVX1 U41597 ( .A(n40260), .Y(n40538) );
  OR2X1 U41598 ( .A(n40539), .B(n40540), .Y(n69242) );
  OR2X1 U41599 ( .A(n37367), .B(n68890), .Y(n40539) );
  AND2X1 U41600 ( .A(n43653), .B(n68891), .Y(n40540) );
  OR2X1 U41601 ( .A(n72726), .B(n72725), .Y(n40541) );
  OR2X1 U41602 ( .A(n43718), .B(n72727), .Y(n40542) );
  AND2X1 U41603 ( .A(n40544), .B(n40545), .Y(n40543) );
  INVX1 U41604 ( .A(n40543), .Y(n72820) );
  NOR2X1 U41605 ( .A(n49220), .B(n49219), .Y(n40544) );
  NOR2X1 U41606 ( .A(n49232), .B(n49231), .Y(n40545) );
  AND2X1 U41607 ( .A(n60319), .B(n60440), .Y(n40547) );
  AND2X1 U41608 ( .A(n60165), .B(n60164), .Y(n40548) );
  NOR2X1 U41609 ( .A(n40550), .B(n40551), .Y(n40549) );
  AND2X1 U41610 ( .A(n60872), .B(n60873), .Y(n40550) );
  AND2X1 U41611 ( .A(n41993), .B(n60874), .Y(n40551) );
  AND2X1 U41612 ( .A(n43772), .B(n43456), .Y(n40552) );
  INVX1 U41613 ( .A(n40552), .Y(n59355) );
  AND2X1 U41614 ( .A(n61160), .B(n61159), .Y(n40553) );
  INVX1 U41615 ( .A(n40553), .Y(n62434) );
  AND2X1 U41616 ( .A(n3033), .B(n49685), .Y(n40554) );
  INVX1 U41617 ( .A(n40554), .Y(n47314) );
  OR2X1 U41618 ( .A(n40555), .B(n40556), .Y(n71715) );
  OR2X1 U41619 ( .A(n71712), .B(n40456), .Y(n40555) );
  AND2X1 U41620 ( .A(n71714), .B(n71713), .Y(n40556) );
  OR2X1 U41621 ( .A(n40557), .B(n40558), .Y(n69934) );
  AND2X1 U41622 ( .A(n69603), .B(n43636), .Y(n40557) );
  AND2X1 U41623 ( .A(n69602), .B(n69601), .Y(n40558) );
  OR2X1 U41624 ( .A(n43528), .B(n70836), .Y(n70837) );
  OR2X1 U41625 ( .A(n40559), .B(n40560), .Y(n70517) );
  OR2X1 U41626 ( .A(n38423), .B(n39145), .Y(n40559) );
  AND2X1 U41627 ( .A(n70217), .B(n39186), .Y(n40560) );
  AND2X1 U41628 ( .A(n39255), .B(n43513), .Y(n40561) );
  AND2X1 U41629 ( .A(n70780), .B(n43528), .Y(n40562) );
  XOR2X1 U41630 ( .A(n67703), .B(n41382), .Y(n40563) );
  INVX1 U41631 ( .A(n40563), .Y(n67696) );
  OR2X1 U41632 ( .A(n70478), .B(n40153), .Y(n70766) );
  OR2X1 U41633 ( .A(n40564), .B(n40565), .Y(n71151) );
  OR2X1 U41634 ( .A(n41035), .B(n70843), .Y(n40564) );
  AND2X1 U41635 ( .A(n43521), .B(n40320), .Y(n40565) );
  AND2X1 U41636 ( .A(n70792), .B(n70791), .Y(n40566) );
  XOR2X1 U41637 ( .A(n70857), .B(n70858), .Y(n70872) );
  AND2X1 U41638 ( .A(n70817), .B(n43696), .Y(n40567) );
  NOR2X1 U41639 ( .A(n40567), .B(n40568), .Y(n40571) );
  OR2X1 U41640 ( .A(n40569), .B(n39922), .Y(n40568) );
  AND2X1 U41641 ( .A(n70818), .B(n70819), .Y(n40569) );
  NOR2X1 U41642 ( .A(n40570), .B(n40571), .Y(n41030) );
  INVX1 U41643 ( .A(n71141), .Y(n40570) );
  AND2X1 U41644 ( .A(n59282), .B(n59300), .Y(n59296) );
  AND2X1 U41645 ( .A(n40572), .B(n40573), .Y(n49617) );
  OR2X1 U41646 ( .A(n49610), .B(n36915), .Y(n40572) );
  AND2X1 U41647 ( .A(n49613), .B(n49612), .Y(n40573) );
  AND2X1 U41648 ( .A(n45939), .B(n45938), .Y(n40574) );
  INVX1 U41649 ( .A(n40574), .Y(n60234) );
  OR2X1 U41650 ( .A(n40575), .B(n40576), .Y(n49620) );
  OR2X1 U41651 ( .A(n40833), .B(n40834), .Y(n40575) );
  OR2X1 U41652 ( .A(n49619), .B(n49618), .Y(n40576) );
  OR2X1 U41653 ( .A(n59252), .B(n59253), .Y(n59258) );
  AND2X1 U41654 ( .A(n39680), .B(n40390), .Y(n40577) );
  XNOR2X1 U41655 ( .A(n59495), .B(n59536), .Y(n40578) );
  INVX1 U41656 ( .A(n40578), .Y(n59566) );
  XNOR2X1 U41657 ( .A(writeback_exec_idx_w[0]), .B(n42740), .Y(n40579) );
  INVX1 U41658 ( .A(n40579), .Y(n45266) );
  NOR2X1 U41659 ( .A(n40581), .B(n40582), .Y(n40580) );
  INVX1 U41660 ( .A(n40580), .Y(n59511) );
  AND2X1 U41661 ( .A(n36764), .B(n59496), .Y(n40581) );
  AND2X1 U41662 ( .A(n59498), .B(n59497), .Y(n40582) );
  NOR2X1 U41663 ( .A(n40584), .B(n40585), .Y(n40583) );
  INVX1 U41664 ( .A(n40583), .Y(n59386) );
  AND2X1 U41665 ( .A(n59436), .B(n59364), .Y(n40584) );
  AND2X1 U41666 ( .A(n59366), .B(n59365), .Y(n40585) );
  OR2X1 U41667 ( .A(n46231), .B(n46394), .Y(n49573) );
  OR2X1 U41668 ( .A(n42822), .B(n40371), .Y(n59146) );
  NOR2X1 U41669 ( .A(n40587), .B(n40588), .Y(n40586) );
  INVX1 U41670 ( .A(n40586), .Y(n59949) );
  AND2X1 U41671 ( .A(n59743), .B(n36770), .Y(n40587) );
  AND2X1 U41672 ( .A(n59746), .B(n59745), .Y(n40588) );
  OR2X1 U41673 ( .A(n40589), .B(n43777), .Y(n59689) );
  INVX1 U41674 ( .A(n63222), .Y(n40589) );
  AND2X1 U41675 ( .A(n45176), .B(n45610), .Y(n40590) );
  INVX1 U41676 ( .A(n40590), .Y(n46006) );
  NAND2X1 U41677 ( .A(n47291), .B(n40591), .Y(n42337) );
  NOR2X1 U41678 ( .A(n40592), .B(n47292), .Y(n40591) );
  OR2X1 U41679 ( .A(n47290), .B(n47289), .Y(n40592) );
  NOR2X1 U41680 ( .A(n40604), .B(n42739), .Y(n40593) );
  AND2X1 U41681 ( .A(n42671), .B(n46014), .Y(n40594) );
  INVX1 U41682 ( .A(n40594), .Y(n46726) );
  AND2X1 U41683 ( .A(n60989), .B(n60988), .Y(n40595) );
  INVX1 U41684 ( .A(n40595), .Y(n61215) );
  OR2X1 U41685 ( .A(n60584), .B(n36787), .Y(n60585) );
  AND2X1 U41686 ( .A(n59197), .B(n59200), .Y(n40596) );
  INVX1 U41687 ( .A(n40596), .Y(n59293) );
  AND2X1 U41688 ( .A(n59353), .B(n59350), .Y(n40597) );
  INVX1 U41689 ( .A(n40597), .Y(n59290) );
  XNOR2X1 U41690 ( .A(n36764), .B(n40599), .Y(n40598) );
  OR2X1 U41691 ( .A(n59577), .B(n59576), .Y(n40599) );
  OR2X1 U41692 ( .A(n40600), .B(n40407), .Y(n46314) );
  NOR2X1 U41693 ( .A(n40602), .B(n40603), .Y(n40601) );
  AND2X1 U41694 ( .A(n59688), .B(n59690), .Y(n40602) );
  AND2X1 U41695 ( .A(n59693), .B(n59692), .Y(n40603) );
  OR2X1 U41696 ( .A(n40604), .B(n42740), .Y(n46927) );
  OR2X1 U41697 ( .A(opcode_opcode_w[21]), .B(n42814), .Y(n40604) );
  AND2X1 U41698 ( .A(n63347), .B(n62868), .Y(n40605) );
  INVX1 U41699 ( .A(n40605), .Y(n63340) );
  AND2X1 U41700 ( .A(n43773), .B(n44070), .Y(n40606) );
  INVX1 U41701 ( .A(n40606), .Y(n59395) );
  AND2X1 U41702 ( .A(n42750), .B(n42761), .Y(n40607) );
  NOR2X1 U41703 ( .A(n40609), .B(n40610), .Y(n40608) );
  AND2X1 U41704 ( .A(n61417), .B(n61418), .Y(n40609) );
  AND2X1 U41705 ( .A(n41976), .B(n61419), .Y(n40610) );
  NOR2X1 U41706 ( .A(n40612), .B(n40613), .Y(n40611) );
  AND2X1 U41707 ( .A(n60498), .B(n60784), .Y(n40612) );
  AND2X1 U41708 ( .A(n60783), .B(n60500), .Y(n40613) );
  NOR2X1 U41709 ( .A(n40615), .B(n40616), .Y(n40614) );
  AND2X1 U41710 ( .A(n60246), .B(n38695), .Y(n40615) );
  AND2X1 U41711 ( .A(n60249), .B(n60248), .Y(n40616) );
  OR2X1 U41712 ( .A(n60011), .B(n36786), .Y(n59809) );
  OR2X1 U41713 ( .A(n40617), .B(n40618), .Y(n47336) );
  OR2X1 U41714 ( .A(n47335), .B(n47334), .Y(n40617) );
  AND2X1 U41715 ( .A(n3025), .B(n57613), .Y(n40618) );
  INVX1 U41716 ( .A(n40619), .Y(n59244) );
  XNOR2X1 U41717 ( .A(n36787), .B(n40621), .Y(n40620) );
  INVX1 U41718 ( .A(n40620), .Y(n60582) );
  XOR2X1 U41719 ( .A(n60584), .B(n41499), .Y(n40621) );
  NOR2X1 U41720 ( .A(n40623), .B(n40624), .Y(n40622) );
  AND2X1 U41721 ( .A(n59511), .B(n59512), .Y(n40623) );
  AND2X1 U41722 ( .A(n59514), .B(n59513), .Y(n40624) );
  AND2X1 U41723 ( .A(n59798), .B(n59797), .Y(n40625) );
  INVX1 U41724 ( .A(n40625), .Y(n60005) );
  OR2X1 U41725 ( .A(n59231), .B(n39714), .Y(n59686) );
  OR2X1 U41726 ( .A(n39017), .B(n60319), .Y(n60164) );
  NOR2X1 U41727 ( .A(n43459), .B(n43778), .Y(n40626) );
  INVX1 U41728 ( .A(n40626), .Y(n59684) );
  INVX1 U41729 ( .A(n43456), .Y(n40627) );
  NOR2X1 U41730 ( .A(n40629), .B(n40630), .Y(n40628) );
  AND2X1 U41731 ( .A(n59211), .B(n59212), .Y(n40629) );
  AND2X1 U41732 ( .A(n59214), .B(n59213), .Y(n40630) );
  OR2X1 U41733 ( .A(n40631), .B(n59147), .Y(n59124) );
  OR2X1 U41734 ( .A(n59148), .B(n59149), .Y(n40631) );
  NOR2X1 U41735 ( .A(n40633), .B(n40634), .Y(n40632) );
  INVX1 U41736 ( .A(n40632), .Y(n60847) );
  AND2X1 U41737 ( .A(n61324), .B(n60844), .Y(n40633) );
  AND2X1 U41738 ( .A(n41913), .B(n60846), .Y(n40634) );
  NOR2X1 U41739 ( .A(n40636), .B(n40637), .Y(n40635) );
  INVX1 U41740 ( .A(n40635), .Y(n60102) );
  AND2X1 U41741 ( .A(n60133), .B(n60134), .Y(n40636) );
  AND2X1 U41742 ( .A(n41819), .B(n60010), .Y(n40637) );
  NOR2X1 U41743 ( .A(n40639), .B(n40640), .Y(n40638) );
  AND2X1 U41744 ( .A(n59308), .B(n59309), .Y(n40639) );
  AND2X1 U41745 ( .A(n59311), .B(n59310), .Y(n40640) );
  OR2X1 U41746 ( .A(n59597), .B(n40598), .Y(n59578) );
  AND2X1 U41747 ( .A(n3024), .B(n40537), .Y(n40641) );
  INVX1 U41748 ( .A(n40641), .Y(n47332) );
  OR2X1 U41749 ( .A(n59785), .B(n59619), .Y(n59620) );
  OR2X1 U41750 ( .A(n36600), .B(n42866), .Y(n49605) );
  OR2X1 U41751 ( .A(n45255), .B(n45619), .Y(n42780) );
  OR2X1 U41752 ( .A(n40642), .B(n49610), .Y(n47328) );
  NOR2X1 U41753 ( .A(n40644), .B(n40645), .Y(n40643) );
  AND2X1 U41754 ( .A(n60370), .B(n60368), .Y(n40644) );
  AND2X1 U41755 ( .A(n41851), .B(n60140), .Y(n40645) );
  XOR2X1 U41756 ( .A(n63612), .B(n63146), .Y(n63626) );
  AND2X1 U41757 ( .A(n59866), .B(n59865), .Y(n40646) );
  OR2X1 U41758 ( .A(n40647), .B(n40648), .Y(n59697) );
  INVX1 U41759 ( .A(n41779), .Y(n40647) );
  AND2X1 U41760 ( .A(n40662), .B(n59696), .Y(n40648) );
  OR2X1 U41761 ( .A(n59648), .B(n59649), .Y(n59650) );
  OR2X1 U41762 ( .A(n38807), .B(n38661), .Y(n46019) );
  NOR2X1 U41763 ( .A(n40650), .B(n40651), .Y(n40649) );
  AND2X1 U41764 ( .A(n59827), .B(n60031), .Y(n40650) );
  AND2X1 U41765 ( .A(n41869), .B(n59829), .Y(n40651) );
  AND2X1 U41766 ( .A(n2233), .B(n39318), .Y(n40652) );
  INVX1 U41767 ( .A(n40652), .Y(n47274) );
  NOR2X1 U41768 ( .A(n40654), .B(n40655), .Y(n40653) );
  INVX1 U41769 ( .A(n40653), .Y(n59601) );
  AND2X1 U41770 ( .A(n59618), .B(n59616), .Y(n40654) );
  AND2X1 U41771 ( .A(n41774), .B(n59552), .Y(n40655) );
  NOR2X1 U41772 ( .A(n40657), .B(n40658), .Y(n40656) );
  AND2X1 U41773 ( .A(n59735), .B(n38765), .Y(n40657) );
  AND2X1 U41774 ( .A(n59740), .B(n59739), .Y(n40658) );
  NOR2X1 U41775 ( .A(n40660), .B(n40661), .Y(n40659) );
  INVX1 U41776 ( .A(n40659), .Y(n59985) );
  AND2X1 U41777 ( .A(n36786), .B(n60011), .Y(n40660) );
  AND2X1 U41778 ( .A(n41815), .B(n59809), .Y(n40661) );
  AND2X1 U41779 ( .A(n59223), .B(n59222), .Y(n40662) );
  INVX1 U41780 ( .A(n40662), .Y(n59694) );
  NOR2X1 U41781 ( .A(n40664), .B(n40665), .Y(n40663) );
  AND2X1 U41782 ( .A(n59925), .B(n59923), .Y(n40664) );
  AND2X1 U41783 ( .A(n59928), .B(n59927), .Y(n40665) );
  NOR2X1 U41784 ( .A(n40667), .B(n40668), .Y(n40666) );
  AND2X1 U41785 ( .A(n59632), .B(n59819), .Y(n40667) );
  AND2X1 U41786 ( .A(n41839), .B(n59634), .Y(n40668) );
  INVX1 U41787 ( .A(n15442), .Y(n40669) );
  INVX1 U41788 ( .A(n43567), .Y(n40670) );
  AND2X1 U41789 ( .A(n57893), .B(n55820), .Y(n56763) );
  INVX1 U41790 ( .A(n56763), .Y(n40671) );
  INVX1 U41791 ( .A(n56763), .Y(n40672) );
  INVX1 U41792 ( .A(n56763), .Y(n40673) );
  INVX1 U41793 ( .A(n73510), .Y(n40674) );
  AND2X1 U41794 ( .A(n57993), .B(n58179), .Y(n58084) );
  INVX1 U41795 ( .A(n58084), .Y(n40675) );
  INVX1 U41796 ( .A(n58084), .Y(n40676) );
  INVX1 U41797 ( .A(n58084), .Y(n40677) );
  NAND2X1 U41798 ( .A(n16342), .B(n73572), .Y(n40678) );
  NAND2X1 U41799 ( .A(n56998), .B(n56824), .Y(n40679) );
  NAND2X1 U41800 ( .A(n56998), .B(n56824), .Y(n40680) );
  AND2X1 U41801 ( .A(n73539), .B(n73503), .Y(n24967) );
  INVX1 U41802 ( .A(n24967), .Y(n40681) );
  INVX1 U41803 ( .A(n24967), .Y(n40682) );
  INVX1 U41804 ( .A(n43615), .Y(n40683) );
  INVX1 U41805 ( .A(n58576), .Y(n40684) );
  NAND2X1 U41806 ( .A(n45520), .B(n39502), .Y(n40685) );
  AND2X1 U41807 ( .A(n55820), .B(n57895), .Y(n56764) );
  INVX1 U41808 ( .A(n56764), .Y(n40686) );
  INVX1 U41809 ( .A(n56764), .Y(n40687) );
  INVX1 U41810 ( .A(n56764), .Y(n40688) );
  AND2X1 U41811 ( .A(n57316), .B(n73523), .Y(n58761) );
  INVX1 U41812 ( .A(n58761), .Y(n40689) );
  INVX1 U41813 ( .A(n58761), .Y(n40690) );
  INVX1 U41814 ( .A(n58761), .Y(n40691) );
  AND2X1 U41815 ( .A(n57991), .B(n58179), .Y(n58078) );
  INVX1 U41816 ( .A(n58078), .Y(n40692) );
  INVX1 U41817 ( .A(n58078), .Y(n40693) );
  INVX1 U41818 ( .A(n58078), .Y(n40694) );
  AND2X1 U41819 ( .A(n40695), .B(n40952), .Y(n40944) );
  INVX1 U41820 ( .A(n71697), .Y(n40695) );
  NOR2X1 U41821 ( .A(n41013), .B(n40227), .Y(n69197) );
  NOR2X1 U41822 ( .A(n66509), .B(n40696), .Y(n66610) );
  NAND2X1 U41823 ( .A(n66609), .B(n66608), .Y(n40696) );
  NOR2X1 U41824 ( .A(n41081), .B(n40697), .Y(n70207) );
  NAND2X1 U41825 ( .A(n70206), .B(n70205), .Y(n40697) );
  NOR2X1 U41826 ( .A(n41059), .B(n40698), .Y(n67928) );
  INVX1 U41827 ( .A(n67927), .Y(n40698) );
  XNOR2X1 U41828 ( .A(n40699), .B(n70438), .Y(n70889) );
  NOR2X1 U41829 ( .A(n70241), .B(n39962), .Y(n40699) );
  XOR2X1 U41830 ( .A(n71182), .B(n71172), .Y(n71177) );
  AND2X1 U41831 ( .A(n40700), .B(n40701), .Y(n60217) );
  NAND2X1 U41832 ( .A(n60212), .B(n36734), .Y(n40700) );
  NAND2X1 U41833 ( .A(n60215), .B(n60214), .Y(n40701) );
  NOR2X1 U41834 ( .A(n40702), .B(n41163), .Y(n67924) );
  INVX1 U41835 ( .A(n67922), .Y(n40702) );
  XNOR2X1 U41836 ( .A(n40703), .B(n40704), .Y(n70144) );
  NOR2X1 U41837 ( .A(n69624), .B(n69623), .Y(n40703) );
  XNOR2X1 U41838 ( .A(n70136), .B(n71794), .Y(n40704) );
  XNOR2X1 U41839 ( .A(n41030), .B(n37393), .Y(n71126) );
  XNOR2X1 U41840 ( .A(n41010), .B(n40705), .Y(n71109) );
  XOR2X1 U41841 ( .A(n70508), .B(n70476), .Y(n40705) );
  XNOR2X1 U41842 ( .A(n40706), .B(n68494), .Y(n68590) );
  NOR2X1 U41843 ( .A(n68269), .B(n68270), .Y(n40706) );
  AND2X1 U41844 ( .A(n40707), .B(n40708), .Y(n41023) );
  NAND2X1 U41845 ( .A(n69210), .B(n69209), .Y(n40708) );
  XOR2X1 U41846 ( .A(n71115), .B(n40709), .Y(n41028) );
  XNOR2X1 U41847 ( .A(n71114), .B(n43679), .Y(n40709) );
  NOR2X1 U41848 ( .A(n68581), .B(n68580), .Y(n40710) );
  NAND2X1 U41849 ( .A(n40711), .B(n43523), .Y(n70211) );
  INVX1 U41850 ( .A(n70209), .Y(n40711) );
  XOR2X1 U41851 ( .A(n40712), .B(n40986), .Y(n70543) );
  XNOR2X1 U41852 ( .A(n70888), .B(n70542), .Y(n40712) );
  NAND2X1 U41853 ( .A(n40713), .B(n71724), .Y(n71413) );
  XNOR2X1 U41854 ( .A(n71413), .B(n36778), .Y(n71422) );
  XNOR2X1 U41855 ( .A(n40714), .B(n69540), .Y(n70167) );
  INVX1 U41856 ( .A(n69885), .Y(n40714) );
  XOR2X1 U41857 ( .A(n71176), .B(n40715), .Y(n71748) );
  XNOR2X1 U41858 ( .A(n71168), .B(n71172), .Y(n40715) );
  INVX1 U41859 ( .A(n66576), .Y(n40716) );
  NOR2X1 U41860 ( .A(n40717), .B(n40718), .Y(n65601) );
  INVX1 U41861 ( .A(n65595), .Y(n40717) );
  NOR2X1 U41862 ( .A(n43678), .B(n65596), .Y(n40718) );
  NAND2X1 U41863 ( .A(n43665), .B(n40719), .Y(n68559) );
  INVX1 U41864 ( .A(n68249), .Y(n40719) );
  XOR2X1 U41865 ( .A(n60213), .B(n40720), .Y(n59926) );
  NOR2X1 U41866 ( .A(n59723), .B(n59722), .Y(n40720) );
  XOR2X1 U41867 ( .A(n68241), .B(n40721), .Y(n68245) );
  XNOR2X1 U41868 ( .A(n68243), .B(n68242), .Y(n40721) );
  XOR2X1 U41869 ( .A(n67860), .B(n40722), .Y(n67869) );
  XNOR2X1 U41870 ( .A(n70560), .B(n38725), .Y(n40722) );
  XOR2X1 U41871 ( .A(n66617), .B(n40723), .Y(n66887) );
  XNOR2X1 U41872 ( .A(n66616), .B(n67993), .Y(n40723) );
  XOR2X1 U41873 ( .A(n65552), .B(n40724), .Y(n65557) );
  XNOR2X1 U41874 ( .A(n65553), .B(n43523), .Y(n40724) );
  XOR2X1 U41875 ( .A(n64217), .B(n40725), .Y(n64045) );
  XNOR2X1 U41876 ( .A(n63870), .B(n64202), .Y(n40725) );
  NAND2X1 U41877 ( .A(n43677), .B(n40726), .Y(n66573) );
  INVX1 U41878 ( .A(n66255), .Y(n40726) );
  XOR2X1 U41879 ( .A(n70589), .B(n40727), .Y(n70729) );
  NOR2X1 U41880 ( .A(n70419), .B(n70418), .Y(n40727) );
  NAND2X1 U41881 ( .A(n43506), .B(n40728), .Y(n66921) );
  INVX1 U41882 ( .A(n66572), .Y(n40728) );
  NOR2X1 U41883 ( .A(n40729), .B(n40730), .Y(n68395) );
  INVX1 U41884 ( .A(n68402), .Y(n40729) );
  NAND2X1 U41885 ( .A(n68401), .B(n68130), .Y(n40730) );
  XOR2X1 U41886 ( .A(n67595), .B(n40731), .Y(n67244) );
  XNOR2X1 U41887 ( .A(n67606), .B(n43693), .Y(n40731) );
  XOR2X1 U41888 ( .A(n63971), .B(n40732), .Y(n64274) );
  XNOR2X1 U41889 ( .A(n63969), .B(n43678), .Y(n40732) );
  XOR2X1 U41890 ( .A(n69044), .B(n40733), .Y(n68692) );
  XNOR2X1 U41891 ( .A(n68687), .B(n69041), .Y(n40733) );
  XOR2X1 U41892 ( .A(n40734), .B(n66375), .Y(n66743) );
  XNOR2X1 U41893 ( .A(n66366), .B(n66723), .Y(n40734) );
  NOR2X1 U41894 ( .A(n40735), .B(n40736), .Y(n70328) );
  INVX1 U41895 ( .A(n70321), .Y(n40735) );
  NAND2X1 U41896 ( .A(n70326), .B(n70325), .Y(n40736) );
  OR2X1 U41897 ( .A(n59336), .B(n36771), .Y(n59371) );
  XOR2X1 U41898 ( .A(n40737), .B(n66984), .Y(n66972) );
  XNOR2X1 U41899 ( .A(n66472), .B(n66471), .Y(n40737) );
  XNOR2X1 U41900 ( .A(n66963), .B(n40738), .Y(n67546) );
  XOR2X1 U41901 ( .A(n66849), .B(n66848), .Y(n40738) );
  XOR2X1 U41902 ( .A(n69205), .B(n40739), .Y(n69514) );
  NOR2X1 U41903 ( .A(n68925), .B(n68926), .Y(n40739) );
  AND2X1 U41904 ( .A(n40415), .B(n66946), .Y(n41319) );
  XNOR2X1 U41905 ( .A(n63353), .B(n40740), .Y(n62864) );
  XNOR2X1 U41906 ( .A(n63355), .B(n63356), .Y(n40740) );
  NOR2X1 U41907 ( .A(n67272), .B(n43672), .Y(n40741) );
  NAND2X1 U41908 ( .A(n67634), .B(n67631), .Y(n40742) );
  NAND2X1 U41909 ( .A(n40743), .B(n40744), .Y(n70161) );
  NAND2X1 U41910 ( .A(n69595), .B(n69594), .Y(n40743) );
  NAND2X1 U41911 ( .A(n69596), .B(n43656), .Y(n40744) );
  XNOR2X1 U41912 ( .A(n68928), .B(n43542), .Y(n40745) );
  NOR2X1 U41913 ( .A(n40746), .B(n40747), .Y(n41352) );
  INVX1 U41914 ( .A(n70155), .Y(n40746) );
  AND2X1 U41915 ( .A(n70154), .B(n70153), .Y(n40747) );
  XOR2X1 U41916 ( .A(n67630), .B(n40748), .Y(n41320) );
  XNOR2X1 U41917 ( .A(n67629), .B(n67869), .Y(n40748) );
  OR2X1 U41918 ( .A(n36716), .B(n40749), .Y(n64972) );
  NAND2X1 U41919 ( .A(n64692), .B(n64691), .Y(n40749) );
  XNOR2X1 U41920 ( .A(n63014), .B(n40750), .Y(n62509) );
  NOR2X1 U41921 ( .A(n62408), .B(n62407), .Y(n40750) );
  NAND2X1 U41922 ( .A(n40752), .B(n40751), .Y(n63992) );
  INVX1 U41923 ( .A(n63991), .Y(n40751) );
  NAND2X1 U41924 ( .A(n40753), .B(n40754), .Y(n59848) );
  NAND2X1 U41925 ( .A(n59977), .B(n59976), .Y(n40753) );
  NAND2X1 U41926 ( .A(n59975), .B(n59843), .Y(n40754) );
  XOR2X1 U41927 ( .A(n67218), .B(n40755), .Y(n41368) );
  XNOR2X1 U41928 ( .A(n67217), .B(n43633), .Y(n40755) );
  NOR2X1 U41929 ( .A(n40756), .B(n61063), .Y(n61064) );
  INVX1 U41930 ( .A(n61066), .Y(n40756) );
  XOR2X1 U41931 ( .A(n64677), .B(n40757), .Y(n64668) );
  XNOR2X1 U41932 ( .A(n64502), .B(n64675), .Y(n40757) );
  XOR2X1 U41933 ( .A(n40758), .B(n66799), .Y(n66816) );
  XNOR2X1 U41934 ( .A(n66798), .B(n41407), .Y(n40758) );
  XOR2X1 U41935 ( .A(n68986), .B(n40759), .Y(n68964) );
  XNOR2X1 U41936 ( .A(n69450), .B(n68991), .Y(n40759) );
  XNOR2X1 U41937 ( .A(n40760), .B(n41352), .Y(n70458) );
  XNOR2X1 U41938 ( .A(n70215), .B(n43633), .Y(n40760) );
  NAND2X1 U41939 ( .A(n40761), .B(n44000), .Y(n65493) );
  INVX1 U41940 ( .A(n65159), .Y(n40761) );
  XNOR2X1 U41941 ( .A(n64512), .B(n38129), .Y(n40762) );
  XOR2X1 U41942 ( .A(n40763), .B(n68934), .Y(n68785) );
  XNOR2X1 U41943 ( .A(n68932), .B(n43593), .Y(n40763) );
  XOR2X1 U41944 ( .A(n40764), .B(n64990), .Y(n65315) );
  XNOR2X1 U41945 ( .A(n64983), .B(n64989), .Y(n40764) );
  XOR2X1 U41946 ( .A(n65099), .B(n65110), .Y(n40765) );
  NAND2X1 U41947 ( .A(n40766), .B(n43549), .Y(n67203) );
  INVX1 U41948 ( .A(n66526), .Y(n40766) );
  XNOR2X1 U41949 ( .A(n64369), .B(n40767), .Y(n64201) );
  XOR2X1 U41950 ( .A(n64825), .B(n64200), .Y(n40767) );
  AND2X1 U41951 ( .A(n40768), .B(n66187), .Y(n41376) );
  NAND2X1 U41952 ( .A(n65464), .B(n65463), .Y(n40768) );
  XOR2X1 U41953 ( .A(n40769), .B(n65303), .Y(n41435) );
  XNOR2X1 U41954 ( .A(n65305), .B(n65304), .Y(n40769) );
  NOR2X1 U41955 ( .A(n43714), .B(n40982), .Y(n40770) );
  NAND2X1 U41956 ( .A(n43705), .B(n68529), .Y(n40771) );
  NAND2X1 U41957 ( .A(n68530), .B(n68531), .Y(n40772) );
  XOR2X1 U41958 ( .A(n40773), .B(n66755), .Y(n66362) );
  XNOR2X1 U41959 ( .A(n66745), .B(n66143), .Y(n40773) );
  XOR2X1 U41960 ( .A(n40774), .B(n70033), .Y(n70047) );
  XNOR2X1 U41961 ( .A(n70023), .B(n69784), .Y(n40774) );
  XOR2X1 U41962 ( .A(n40775), .B(n66139), .Y(n66384) );
  XNOR2X1 U41963 ( .A(n66123), .B(n71847), .Y(n40775) );
  NOR2X1 U41964 ( .A(n40776), .B(n40777), .Y(n69131) );
  INVX1 U41965 ( .A(n69125), .Y(n40776) );
  NOR2X1 U41966 ( .A(n69126), .B(n69127), .Y(n40777) );
  XOR2X1 U41967 ( .A(n40778), .B(n68351), .Y(n68379) );
  XNOR2X1 U41968 ( .A(n68358), .B(n41515), .Y(n40778) );
  NOR2X1 U41969 ( .A(n68661), .B(n40779), .Y(n68668) );
  NAND2X1 U41970 ( .A(n68667), .B(n68666), .Y(n40779) );
  XOR2X1 U41971 ( .A(n70990), .B(n40780), .Y(n71028) );
  NOR2X1 U41972 ( .A(n70659), .B(n70658), .Y(n40780) );
  NAND2X1 U41973 ( .A(n66019), .B(n36586), .Y(n40781) );
  XOR2X1 U41974 ( .A(n40782), .B(n64345), .Y(n64497) );
  XNOR2X1 U41975 ( .A(n64344), .B(n64346), .Y(n40782) );
  XOR2X1 U41976 ( .A(n40783), .B(n64039), .Y(n64028) );
  XNOR2X1 U41977 ( .A(n64038), .B(n41566), .Y(n40783) );
  XOR2X1 U41978 ( .A(n64312), .B(n40784), .Y(n63990) );
  XNOR2X1 U41979 ( .A(n64645), .B(n64311), .Y(n40784) );
  XOR2X1 U41980 ( .A(n66205), .B(n40785), .Y(n66032) );
  XNOR2X1 U41981 ( .A(n66023), .B(n66207), .Y(n40785) );
  XOR2X1 U41982 ( .A(n40786), .B(n62535), .Y(n62368) );
  XNOR2X1 U41983 ( .A(n62537), .B(n62534), .Y(n40786) );
  XOR2X1 U41984 ( .A(n63461), .B(n40787), .Y(n63905) );
  XNOR2X1 U41985 ( .A(n63462), .B(n41992), .Y(n40787) );
  XOR2X1 U41986 ( .A(n64866), .B(n64865), .Y(n41609) );
  XOR2X1 U41987 ( .A(n68067), .B(n40788), .Y(n68739) );
  XNOR2X1 U41988 ( .A(n68178), .B(n68179), .Y(n40788) );
  XNOR2X1 U41989 ( .A(n40789), .B(n65269), .Y(n65174) );
  XOR2X1 U41990 ( .A(n42067), .B(n65257), .Y(n40789) );
  XOR2X1 U41991 ( .A(n40790), .B(n69817), .Y(n41638) );
  NOR2X1 U41992 ( .A(n69652), .B(n69651), .Y(n40790) );
  XOR2X1 U41993 ( .A(n63988), .B(n40791), .Y(n64299) );
  XNOR2X1 U41994 ( .A(n63925), .B(n63924), .Y(n40791) );
  XOR2X1 U41995 ( .A(n40792), .B(n59743), .Y(n59749) );
  XNOR2X1 U41996 ( .A(n59744), .B(n36770), .Y(n40792) );
  XOR2X1 U41997 ( .A(n63743), .B(n40793), .Y(n41644) );
  XNOR2X1 U41998 ( .A(n63653), .B(n63652), .Y(n40793) );
  NAND2X1 U41999 ( .A(n40795), .B(n40794), .Y(n62378) );
  NAND2X1 U42000 ( .A(n41930), .B(n61265), .Y(n40794) );
  NAND2X1 U42001 ( .A(n61267), .B(n61266), .Y(n40795) );
  XOR2X1 U42002 ( .A(n40796), .B(n66997), .Y(n41633) );
  XNOR2X1 U42003 ( .A(n67011), .B(n67520), .Y(n40796) );
  XOR2X1 U42004 ( .A(n61117), .B(n40797), .Y(n61100) );
  XNOR2X1 U42005 ( .A(n61078), .B(n61077), .Y(n40797) );
  XOR2X1 U42006 ( .A(n63430), .B(n40798), .Y(n63428) );
  XNOR2X1 U42007 ( .A(n63434), .B(n42078), .Y(n40798) );
  XOR2X1 U42008 ( .A(n64301), .B(n40799), .Y(n63986) );
  XNOR2X1 U42009 ( .A(n64299), .B(n64296), .Y(n40799) );
  NOR2X1 U42010 ( .A(n40800), .B(n65352), .Y(n64995) );
  INVX1 U42011 ( .A(n65353), .Y(n40800) );
  XOR2X1 U42012 ( .A(n59419), .B(n40801), .Y(n59420) );
  NOR2X1 U42013 ( .A(n59418), .B(n59417), .Y(n40801) );
  XOR2X1 U42014 ( .A(n63667), .B(n40802), .Y(n63675) );
  XNOR2X1 U42015 ( .A(n63668), .B(n42032), .Y(n40802) );
  XOR2X1 U42016 ( .A(n66832), .B(n40803), .Y(n66664) );
  XNOR2X1 U42017 ( .A(n66833), .B(n66834), .Y(n40803) );
  XOR2X1 U42018 ( .A(n40279), .B(n40804), .Y(n62364) );
  XNOR2X1 U42019 ( .A(n63034), .B(n63032), .Y(n40804) );
  XNOR2X1 U42020 ( .A(n40805), .B(n71630), .Y(n71631) );
  XOR2X1 U42021 ( .A(n71629), .B(n41664), .Y(n40805) );
  XOR2X1 U42022 ( .A(n71487), .B(n40806), .Y(n71479) );
  XNOR2X1 U42023 ( .A(n42998), .B(n71596), .Y(n40806) );
  XOR2X1 U42024 ( .A(n40807), .B(n65390), .Y(n65388) );
  XNOR2X1 U42025 ( .A(n65378), .B(n65392), .Y(n40807) );
  NAND2X1 U42026 ( .A(n41532), .B(n40808), .Y(n49804) );
  NAND2X1 U42027 ( .A(n49803), .B(n49802), .Y(n40808) );
  NAND2X1 U42028 ( .A(n40552), .B(n59356), .Y(n59350) );
  XNOR2X1 U42029 ( .A(n64982), .B(n40809), .Y(n64977) );
  XOR2X1 U42030 ( .A(n64979), .B(n64981), .Y(n40809) );
  NOR2X1 U42031 ( .A(n40810), .B(n65294), .Y(n65302) );
  INVX1 U42032 ( .A(n65299), .Y(n40810) );
  XOR2X1 U42033 ( .A(n63602), .B(n40811), .Y(n63336) );
  XNOR2X1 U42034 ( .A(n63599), .B(n63477), .Y(n40811) );
  NAND2X1 U42035 ( .A(n40812), .B(n40813), .Y(n69448) );
  INVX1 U42036 ( .A(n68619), .Y(n40812) );
  NAND2X1 U42037 ( .A(n68626), .B(n68625), .Y(n40813) );
  XNOR2X1 U42038 ( .A(n59339), .B(n40814), .Y(n59419) );
  XNOR2X1 U42039 ( .A(n59355), .B(n59338), .Y(n40814) );
  XOR2X1 U42040 ( .A(n64777), .B(n40815), .Y(n64130) );
  XNOR2X1 U42041 ( .A(n64064), .B(n64413), .Y(n40815) );
  NOR2X1 U42042 ( .A(n40817), .B(n40816), .Y(n48967) );
  INVX1 U42043 ( .A(n57672), .Y(n40816) );
  NOR2X1 U42044 ( .A(n48966), .B(n42194), .Y(n40817) );
  NOR2X1 U42045 ( .A(n40818), .B(n40819), .Y(n57795) );
  INVX1 U42046 ( .A(n57793), .Y(n40818) );
  NOR2X1 U42047 ( .A(n31289), .B(n42046), .Y(n40819) );
  NOR2X1 U42048 ( .A(n40820), .B(n42196), .Y(n31654) );
  INVX1 U42049 ( .A(n57677), .Y(n40820) );
  XOR2X1 U42050 ( .A(n59881), .B(n40821), .Y(n59875) );
  XNOR2X1 U42051 ( .A(n59879), .B(n59677), .Y(n40821) );
  NAND2X1 U42052 ( .A(n38493), .B(n39853), .Y(n63824) );
  XOR2X1 U42053 ( .A(n59679), .B(n40822), .Y(n59691) );
  XNOR2X1 U42054 ( .A(n59230), .B(n59229), .Y(n40822) );
  XOR2X1 U42055 ( .A(n60617), .B(n40823), .Y(n60631) );
  XNOR2X1 U42056 ( .A(n60618), .B(n60245), .Y(n40823) );
  NAND2X1 U42057 ( .A(n63821), .B(n36781), .Y(n45291) );
  OR2X1 U42058 ( .A(n40824), .B(n42798), .Y(n62895) );
  NOR2X1 U42059 ( .A(n61178), .B(n61177), .Y(n40824) );
  XNOR2X1 U42060 ( .A(n40825), .B(n50027), .Y(n50229) );
  XNOR2X1 U42061 ( .A(n44057), .B(n44636), .Y(n40825) );
  XOR2X1 U42062 ( .A(n50169), .B(n40826), .Y(n50170) );
  XNOR2X1 U42063 ( .A(n50168), .B(n50167), .Y(n40826) );
  XOR2X1 U42064 ( .A(n50152), .B(n40827), .Y(n50153) );
  XNOR2X1 U42065 ( .A(n50151), .B(n50150), .Y(n40827) );
  XOR2X1 U42066 ( .A(n50312), .B(n40828), .Y(n50313) );
  XNOR2X1 U42067 ( .A(n50311), .B(n50310), .Y(n40828) );
  XOR2X1 U42068 ( .A(n54972), .B(n40829), .Y(n54973) );
  XNOR2X1 U42069 ( .A(n54971), .B(n54970), .Y(n40829) );
  NAND2X1 U42070 ( .A(n40830), .B(n40831), .Y(n46894) );
  NOR2X1 U42071 ( .A(n46854), .B(n46853), .Y(n40830) );
  NAND2X1 U42072 ( .A(n40490), .B(n46893), .Y(n40831) );
  NAND2X1 U42073 ( .A(n49627), .B(n49626), .Y(n49628) );
  NOR2X1 U42074 ( .A(n47342), .B(n40832), .Y(n47343) );
  INVX1 U42075 ( .A(n42334), .Y(n40832) );
  NAND2X1 U42076 ( .A(n49586), .B(n49585), .Y(n40833) );
  NAND2X1 U42077 ( .A(n49598), .B(n49597), .Y(n40834) );
  OR2X1 U42078 ( .A(n39195), .B(n40870), .Y(n49593) );
  NAND2X1 U42079 ( .A(n40835), .B(n40836), .Y(n61187) );
  NOR2X1 U42080 ( .A(n45218), .B(n45217), .Y(n40835) );
  NOR2X1 U42081 ( .A(n45249), .B(n45248), .Y(n40836) );
  NAND2X1 U42082 ( .A(n40837), .B(n40838), .Y(n51965) );
  NAND2X1 U42083 ( .A(n50038), .B(n50037), .Y(n40837) );
  NAND2X1 U42084 ( .A(n50041), .B(n50040), .Y(n40838) );
  NAND2X1 U42085 ( .A(n40839), .B(n40840), .Y(n54438) );
  NAND2X1 U42086 ( .A(n43307), .B(n54431), .Y(n40839) );
  NAND2X1 U42087 ( .A(n43312), .B(n54432), .Y(n40840) );
  NOR2X1 U42088 ( .A(n40842), .B(n45292), .Y(n40841) );
  INVX1 U42089 ( .A(n36237), .Y(n40842) );
  AND2X1 U42090 ( .A(n29623), .B(n40935), .Y(n40843) );
  AND2X1 U42091 ( .A(n46787), .B(n42878), .Y(n40844) );
  AND2X1 U42092 ( .A(n46657), .B(n42877), .Y(n40845) );
  NOR2X1 U42093 ( .A(n40846), .B(n40847), .Y(n46725) );
  NAND2X1 U42094 ( .A(n40499), .B(n40035), .Y(n40847) );
  NAND2X1 U42095 ( .A(n44982), .B(n38919), .Y(n58820) );
  NOR2X1 U42096 ( .A(n40848), .B(n40849), .Y(n47294) );
  NOR2X1 U42097 ( .A(n39354), .B(n37153), .Y(n40848) );
  NOR2X1 U42098 ( .A(n43092), .B(n40360), .Y(n40849) );
  NOR2X1 U42099 ( .A(n40850), .B(n40851), .Y(n45656) );
  NOR2X1 U42100 ( .A(n40852), .B(n40853), .Y(n45652) );
  NAND2X1 U42101 ( .A(n42785), .B(n36665), .Y(n40853) );
  NOR2X1 U42102 ( .A(n47303), .B(n36748), .Y(n47305) );
  NOR2X1 U42103 ( .A(n40854), .B(n42911), .Y(n46586) );
  NAND2X1 U42104 ( .A(n40499), .B(n46736), .Y(n40855) );
  NOR2X1 U42105 ( .A(n40856), .B(n45507), .Y(n46544) );
  NOR2X1 U42106 ( .A(n40858), .B(n42911), .Y(n46407) );
  NOR2X1 U42107 ( .A(n40859), .B(n40860), .Y(n46052) );
  OR2X1 U42108 ( .A(n40508), .B(n42693), .Y(n40860) );
  NOR2X1 U42109 ( .A(n40861), .B(n40862), .Y(n46378) );
  NAND2X1 U42110 ( .A(n42146), .B(n40404), .Y(n40862) );
  NOR2X1 U42111 ( .A(n40863), .B(n40864), .Y(n47677) );
  NAND2X1 U42112 ( .A(n48199), .B(n42673), .Y(n40864) );
  NOR2X1 U42113 ( .A(n40865), .B(n40866), .Y(n45498) );
  NAND2X1 U42114 ( .A(n42749), .B(n42760), .Y(n40866) );
  NOR2X1 U42115 ( .A(n40867), .B(n40868), .Y(n46061) );
  OR2X1 U42116 ( .A(n42694), .B(n42867), .Y(n40868) );
  NOR2X1 U42117 ( .A(n40869), .B(n42866), .Y(n45494) );
  NAND2X1 U42118 ( .A(n40454), .B(n42749), .Y(n40870) );
  NOR2X1 U42119 ( .A(n40871), .B(n40872), .Y(n47680) );
  NAND2X1 U42120 ( .A(n39810), .B(n43019), .Y(n40872) );
  NOR2X1 U42121 ( .A(n40873), .B(n40874), .Y(n46976) );
  NOR2X1 U42122 ( .A(n39354), .B(n37155), .Y(n40873) );
  NOR2X1 U42123 ( .A(n40360), .B(n43154), .Y(n40874) );
  NOR2X1 U42124 ( .A(n40875), .B(n40876), .Y(n45242) );
  NAND2X1 U42125 ( .A(n46216), .B(n36665), .Y(n40876) );
  NOR2X1 U42126 ( .A(n40877), .B(n40878), .Y(n45193) );
  NAND2X1 U42127 ( .A(n46049), .B(n38947), .Y(n40878) );
  NOR2X1 U42128 ( .A(n40879), .B(n40880), .Y(n47659) );
  NAND2X1 U42129 ( .A(n48199), .B(n58130), .Y(n40880) );
  NOR2X1 U42130 ( .A(n40881), .B(n40882), .Y(n48359) );
  NAND2X1 U42131 ( .A(n40448), .B(n43017), .Y(n40882) );
  NOR2X1 U42132 ( .A(n40883), .B(n40896), .Y(n45740) );
  NOR2X1 U42133 ( .A(n40884), .B(n45870), .Y(n45196) );
  NOR2X1 U42134 ( .A(n40885), .B(n40886), .Y(n45284) );
  NAND2X1 U42135 ( .A(n51983), .B(n46216), .Y(n40886) );
  NOR2X1 U42136 ( .A(n40887), .B(n40888), .Y(n45646) );
  NAND2X1 U42137 ( .A(n42697), .B(n42771), .Y(n40888) );
  NOR2X1 U42138 ( .A(n40889), .B(n40890), .Y(n46036) );
  OR2X1 U42139 ( .A(n45632), .B(n39195), .Y(n40890) );
  NOR2X1 U42140 ( .A(n40891), .B(n40892), .Y(n46035) );
  OR2X1 U42141 ( .A(n42866), .B(n39196), .Y(n40892) );
  NOR2X1 U42142 ( .A(n40893), .B(n40894), .Y(n47645) );
  NAND2X1 U42143 ( .A(n48205), .B(n58130), .Y(n40894) );
  NOR2X1 U42144 ( .A(n40895), .B(n40896), .Y(n45641) );
  NAND2X1 U42145 ( .A(n39198), .B(n42771), .Y(n40896) );
  NOR2X1 U42146 ( .A(n40897), .B(n40898), .Y(n45283) );
  NAND2X1 U42147 ( .A(n38537), .B(n46054), .Y(n40898) );
  NOR2X1 U42148 ( .A(n40899), .B(n40900), .Y(n46042) );
  OR2X1 U42149 ( .A(n45200), .B(n42693), .Y(n40900) );
  NOR2X1 U42150 ( .A(n40901), .B(n40902), .Y(n48387) );
  NAND2X1 U42151 ( .A(n42742), .B(n42673), .Y(n40902) );
  NOR2X1 U42152 ( .A(n40903), .B(n46030), .Y(n46187) );
  NOR2X1 U42153 ( .A(n40904), .B(n40905), .Y(n46041) );
  OR2X1 U42154 ( .A(n42764), .B(n40534), .Y(n40905) );
  NOR2X1 U42155 ( .A(n40906), .B(n40907), .Y(n45192) );
  NAND2X1 U42156 ( .A(n42699), .B(n42774), .Y(n40907) );
  NOR2X1 U42157 ( .A(n40908), .B(n40909), .Y(n45229) );
  NAND2X1 U42158 ( .A(n39197), .B(n42771), .Y(n40909) );
  AND2X1 U42159 ( .A(n40910), .B(n40911), .Y(n42515) );
  NAND2X1 U42160 ( .A(writeback_exec_value_w[4]), .B(n43026), .Y(n40910) );
  NAND2X1 U42161 ( .A(n38271), .B(n48452), .Y(n40911) );
  AND2X1 U42162 ( .A(n40912), .B(n40453), .Y(n42516) );
  NOR2X1 U42163 ( .A(n39115), .B(n36599), .Y(n40912) );
  NAND2X1 U42164 ( .A(n40913), .B(n40914), .Y(mem_i_pc_o[2]) );
  NOR2X1 U42165 ( .A(n54433), .B(n54438), .Y(n40913) );
  OR2X1 U42166 ( .A(n1760), .B(n42846), .Y(n40914) );
  NOR2X1 U42167 ( .A(n40915), .B(n40916), .Y(n50037) );
  NOR2X1 U42168 ( .A(opcode_instr_w_24), .B(n50033), .Y(n40915) );
  NOR2X1 U42169 ( .A(n50036), .B(n50040), .Y(n40916) );
  NOR2X1 U42170 ( .A(opcode_instr_w[12]), .B(n40917), .Y(n50661) );
  NAND2X1 U42171 ( .A(n40918), .B(n40919), .Y(n56824) );
  NOR2X1 U42172 ( .A(n54897), .B(n50669), .Y(n40918) );
  NOR2X1 U42173 ( .A(n40920), .B(n40921), .Y(n44971) );
  NOR2X1 U42174 ( .A(n43032), .B(n40249), .Y(n40920) );
  OR2X1 U42175 ( .A(n1852), .B(n40922), .Y(n27964) );
  OR2X1 U42176 ( .A(opcode_instr_w_45), .B(n29634), .Y(n40922) );
  AND2X1 U42177 ( .A(n40923), .B(u_csr_csr_mie_q_1), .Y(n29607) );
  OR2X1 U42178 ( .A(n40924), .B(u_muldiv_q_mask_q[7]), .Y(n29546) );
  OR2X1 U42179 ( .A(u_muldiv_q_mask_q[9]), .B(u_muldiv_q_mask_q[8]), .Y(n40924) );
  OR2X1 U42180 ( .A(n40925), .B(opcode_instr_w_46), .Y(n24367) );
  AND2X1 U42181 ( .A(n40926), .B(n40927), .Y(n29538) );
  NOR2X1 U42182 ( .A(u_muldiv_q_mask_q[25]), .B(u_muldiv_q_mask_q[26]), .Y(
        n40926) );
  NOR2X1 U42183 ( .A(u_muldiv_q_mask_q[23]), .B(u_muldiv_q_mask_q[24]), .Y(
        n40927) );
  AND2X1 U42184 ( .A(n40928), .B(n40929), .Y(n29539) );
  NOR2X1 U42185 ( .A(u_muldiv_q_mask_q[29]), .B(u_muldiv_q_mask_q[2]), .Y(
        n40928) );
  NOR2X1 U42186 ( .A(u_muldiv_q_mask_q[27]), .B(u_muldiv_q_mask_q[28]), .Y(
        n40929) );
  AND2X1 U42187 ( .A(n43013), .B(n40930), .Y(n42579) );
  AND2X1 U42188 ( .A(n50858), .B(n40931), .Y(n42609) );
  NOR2X1 U42189 ( .A(n8810), .B(n40932), .Y(n28550) );
  NOR2X1 U42190 ( .A(n1887), .B(n40933), .Y(n28551) );
  NAND2X1 U42191 ( .A(opcode_instr_w[5]), .B(n40934), .Y(n58539) );
  AND2X1 U42192 ( .A(n34489), .B(n35891), .Y(n40935) );
  OR2X1 U42193 ( .A(n40936), .B(mem_d_resp_tag_i[4]), .Y(n45025) );
  OR2X1 U42194 ( .A(mem_d_resp_tag_i[0]), .B(n45297), .Y(n40936) );
  AND2X1 U42195 ( .A(n36248), .B(n45163), .Y(n40937) );
  AND2X1 U42196 ( .A(n36163), .B(n73527), .Y(n40938) );
  AND2X1 U42197 ( .A(n46094), .B(n42876), .Y(n40939) );
  AND2X1 U42198 ( .A(n45382), .B(n42877), .Y(n40940) );
  AND2X1 U42199 ( .A(n46245), .B(n42877), .Y(n40941) );
  AND2X1 U42200 ( .A(n42876), .B(n45273), .Y(n40942) );
  INVX1 U42201 ( .A(n42615), .Y(n40943) );
  XOR2X1 U42202 ( .A(n40168), .B(n67935), .Y(n67947) );
  XOR2X1 U42203 ( .A(n71733), .B(n39412), .Y(n72677) );
  XNOR2X1 U42204 ( .A(n70524), .B(n70827), .Y(n70508) );
  AND2X1 U42205 ( .A(n61027), .B(n61026), .Y(n40945) );
  XOR2X1 U42206 ( .A(n71178), .B(n71185), .Y(n71181) );
  XOR2X1 U42207 ( .A(n38619), .B(n40948), .Y(n40946) );
  XOR2X1 U42208 ( .A(n70144), .B(n39153), .Y(n70145) );
  AND2X1 U42209 ( .A(n64996), .B(n64812), .Y(n40947) );
  AND2X1 U42210 ( .A(n63583), .B(n63851), .Y(n40948) );
  XNOR2X1 U42211 ( .A(n67052), .B(n67076), .Y(n67055) );
  OR2X1 U42212 ( .A(n69282), .B(n40949), .Y(n69258) );
  INVX1 U42213 ( .A(n69198), .Y(n40949) );
  XOR2X1 U42214 ( .A(n69601), .B(n69597), .Y(n70453) );
  NAND2X1 U42215 ( .A(n71153), .B(n40950), .Y(n71435) );
  AND2X1 U42216 ( .A(n71154), .B(n71152), .Y(n40950) );
  XOR2X1 U42217 ( .A(n71114), .B(n71115), .Y(n71116) );
  AND2X1 U42218 ( .A(n39952), .B(n67982), .Y(n40951) );
  XOR2X1 U42219 ( .A(n72097), .B(n38399), .Y(n72666) );
  XNOR2X1 U42220 ( .A(n71699), .B(n71698), .Y(n40952) );
  XNOR2X1 U42221 ( .A(n66936), .B(n66937), .Y(n66938) );
  AND2X1 U42222 ( .A(n67294), .B(n67291), .Y(n40953) );
  XOR2X1 U42223 ( .A(n67287), .B(n40953), .Y(n67290) );
  XNOR2X1 U42224 ( .A(n69248), .B(n68819), .Y(n68820) );
  AND2X1 U42225 ( .A(n40949), .B(n69192), .Y(n40954) );
  XOR2X1 U42226 ( .A(n71163), .B(n71162), .Y(n40955) );
  AND2X1 U42227 ( .A(n38160), .B(n70776), .Y(n40956) );
  AND2X1 U42228 ( .A(n37377), .B(n60263), .Y(n40957) );
  XNOR2X1 U42229 ( .A(n68830), .B(n68829), .Y(n69543) );
  NAND2X1 U42230 ( .A(n68884), .B(n40958), .Y(n68825) );
  AND2X1 U42231 ( .A(n68885), .B(n68886), .Y(n40958) );
  AND2X1 U42232 ( .A(n69529), .B(n69528), .Y(n40959) );
  XNOR2X1 U42233 ( .A(n67255), .B(n67256), .Y(n67264) );
  AND2X1 U42234 ( .A(n62884), .B(n62883), .Y(n40960) );
  AND2X1 U42235 ( .A(n67939), .B(n40961), .Y(n67941) );
  OR2X1 U42236 ( .A(n40962), .B(n67940), .Y(n40961) );
  AND2X1 U42237 ( .A(n39760), .B(n67581), .Y(n40962) );
  AND2X1 U42238 ( .A(n40963), .B(n69267), .Y(n69265) );
  INVX1 U42239 ( .A(n69264), .Y(n40963) );
  OR2X1 U42240 ( .A(n40964), .B(n67940), .Y(n67586) );
  OR2X1 U42241 ( .A(n40962), .B(n67582), .Y(n40964) );
  XNOR2X1 U42242 ( .A(n67625), .B(n67618), .Y(n67620) );
  XNOR2X1 U42243 ( .A(n71414), .B(n40965), .Y(n71405) );
  XNOR2X1 U42244 ( .A(n72101), .B(n71404), .Y(n40965) );
  XNOR2X1 U42245 ( .A(n70765), .B(n40966), .Y(n71115) );
  XNOR2X1 U42246 ( .A(n71173), .B(n70764), .Y(n40966) );
  XNOR2X1 U42247 ( .A(n67575), .B(n67576), .Y(n67642) );
  XOR2X1 U42248 ( .A(n68549), .B(n41072), .Y(n68551) );
  NAND2X1 U42249 ( .A(n71762), .B(n40967), .Y(n71782) );
  AND2X1 U42250 ( .A(n71764), .B(n71763), .Y(n40967) );
  AND2X1 U42251 ( .A(n68872), .B(n40968), .Y(n68874) );
  AND2X1 U42252 ( .A(n41060), .B(n68873), .Y(n40968) );
  XNOR2X1 U42253 ( .A(n66529), .B(n66530), .Y(n66536) );
  XOR2X1 U42254 ( .A(n63008), .B(n62392), .Y(n62396) );
  XOR2X1 U42255 ( .A(n69875), .B(n69536), .Y(n69538) );
  XOR2X1 U42256 ( .A(n41128), .B(n66896), .Y(n40969) );
  AND2X1 U42257 ( .A(n67953), .B(n40970), .Y(n68210) );
  AND2X1 U42258 ( .A(n67954), .B(n67955), .Y(n40970) );
  XOR2X1 U42259 ( .A(n70775), .B(n70528), .Y(n70827) );
  XNOR2X1 U42260 ( .A(n69588), .B(n69534), .Y(n69535) );
  XOR2X1 U42261 ( .A(n41105), .B(n41108), .Y(n40971) );
  XNOR2X1 U42262 ( .A(n67231), .B(n67232), .Y(n67247) );
  XNOR2X1 U42263 ( .A(n70478), .B(n40972), .Y(n70178) );
  XNOR2X1 U42264 ( .A(n71402), .B(n70212), .Y(n40972) );
  AND2X1 U42265 ( .A(n64451), .B(n65025), .Y(n40973) );
  AND2X1 U42266 ( .A(n64451), .B(n40974), .Y(n65028) );
  XNOR2X1 U42267 ( .A(n68241), .B(n40975), .Y(n68516) );
  XOR2X1 U42268 ( .A(n68249), .B(n70762), .Y(n40975) );
  AND2X1 U42269 ( .A(n65100), .B(n65101), .Y(n65102) );
  XOR2X1 U42270 ( .A(n64454), .B(n65010), .Y(n64811) );
  XNOR2X1 U42271 ( .A(n71187), .B(n40977), .Y(n40976) );
  XOR2X1 U42272 ( .A(n70760), .B(n70885), .Y(n40977) );
  AND2X1 U42273 ( .A(n66175), .B(n66176), .Y(n40978) );
  XNOR2X1 U42274 ( .A(n65966), .B(n65960), .Y(n65963) );
  AND2X1 U42275 ( .A(n70120), .B(n70220), .Y(n40979) );
  XOR2X1 U42276 ( .A(n41104), .B(n70442), .Y(n70446) );
  OR2X1 U42277 ( .A(n68454), .B(n68453), .Y(n40980) );
  AND2X1 U42278 ( .A(n66175), .B(n66177), .Y(n40981) );
  AND2X1 U42279 ( .A(n68544), .B(n68545), .Y(n68547) );
  NOR2X1 U42280 ( .A(n38062), .B(n69571), .Y(n40982) );
  OR2X1 U42281 ( .A(n40990), .B(n64391), .Y(n40983) );
  XNOR2X1 U42282 ( .A(n66682), .B(n66322), .Y(n66438) );
  AND2X1 U42283 ( .A(n64207), .B(n64208), .Y(n64210) );
  XOR2X1 U42284 ( .A(n64721), .B(n40973), .Y(n65019) );
  XOR2X1 U42285 ( .A(n36657), .B(n41171), .Y(n40984) );
  XNOR2X1 U42286 ( .A(n65009), .B(n65035), .Y(n40985) );
  AND2X1 U42287 ( .A(n70549), .B(n70548), .Y(n40986) );
  NAND2X1 U42288 ( .A(n65715), .B(n40987), .Y(n65714) );
  AND2X1 U42289 ( .A(n65716), .B(n65717), .Y(n40987) );
  AND2X1 U42290 ( .A(n63580), .B(n63581), .Y(n40988) );
  NAND2X1 U42291 ( .A(n67019), .B(n40989), .Y(n67328) );
  AND2X1 U42292 ( .A(n67021), .B(n67020), .Y(n40989) );
  XOR2X1 U42293 ( .A(n71212), .B(n71204), .Y(n71208) );
  XOR2X1 U42294 ( .A(n41193), .B(n70576), .Y(n70564) );
  XNOR2X1 U42295 ( .A(n65363), .B(n65367), .Y(n65370) );
  AND2X1 U42296 ( .A(n64384), .B(n64383), .Y(n40990) );
  AND2X1 U42297 ( .A(n63794), .B(n63795), .Y(n40991) );
  AND2X1 U42298 ( .A(n63580), .B(n63582), .Y(n40992) );
  XOR2X1 U42299 ( .A(n66680), .B(n39968), .Y(n66686) );
  XOR2X1 U42300 ( .A(n71198), .B(n71206), .Y(n71199) );
  XOR2X1 U42301 ( .A(n66417), .B(n66093), .Y(n66098) );
  AND2X1 U42302 ( .A(n68969), .B(n40993), .Y(n68972) );
  OR2X1 U42303 ( .A(n38986), .B(n68971), .Y(n40993) );
  AND2X1 U42304 ( .A(n66785), .B(n66784), .Y(n40994) );
  XOR2X1 U42305 ( .A(n71442), .B(n71445), .Y(n71446) );
  XOR2X1 U42306 ( .A(n68086), .B(n67783), .Y(n68419) );
  XNOR2X1 U42307 ( .A(n72077), .B(n40995), .Y(n72082) );
  XOR2X1 U42308 ( .A(n72081), .B(n72080), .Y(n40995) );
  XOR2X1 U42309 ( .A(n68428), .B(n68427), .Y(n68710) );
  XNOR2X1 U42310 ( .A(n65031), .B(n65088), .Y(n65036) );
  XOR2X1 U42311 ( .A(n64727), .B(n40996), .Y(n65026) );
  AND2X1 U42312 ( .A(n64751), .B(n64750), .Y(n40996) );
  OR2X1 U42313 ( .A(n67441), .B(n40997), .Y(n67076) );
  AND2X1 U42314 ( .A(n66716), .B(n67077), .Y(n40997) );
  AND2X1 U42315 ( .A(n65436), .B(n65435), .Y(n40998) );
  XOR2X1 U42316 ( .A(n39102), .B(n65804), .Y(n40999) );
  XNOR2X1 U42317 ( .A(n67712), .B(n67705), .Y(n67709) );
  AND2X1 U42318 ( .A(n65729), .B(n65736), .Y(n41000) );
  AND2X1 U42319 ( .A(n67725), .B(n67436), .Y(n41001) );
  XNOR2X1 U42320 ( .A(n68084), .B(n68085), .Y(n68324) );
  XNOR2X1 U42321 ( .A(n65552), .B(n41002), .Y(n65201) );
  XNOR2X1 U42322 ( .A(n65553), .B(n71402), .Y(n41002) );
  AND2X1 U42323 ( .A(n68132), .B(n68131), .Y(n41003) );
  AND2X1 U42324 ( .A(n69388), .B(n69052), .Y(n41004) );
  AND2X1 U42325 ( .A(n68350), .B(n69055), .Y(n41005) );
  XOR2X1 U42326 ( .A(n66742), .B(n67090), .Y(n66394) );
  NOR2X1 U42327 ( .A(n67771), .B(n67772), .Y(n41006) );
  XNOR2X1 U42328 ( .A(n68088), .B(n68383), .Y(n68339) );
  XOR2X1 U42329 ( .A(n70327), .B(n70330), .Y(n70336) );
  OR2X1 U42330 ( .A(n41007), .B(n38368), .Y(n66964) );
  OR2X1 U42331 ( .A(n39929), .B(n39300), .Y(n41007) );
  OR2X1 U42332 ( .A(n41008), .B(n41009), .Y(n67650) );
  AND2X1 U42333 ( .A(n43536), .B(n67569), .Y(n41008) );
  AND2X1 U42334 ( .A(n43536), .B(n67646), .Y(n41009) );
  AND2X1 U42335 ( .A(n70214), .B(n70837), .Y(n41010) );
  XNOR2X1 U42336 ( .A(n69934), .B(n41011), .Y(n69877) );
  XNOR2X1 U42337 ( .A(n39858), .B(n69862), .Y(n41011) );
  AND2X1 U42338 ( .A(n68594), .B(n41012), .Y(n68592) );
  INVX1 U42339 ( .A(n43560), .Y(n41012) );
  AND2X1 U42340 ( .A(n40235), .B(n43559), .Y(n41013) );
  NOR2X1 U42341 ( .A(n41015), .B(n41016), .Y(n41014) );
  OR2X1 U42342 ( .A(n71421), .B(n72102), .Y(n41015) );
  AND2X1 U42343 ( .A(n71422), .B(n72098), .Y(n41016) );
  XOR2X1 U42344 ( .A(n72105), .B(n41014), .Y(n72646) );
  XOR2X1 U42345 ( .A(n69513), .B(n69514), .Y(n69524) );
  AND2X1 U42346 ( .A(n69926), .B(n69871), .Y(n41017) );
  AND2X1 U42347 ( .A(n71142), .B(n71141), .Y(n41018) );
  AND2X1 U42348 ( .A(n70507), .B(n71152), .Y(n41020) );
  OR2X1 U42349 ( .A(n59438), .B(n59510), .Y(n59439) );
  OR2X1 U42350 ( .A(n43528), .B(n70780), .Y(n70840) );
  XOR2X1 U42351 ( .A(n71430), .B(n71149), .Y(n71706) );
  OR2X1 U42352 ( .A(n41021), .B(n41022), .Y(n68903) );
  AND2X1 U42353 ( .A(n68565), .B(n68564), .Y(n41021) );
  AND2X1 U42354 ( .A(n68569), .B(n68910), .Y(n41022) );
  AND2X1 U42355 ( .A(n67283), .B(n41024), .Y(n67286) );
  AND2X1 U42356 ( .A(n67285), .B(n67284), .Y(n41024) );
  XNOR2X1 U42357 ( .A(n67980), .B(n41026), .Y(n68572) );
  XNOR2X1 U42358 ( .A(n67983), .B(n67979), .Y(n41026) );
  NOR2X1 U42359 ( .A(n36570), .B(n40561), .Y(n41027) );
  OR2X1 U42360 ( .A(n41029), .B(n40395), .Y(n72715) );
  OR2X1 U42361 ( .A(n36569), .B(n41273), .Y(n41029) );
  OR2X1 U42362 ( .A(n68515), .B(n41031), .Y(n68884) );
  OR2X1 U42363 ( .A(n39888), .B(n68517), .Y(n41031) );
  XOR2X1 U42364 ( .A(n66506), .B(n65884), .Y(n66224) );
  AND2X1 U42365 ( .A(n66225), .B(n39851), .Y(n41032) );
  AND2X1 U42366 ( .A(n69889), .B(n69890), .Y(n41033) );
  XNOR2X1 U42367 ( .A(n36752), .B(n69537), .Y(n69244) );
  XNOR2X1 U42368 ( .A(n67623), .B(n67624), .Y(n67886) );
  XOR2X1 U42369 ( .A(n67217), .B(n67218), .Y(n67219) );
  AND2X1 U42370 ( .A(n68911), .B(n68910), .Y(n41034) );
  XNOR2X1 U42371 ( .A(n40421), .B(n67983), .Y(n67990) );
  AND2X1 U42372 ( .A(n71158), .B(n70842), .Y(n41035) );
  AND2X1 U42373 ( .A(n68212), .B(n68237), .Y(n41036) );
  XOR2X1 U42374 ( .A(n72098), .B(n71713), .Y(n72106) );
  XOR2X1 U42375 ( .A(n65287), .B(n65480), .Y(n41037) );
  OR2X1 U42376 ( .A(n61128), .B(n41038), .Y(n62412) );
  AND2X1 U42377 ( .A(n38508), .B(n36755), .Y(n41038) );
  AND2X1 U42378 ( .A(n39423), .B(n38981), .Y(n63001) );
  XOR2X1 U42379 ( .A(n39362), .B(n41039), .Y(n70478) );
  XOR2X1 U42380 ( .A(n69884), .B(n43654), .Y(n41039) );
  XNOR2X1 U42381 ( .A(n70477), .B(n41040), .Y(n70504) );
  XOR2X1 U42382 ( .A(n70478), .B(n43524), .Y(n41040) );
  OR2X1 U42383 ( .A(n38930), .B(n41041), .Y(n71169) );
  AND2X1 U42384 ( .A(n70765), .B(n71106), .Y(n41041) );
  NOR2X1 U42385 ( .A(n41043), .B(n41044), .Y(n41042) );
  AND2X1 U42386 ( .A(n43642), .B(n70461), .Y(n41043) );
  AND2X1 U42387 ( .A(n43642), .B(n70466), .Y(n41044) );
  OR2X1 U42388 ( .A(n43669), .B(n66597), .Y(n67223) );
  AND2X1 U42389 ( .A(n67275), .B(n67274), .Y(n41045) );
  AND2X1 U42390 ( .A(n69921), .B(n70467), .Y(n41046) );
  AND2X1 U42391 ( .A(n43521), .B(n71696), .Y(n41047) );
  OR2X1 U42392 ( .A(n71173), .B(n41048), .Y(n70847) );
  AND2X1 U42393 ( .A(n43642), .B(n70846), .Y(n41048) );
  AND2X1 U42394 ( .A(n69528), .B(n69529), .Y(n68907) );
  XOR2X1 U42395 ( .A(n43546), .B(n67961), .Y(n67963) );
  AND2X1 U42396 ( .A(n67203), .B(n67209), .Y(n41049) );
  OR2X1 U42397 ( .A(n41050), .B(n41051), .Y(n67884) );
  AND2X1 U42398 ( .A(n40142), .B(n67267), .Y(n41050) );
  AND2X1 U42399 ( .A(n67271), .B(n67270), .Y(n41051) );
  XOR2X1 U42400 ( .A(n69861), .B(n66605), .Y(n66527) );
  XNOR2X1 U42401 ( .A(n67222), .B(n66587), .Y(n66588) );
  AND2X1 U42402 ( .A(n43545), .B(n66517), .Y(n41052) );
  XNOR2X1 U42403 ( .A(n59926), .B(n41053), .Y(n59932) );
  OR2X1 U42404 ( .A(n59734), .B(n59733), .Y(n41053) );
  XOR2X1 U42405 ( .A(n69918), .B(n69589), .Y(n69596) );
  NOR2X1 U42406 ( .A(n41055), .B(n41056), .Y(n41054) );
  AND2X1 U42407 ( .A(n43677), .B(n69545), .Y(n41055) );
  AND2X1 U42408 ( .A(n69549), .B(n68865), .Y(n41056) );
  AND2X1 U42409 ( .A(n67965), .B(n67966), .Y(n41057) );
  XOR2X1 U42410 ( .A(n68858), .B(n68857), .Y(n69546) );
  XOR2X1 U42411 ( .A(n41058), .B(n67228), .Y(n67585) );
  OR2X1 U42412 ( .A(n67268), .B(n41316), .Y(n41058) );
  AND2X1 U42413 ( .A(n67616), .B(n67617), .Y(n41059) );
  AND2X1 U42414 ( .A(n68824), .B(n68823), .Y(n41060) );
  AND2X1 U42415 ( .A(n62489), .B(n62491), .Y(n41061) );
  XNOR2X1 U42416 ( .A(n66931), .B(n41062), .Y(n66929) );
  XNOR2X1 U42417 ( .A(n66932), .B(n66893), .Y(n41062) );
  XNOR2X1 U42418 ( .A(n65177), .B(n65178), .Y(n65180) );
  XOR2X1 U42419 ( .A(n66932), .B(n66934), .Y(n66935) );
  XOR2X1 U42420 ( .A(n69605), .B(n41063), .Y(n69597) );
  XNOR2X1 U42421 ( .A(n69940), .B(n69512), .Y(n41063) );
  AND2X1 U42422 ( .A(n67274), .B(n67275), .Y(n41064) );
  AND2X1 U42423 ( .A(n66267), .B(n66266), .Y(n66270) );
  XNOR2X1 U42424 ( .A(n67884), .B(n41065), .Y(n67626) );
  XNOR2X1 U42425 ( .A(n67624), .B(n67580), .Y(n41065) );
  NAND2X1 U42426 ( .A(n67283), .B(n41066), .Y(n67862) );
  AND2X1 U42427 ( .A(n67284), .B(n67285), .Y(n41066) );
  XOR2X1 U42428 ( .A(n68803), .B(n68802), .Y(n68809) );
  XNOR2X1 U42429 ( .A(n41067), .B(n36694), .Y(n67655) );
  OR2X1 U42430 ( .A(n66948), .B(n66947), .Y(n41067) );
  XNOR2X1 U42431 ( .A(n70826), .B(n70823), .Y(n71104) );
  AND2X1 U42432 ( .A(n66272), .B(n66598), .Y(n41068) );
  XNOR2X1 U42433 ( .A(n41299), .B(n41069), .Y(n72101) );
  XNOR2X1 U42434 ( .A(n71698), .B(n71403), .Y(n41069) );
  AND2X1 U42435 ( .A(n72110), .B(n36565), .Y(n41070) );
  XOR2X1 U42436 ( .A(n66512), .B(n66513), .Y(n66526) );
  XOR2X1 U42437 ( .A(n66617), .B(n66613), .Y(n66614) );
  XOR2X1 U42438 ( .A(n68825), .B(n68826), .Y(n68873) );
  OR2X1 U42439 ( .A(n66494), .B(n39171), .Y(n66873) );
  XOR2X1 U42440 ( .A(n66513), .B(n66216), .Y(n41071) );
  AND2X1 U42441 ( .A(n68559), .B(n68558), .Y(n41072) );
  XOR2X1 U42442 ( .A(n68880), .B(n68881), .Y(n68891) );
  AND2X1 U42443 ( .A(n39725), .B(n71688), .Y(n41073) );
  XOR2X1 U42444 ( .A(n68511), .B(n68553), .Y(n68512) );
  XOR2X1 U42445 ( .A(n63152), .B(n63154), .Y(n63162) );
  XOR2X1 U42446 ( .A(n68505), .B(n68506), .Y(n68570) );
  OR2X1 U42447 ( .A(n39320), .B(n65904), .Y(n65179) );
  AND2X1 U42448 ( .A(n65193), .B(n65541), .Y(n41074) );
  NAND2X1 U42449 ( .A(n68005), .B(n41075), .Y(n68196) );
  AND2X1 U42450 ( .A(n68008), .B(n68004), .Y(n41075) );
  XOR2X1 U42451 ( .A(n66928), .B(n66894), .Y(n66926) );
  XNOR2X1 U42452 ( .A(n70534), .B(n70526), .Y(n70527) );
  XNOR2X1 U42453 ( .A(n66257), .B(n66258), .Y(n41076) );
  OR2X1 U42454 ( .A(n41077), .B(n70470), .Y(n70776) );
  OR2X1 U42455 ( .A(n70469), .B(n70468), .Y(n41077) );
  AND2X1 U42456 ( .A(n65246), .B(n65900), .Y(n41078) );
  NOR2X1 U42457 ( .A(n43668), .B(n64873), .Y(n41079) );
  AND2X1 U42458 ( .A(n41080), .B(n67639), .Y(n67870) );
  OR2X1 U42459 ( .A(n67577), .B(n67640), .Y(n41080) );
  XOR2X1 U42460 ( .A(n69245), .B(n69216), .Y(n69551) );
  AND2X1 U42461 ( .A(n70181), .B(n43505), .Y(n41081) );
  AND2X1 U42462 ( .A(n66589), .B(n41082), .Y(n66591) );
  INVX1 U42463 ( .A(n41335), .Y(n41082) );
  XOR2X1 U42464 ( .A(n68815), .B(n68893), .Y(n68816) );
  NAND2X1 U42465 ( .A(n62877), .B(n41083), .Y(n62880) );
  AND2X1 U42466 ( .A(n62879), .B(n62878), .Y(n41083) );
  XNOR2X1 U42467 ( .A(n70465), .B(n41084), .Y(n70471) );
  XNOR2X1 U42468 ( .A(n70459), .B(n70156), .Y(n41084) );
  XNOR2X1 U42469 ( .A(n65910), .B(n65911), .Y(n65915) );
  OR2X1 U42470 ( .A(n43647), .B(n68211), .Y(n68239) );
  AND2X1 U42471 ( .A(n62489), .B(n62490), .Y(n41085) );
  XNOR2X1 U42472 ( .A(n62428), .B(n41086), .Y(n62490) );
  OR2X1 U42473 ( .A(n61214), .B(n61213), .Y(n41086) );
  OR2X1 U42474 ( .A(n41087), .B(n69255), .Y(n69584) );
  AND2X1 U42475 ( .A(n69249), .B(n69250), .Y(n41087) );
  AND2X1 U42476 ( .A(n67293), .B(n41088), .Y(n67628) );
  OR2X1 U42477 ( .A(n67297), .B(n67296), .Y(n41088) );
  XOR2X1 U42478 ( .A(n67931), .B(n67930), .Y(n67932) );
  AND2X1 U42479 ( .A(n61007), .B(n61008), .Y(n61016) );
  AND2X1 U42480 ( .A(n70179), .B(n70178), .Y(n41089) );
  XOR2X1 U42481 ( .A(n67213), .B(n67212), .Y(n67214) );
  XOR2X1 U42482 ( .A(n67860), .B(n67573), .Y(n67638) );
  XOR2X1 U42483 ( .A(n38524), .B(n63762), .Y(n63763) );
  AND2X1 U42484 ( .A(n40382), .B(n64843), .Y(n41090) );
  XNOR2X1 U42485 ( .A(n71176), .B(n41091), .Y(n71161) );
  XNOR2X1 U42486 ( .A(n71182), .B(n71103), .Y(n41091) );
  XOR2X1 U42487 ( .A(n67198), .B(n67199), .Y(n67200) );
  OR2X1 U42488 ( .A(n41092), .B(n72102), .Y(n72103) );
  OR2X1 U42489 ( .A(n43691), .B(n72101), .Y(n41092) );
  XOR2X1 U42490 ( .A(n66581), .B(n66582), .Y(n66583) );
  XNOR2X1 U42491 ( .A(n41093), .B(n70521), .Y(n70523) );
  AND2X1 U42492 ( .A(n70770), .B(n70771), .Y(n41093) );
  AND2X1 U42493 ( .A(n67893), .B(n67892), .Y(n41094) );
  AND2X1 U42494 ( .A(n68861), .B(n68860), .Y(n41095) );
  XNOR2X1 U42495 ( .A(n68487), .B(n41097), .Y(n68007) );
  XNOR2X1 U42496 ( .A(n68464), .B(n67846), .Y(n41097) );
  AND2X1 U42497 ( .A(n43664), .B(n65192), .Y(n41098) );
  XOR2X1 U42498 ( .A(n43692), .B(n41099), .Y(n70795) );
  AND2X1 U42499 ( .A(n70793), .B(n70816), .Y(n41099) );
  XNOR2X1 U42500 ( .A(n70845), .B(n41100), .Y(n70823) );
  XNOR2X1 U42501 ( .A(n70851), .B(n70763), .Y(n41100) );
  XOR2X1 U42502 ( .A(n67658), .B(n66939), .Y(n67567) );
  AND2X1 U42503 ( .A(n70445), .B(n70444), .Y(n41101) );
  XOR2X1 U42504 ( .A(n68566), .B(n68206), .Y(n68242) );
  XNOR2X1 U42505 ( .A(n63178), .B(n41102), .Y(n63268) );
  XNOR2X1 U42506 ( .A(n40241), .B(n63175), .Y(n41102) );
  XNOR2X1 U42507 ( .A(n63268), .B(n41103), .Y(n63283) );
  XNOR2X1 U42508 ( .A(n63269), .B(n63264), .Y(n41103) );
  XOR2X1 U42509 ( .A(n65875), .B(n41427), .Y(n65881) );
  XOR2X1 U42510 ( .A(n68793), .B(n68794), .Y(n69178) );
  AND2X1 U42511 ( .A(n65924), .B(n65925), .Y(n41105) );
  NOR2X1 U42512 ( .A(n43530), .B(n66540), .Y(n41106) );
  AND2X1 U42513 ( .A(n65968), .B(n66259), .Y(n41107) );
  XOR2X1 U42514 ( .A(n60661), .B(n60660), .Y(n60672) );
  XOR2X1 U42515 ( .A(n43644), .B(n65546), .Y(n41108) );
  AND2X1 U42516 ( .A(n65548), .B(n65920), .Y(n41109) );
  AND2X1 U42517 ( .A(n43677), .B(n67247), .Y(n41110) );
  AND2X1 U42518 ( .A(n64051), .B(n64052), .Y(n41111) );
  AND2X1 U42519 ( .A(n67667), .B(n67666), .Y(n41112) );
  XNOR2X1 U42520 ( .A(n68597), .B(n41113), .Y(n68794) );
  XOR2X1 U42521 ( .A(n68785), .B(n70272), .Y(n41113) );
  XOR2X1 U42522 ( .A(n70215), .B(n38192), .Y(n70217) );
  XOR2X1 U42523 ( .A(n63582), .B(n41114), .Y(n63515) );
  XNOR2X1 U42524 ( .A(n63579), .B(n63581), .Y(n41114) );
  XNOR2X1 U42525 ( .A(n68907), .B(n68894), .Y(n69255) );
  AND2X1 U42526 ( .A(n43677), .B(n67891), .Y(n41115) );
  AND2X1 U42527 ( .A(n41392), .B(n71755), .Y(n41116) );
  AND2X1 U42528 ( .A(n68967), .B(n69477), .Y(n41117) );
  XOR2X1 U42529 ( .A(n67706), .B(n67464), .Y(n67702) );
  XOR2X1 U42530 ( .A(n68978), .B(n68970), .Y(n41118) );
  AND2X1 U42531 ( .A(n67000), .B(n66999), .Y(n41119) );
  XOR2X1 U42532 ( .A(n68022), .B(n40027), .Y(n68477) );
  AND2X1 U42533 ( .A(n63332), .B(n63331), .Y(n41120) );
  XNOR2X1 U42534 ( .A(n41121), .B(n66318), .Y(n66314) );
  XOR2X1 U42535 ( .A(n66819), .B(n66820), .Y(n41121) );
  AND2X1 U42536 ( .A(n65706), .B(n65705), .Y(n41122) );
  XOR2X1 U42537 ( .A(n66173), .B(n66463), .Y(n66319) );
  AND2X1 U42538 ( .A(n66083), .B(n66082), .Y(n41123) );
  XOR2X1 U42539 ( .A(n64526), .B(n64874), .Y(n64881) );
  XNOR2X1 U42540 ( .A(n68858), .B(n41125), .Y(n41124) );
  XOR2X1 U42541 ( .A(n68857), .B(n43679), .Y(n41125) );
  XOR2X1 U42542 ( .A(n66258), .B(n66229), .Y(n41126) );
  XNOR2X1 U42543 ( .A(n66177), .B(n65827), .Y(n66197) );
  AND2X1 U42544 ( .A(n66673), .B(n67140), .Y(n41127) );
  XOR2X1 U42545 ( .A(n66582), .B(n66538), .Y(n41128) );
  XOR2X1 U42546 ( .A(n64833), .B(n65119), .Y(n65138) );
  AND2X1 U42547 ( .A(n71087), .B(n71088), .Y(n41129) );
  XOR2X1 U42548 ( .A(n64147), .B(n64146), .Y(n64155) );
  AND2X1 U42549 ( .A(n65486), .B(n65159), .Y(n41130) );
  OR2X1 U42550 ( .A(n36775), .B(n69598), .Y(n69940) );
  AND2X1 U42551 ( .A(n65139), .B(n41131), .Y(n65137) );
  INVX1 U42552 ( .A(n65135), .Y(n41131) );
  AND2X1 U42553 ( .A(n64370), .B(n65124), .Y(n41132) );
  XNOR2X1 U42554 ( .A(n64173), .B(n41133), .Y(n64184) );
  OR2X1 U42555 ( .A(n63861), .B(n63860), .Y(n41133) );
  AND2X1 U42556 ( .A(n69171), .B(n69170), .Y(n41134) );
  XOR2X1 U42557 ( .A(n69858), .B(n70118), .Y(n70136) );
  XNOR2X1 U42558 ( .A(n70756), .B(n70554), .Y(n70557) );
  OR2X1 U42559 ( .A(n70218), .B(n41135), .Y(n70233) );
  AND2X1 U42560 ( .A(n70133), .B(n70135), .Y(n41135) );
  XNOR2X1 U42561 ( .A(n39521), .B(n68959), .Y(n68960) );
  XNOR2X1 U42562 ( .A(n71439), .B(n41136), .Y(n71787) );
  XNOR2X1 U42563 ( .A(n71660), .B(n71438), .Y(n41136) );
  AND2X1 U42564 ( .A(n66895), .B(n66899), .Y(n41137) );
  AND2X1 U42565 ( .A(n68870), .B(n68869), .Y(n41138) );
  XNOR2X1 U42566 ( .A(n41139), .B(n68520), .Y(n68842) );
  AND2X1 U42567 ( .A(n68835), .B(n68834), .Y(n41139) );
  NAND2X1 U42568 ( .A(n71128), .B(n41140), .Y(n70818) );
  OR2X1 U42569 ( .A(n70204), .B(n71133), .Y(n41140) );
  XNOR2X1 U42570 ( .A(n71691), .B(n41141), .Y(n71752) );
  XNOR2X1 U42571 ( .A(n38561), .B(n71689), .Y(n41141) );
  AND2X1 U42572 ( .A(n72137), .B(n72136), .Y(n41142) );
  AND2X1 U42573 ( .A(n70118), .B(n39958), .Y(n41143) );
  XNOR2X1 U42574 ( .A(n41144), .B(n69897), .Y(n70190) );
  AND2X1 U42575 ( .A(n70205), .B(n70206), .Y(n41144) );
  AND2X1 U42576 ( .A(n64845), .B(n64843), .Y(n41145) );
  AND2X1 U42577 ( .A(n67015), .B(n67017), .Y(n41146) );
  AND2X1 U42578 ( .A(n68280), .B(n68782), .Y(n41147) );
  XNOR2X1 U42579 ( .A(n65138), .B(n41148), .Y(n66180) );
  XNOR2X1 U42580 ( .A(n65139), .B(n65135), .Y(n41148) );
  AND2X1 U42581 ( .A(n70119), .B(n70118), .Y(n41149) );
  XNOR2X1 U42582 ( .A(n41150), .B(n66163), .Y(n66177) );
  XOR2X1 U42583 ( .A(n66162), .B(n66171), .Y(n41150) );
  NAND2X1 U42584 ( .A(n64451), .B(n41151), .Y(n64734) );
  AND2X1 U42585 ( .A(n65026), .B(n64733), .Y(n41151) );
  XOR2X1 U42586 ( .A(n38179), .B(n69164), .Y(n69295) );
  XOR2X1 U42587 ( .A(n38047), .B(n69550), .Y(n41152) );
  XOR2X1 U42588 ( .A(n43644), .B(n64914), .Y(n41153) );
  XOR2X1 U42589 ( .A(n65197), .B(n64883), .Y(n64908) );
  AND2X1 U42590 ( .A(n64295), .B(n64294), .Y(n41154) );
  AND2X1 U42591 ( .A(n67029), .B(n67030), .Y(n41155) );
  AND2X1 U42592 ( .A(n64368), .B(n64367), .Y(n41156) );
  NAND2X1 U42593 ( .A(n67812), .B(n41157), .Y(n67825) );
  AND2X1 U42594 ( .A(n67807), .B(n67809), .Y(n41157) );
  AND2X1 U42595 ( .A(n64912), .B(n64911), .Y(n41158) );
  OR2X1 U42596 ( .A(n41159), .B(n41160), .Y(n69220) );
  OR2X1 U42597 ( .A(n41204), .B(n37994), .Y(n41159) );
  AND2X1 U42598 ( .A(n43505), .B(n68838), .Y(n41160) );
  OR2X1 U42599 ( .A(n41161), .B(n41162), .Y(n68839) );
  OR2X1 U42600 ( .A(n41416), .B(n67921), .Y(n41161) );
  AND2X1 U42601 ( .A(n67923), .B(n67924), .Y(n41162) );
  AND2X1 U42602 ( .A(n43507), .B(n67898), .Y(n41163) );
  AND2X1 U42603 ( .A(n68548), .B(n69231), .Y(n41164) );
  XNOR2X1 U42604 ( .A(n67357), .B(n67028), .Y(n41165) );
  XNOR2X1 U42605 ( .A(n66086), .B(n41166), .Y(n66089) );
  OR2X1 U42606 ( .A(n66345), .B(n66344), .Y(n41166) );
  XNOR2X1 U42607 ( .A(n67980), .B(n67859), .Y(n67962) );
  OR2X1 U42608 ( .A(n41167), .B(n68607), .Y(n68608) );
  OR2X1 U42609 ( .A(n43593), .B(n68933), .Y(n41167) );
  XOR2X1 U42610 ( .A(n67897), .B(n41168), .Y(n67925) );
  OR2X1 U42611 ( .A(n41115), .B(n67896), .Y(n41168) );
  XOR2X1 U42612 ( .A(n72084), .B(n71767), .Y(n71791) );
  OR2X1 U42613 ( .A(n65369), .B(n41169), .Y(n65726) );
  AND2X1 U42614 ( .A(n65372), .B(n65371), .Y(n41169) );
  OR2X1 U42615 ( .A(n41170), .B(n67508), .Y(n67510) );
  AND2X1 U42616 ( .A(n67169), .B(n67168), .Y(n41170) );
  XNOR2X1 U42617 ( .A(n41172), .B(n65713), .Y(n41171) );
  XOR2X1 U42618 ( .A(n65723), .B(n65720), .Y(n41172) );
  OR2X1 U42619 ( .A(n65014), .B(n41173), .Y(n65371) );
  AND2X1 U42620 ( .A(n65022), .B(n65021), .Y(n41173) );
  AND2X1 U42621 ( .A(n61011), .B(n41174), .Y(n61014) );
  AND2X1 U42622 ( .A(n61013), .B(n61012), .Y(n41174) );
  XNOR2X1 U42623 ( .A(n64823), .B(n64824), .Y(n65338) );
  AND2X1 U42624 ( .A(n66196), .B(n66197), .Y(n41175) );
  AND2X1 U42625 ( .A(n64381), .B(n64380), .Y(n41176) );
  XNOR2X1 U42626 ( .A(n65603), .B(n41177), .Y(n65596) );
  XOR2X1 U42627 ( .A(n65602), .B(n43524), .Y(n41177) );
  AND2X1 U42628 ( .A(n67015), .B(n67016), .Y(n41178) );
  XNOR2X1 U42629 ( .A(n63521), .B(n41179), .Y(n63582) );
  XNOR2X1 U42630 ( .A(n63524), .B(n63525), .Y(n41179) );
  AND2X1 U42631 ( .A(n68856), .B(n43705), .Y(n41180) );
  XOR2X1 U42632 ( .A(n64709), .B(n65105), .Y(n64710) );
  XNOR2X1 U42633 ( .A(n65368), .B(n41181), .Y(n65360) );
  XNOR2X1 U42634 ( .A(n65739), .B(n65097), .Y(n41181) );
  XOR2X1 U42635 ( .A(n70818), .B(n70493), .Y(n70500) );
  AND2X1 U42636 ( .A(n69292), .B(n69291), .Y(n41182) );
  XOR2X1 U42637 ( .A(n70219), .B(n40979), .Y(n70537) );
  OR2X1 U42638 ( .A(n70097), .B(n41183), .Y(n69822) );
  OR2X1 U42639 ( .A(n43618), .B(n39306), .Y(n41183) );
  AND2X1 U42640 ( .A(n43655), .B(n65196), .Y(n41184) );
  XNOR2X1 U42641 ( .A(n39281), .B(n41186), .Y(n41185) );
  XOR2X1 U42642 ( .A(n65460), .B(n65840), .Y(n41186) );
  AND2X1 U42643 ( .A(n67811), .B(n67808), .Y(n41187) );
  XOR2X1 U42644 ( .A(n64373), .B(n41423), .Y(n41188) );
  XOR2X1 U42645 ( .A(n40984), .B(n65675), .Y(n65676) );
  AND2X1 U42646 ( .A(n63515), .B(n63516), .Y(n41189) );
  AND2X1 U42647 ( .A(n63517), .B(n63515), .Y(n41190) );
  AND2X1 U42648 ( .A(n43676), .B(n65557), .Y(n41191) );
  XNOR2X1 U42649 ( .A(n68759), .B(n41192), .Y(n68456) );
  XNOR2X1 U42650 ( .A(n39570), .B(n68455), .Y(n41192) );
  XNOR2X1 U42651 ( .A(n70436), .B(n41194), .Y(n41193) );
  XOR2X1 U42652 ( .A(n70435), .B(n70434), .Y(n41194) );
  XOR2X1 U42653 ( .A(n69232), .B(n69898), .Y(n69241) );
  XNOR2X1 U42654 ( .A(n68165), .B(n41195), .Y(n68079) );
  XNOR2X1 U42655 ( .A(n68082), .B(n68076), .Y(n41195) );
  AND2X1 U42656 ( .A(n67141), .B(n67140), .Y(n41196) );
  AND2X1 U42657 ( .A(n43706), .B(n69572), .Y(n41197) );
  AND2X1 U42658 ( .A(n63510), .B(n63511), .Y(n41198) );
  XOR2X1 U42659 ( .A(n65723), .B(n65713), .Y(n65719) );
  XOR2X1 U42660 ( .A(n64447), .B(n41199), .Y(n64173) );
  XNOR2X1 U42661 ( .A(n64147), .B(n63850), .Y(n41199) );
  XOR2X1 U42662 ( .A(n67594), .B(n67899), .Y(n67613) );
  XNOR2X1 U42663 ( .A(n71096), .B(n41200), .Y(n71204) );
  XNOR2X1 U42664 ( .A(n71211), .B(n71095), .Y(n41200) );
  OR2X1 U42665 ( .A(n70129), .B(n41201), .Y(n69619) );
  OR2X1 U42666 ( .A(n43536), .B(n69618), .Y(n41201) );
  AND2X1 U42667 ( .A(n63510), .B(n63512), .Y(n41202) );
  XOR2X1 U42668 ( .A(n70889), .B(n70439), .Y(n70440) );
  AND2X1 U42669 ( .A(n67035), .B(n66689), .Y(n41203) );
  XOR2X1 U42670 ( .A(n68615), .B(n39025), .Y(n68705) );
  AND2X1 U42671 ( .A(n43506), .B(n67925), .Y(n41204) );
  AND2X1 U42672 ( .A(n66463), .B(n66462), .Y(n41205) );
  NAND2X1 U42673 ( .A(n68419), .B(n37365), .Y(n68083) );
  XOR2X1 U42674 ( .A(n69432), .B(n69140), .Y(n69438) );
  OR2X1 U42675 ( .A(n67054), .B(n41206), .Y(n67456) );
  AND2X1 U42676 ( .A(n67071), .B(n67070), .Y(n41206) );
  AND2X1 U42677 ( .A(n68161), .B(n68160), .Y(n41207) );
  XOR2X1 U42678 ( .A(n67327), .B(n67473), .Y(n67338) );
  AND2X1 U42679 ( .A(n67332), .B(n41208), .Y(n67335) );
  OR2X1 U42680 ( .A(n67334), .B(n67333), .Y(n41208) );
  AND2X1 U42681 ( .A(n41518), .B(n66462), .Y(n41209) );
  OR2X1 U42682 ( .A(n67789), .B(n67796), .Y(n68172) );
  XOR2X1 U42683 ( .A(n69653), .B(n69677), .Y(n69953) );
  XNOR2X1 U42684 ( .A(n70570), .B(n41210), .Y(n70571) );
  XOR2X1 U42685 ( .A(n70569), .B(n70582), .Y(n41210) );
  XOR2X1 U42686 ( .A(n68223), .B(n36516), .Y(n68529) );
  XOR2X1 U42687 ( .A(n64907), .B(n64887), .Y(n64905) );
  XOR2X1 U42688 ( .A(n36402), .B(n67903), .Y(n67915) );
  XNOR2X1 U42689 ( .A(n63804), .B(n41211), .Y(n63794) );
  XNOR2X1 U42690 ( .A(n64165), .B(n63791), .Y(n41211) );
  XNOR2X1 U42691 ( .A(n41212), .B(n66902), .Y(n66922) );
  AND2X1 U42692 ( .A(n67248), .B(n67249), .Y(n41212) );
  XNOR2X1 U42693 ( .A(n71668), .B(n41213), .Y(n71670) );
  XNOR2X1 U42694 ( .A(n71667), .B(n71666), .Y(n41213) );
  XNOR2X1 U42695 ( .A(n72076), .B(n41214), .Y(n72611) );
  XNOR2X1 U42696 ( .A(n72595), .B(n72075), .Y(n41214) );
  AND2X1 U42697 ( .A(n72173), .B(n41215), .Y(n72063) );
  AND2X1 U42698 ( .A(n72174), .B(n72065), .Y(n41215) );
  XNOR2X1 U42699 ( .A(n38047), .B(n66580), .Y(n41216) );
  AND2X1 U42700 ( .A(n66256), .B(n66578), .Y(n41217) );
  XOR2X1 U42701 ( .A(n66570), .B(n66545), .Y(n66567) );
  XOR2X1 U42702 ( .A(n40324), .B(n65952), .Y(n41218) );
  XOR2X1 U42703 ( .A(n66252), .B(n66236), .Y(n66548) );
  AND2X1 U42704 ( .A(n38224), .B(n66112), .Y(n41220) );
  XNOR2X1 U42705 ( .A(n65086), .B(n65087), .Y(n41221) );
  XOR2X1 U42706 ( .A(n72039), .B(n72054), .Y(n72040) );
  XOR2X1 U42707 ( .A(n66254), .B(n66235), .Y(n66251) );
  AND2X1 U42708 ( .A(n65589), .B(n65590), .Y(n41222) );
  XOR2X1 U42709 ( .A(n64541), .B(n64269), .Y(n64582) );
  XOR2X1 U42710 ( .A(n66919), .B(n66905), .Y(n66917) );
  XNOR2X1 U42711 ( .A(n72039), .B(n41223), .Y(n72079) );
  OR2X1 U42712 ( .A(n71658), .B(n71657), .Y(n41223) );
  XOR2X1 U42713 ( .A(n72627), .B(n72612), .Y(n72615) );
  AND2X1 U42714 ( .A(n65441), .B(n65795), .Y(n41224) );
  AND2X1 U42715 ( .A(n41225), .B(n72562), .Y(n72073) );
  AND2X1 U42716 ( .A(n38169), .B(n43620), .Y(n41225) );
  NOR2X1 U42717 ( .A(n43702), .B(n65205), .Y(n41226) );
  XOR2X1 U42718 ( .A(n64904), .B(n64888), .Y(n65203) );
  XOR2X1 U42719 ( .A(n41485), .B(n69417), .Y(n69433) );
  XNOR2X1 U42720 ( .A(n66703), .B(n66701), .Y(n66690) );
  XOR2X1 U42721 ( .A(n66403), .B(n66101), .Y(n66357) );
  XOR2X1 U42722 ( .A(n72611), .B(n72610), .Y(n72629) );
  NOR2X1 U42723 ( .A(n41228), .B(n66770), .Y(n41227) );
  INVX1 U42724 ( .A(n67073), .Y(n41228) );
  AND2X1 U42725 ( .A(n64273), .B(n64272), .Y(n41229) );
  AND2X1 U42726 ( .A(n65219), .B(n65220), .Y(n65222) );
  XNOR2X1 U42727 ( .A(n64578), .B(n41230), .Y(n64891) );
  XOR2X1 U42728 ( .A(n64577), .B(n43508), .Y(n41230) );
  AND2X1 U42729 ( .A(n65413), .B(n41231), .Y(n65415) );
  OR2X1 U42730 ( .A(n65428), .B(n65414), .Y(n41231) );
  XNOR2X1 U42731 ( .A(n65088), .B(n41232), .Y(n65009) );
  XOR2X1 U42732 ( .A(n65031), .B(n65023), .Y(n41232) );
  AND2X1 U42733 ( .A(n65588), .B(n41233), .Y(n65591) );
  AND2X1 U42734 ( .A(n65589), .B(n65590), .Y(n41233) );
  XNOR2X1 U42735 ( .A(n66546), .B(n41234), .Y(n66554) );
  XOR2X1 U42736 ( .A(n66548), .B(n43693), .Y(n41234) );
  XNOR2X1 U42737 ( .A(n63698), .B(n41235), .Y(n63938) );
  XOR2X1 U42738 ( .A(n63697), .B(n37975), .Y(n41235) );
  XOR2X1 U42739 ( .A(n41236), .B(n68394), .Y(n68683) );
  XOR2X1 U42740 ( .A(n68395), .B(n41521), .Y(n41236) );
  AND2X1 U42741 ( .A(n41237), .B(n68136), .Y(n68137) );
  OR2X1 U42742 ( .A(n68135), .B(n68134), .Y(n41237) );
  XOR2X1 U42743 ( .A(n65788), .B(n66115), .Y(n66400) );
  AND2X1 U42744 ( .A(n72037), .B(n72036), .Y(n41238) );
  AND2X1 U42745 ( .A(n65568), .B(n65569), .Y(n65572) );
  XOR2X1 U42746 ( .A(n64894), .B(n65206), .Y(n64903) );
  XOR2X1 U42747 ( .A(n41004), .B(n69138), .Y(n41239) );
  AND2X1 U42748 ( .A(n66760), .B(n67384), .Y(n41240) );
  AND2X1 U42749 ( .A(n43544), .B(n72595), .Y(n41241) );
  XOR2X1 U42750 ( .A(n69053), .B(n69011), .Y(n69050) );
  AND2X1 U42751 ( .A(n66750), .B(n41242), .Y(n66759) );
  AND2X1 U42752 ( .A(n67110), .B(n66751), .Y(n41242) );
  XOR2X1 U42753 ( .A(n69037), .B(n68680), .Y(n69003) );
  XNOR2X1 U42754 ( .A(n64555), .B(n41243), .Y(n64560) );
  XOR2X1 U42755 ( .A(n64554), .B(n43693), .Y(n41243) );
  XOR2X1 U42756 ( .A(n66378), .B(n66718), .Y(n67090) );
  XNOR2X1 U42757 ( .A(n69706), .B(n41244), .Y(n69786) );
  XNOR2X1 U42758 ( .A(n69697), .B(n69707), .Y(n41244) );
  AND2X1 U42759 ( .A(n69385), .B(n69698), .Y(n41245) );
  XNOR2X1 U42760 ( .A(n69385), .B(n41247), .Y(n41246) );
  XOR2X1 U42761 ( .A(n69698), .B(n69699), .Y(n41247) );
  XOR2X1 U42762 ( .A(n67106), .B(n67396), .Y(n41248) );
  OR2X1 U42763 ( .A(n67407), .B(n41249), .Y(n67100) );
  AND2X1 U42764 ( .A(n67097), .B(n67096), .Y(n41249) );
  XOR2X1 U42765 ( .A(n67101), .B(n68113), .Y(n67402) );
  NOR2X1 U42766 ( .A(n41251), .B(n69057), .Y(n41250) );
  INVX1 U42767 ( .A(n68634), .Y(n41251) );
  OR2X1 U42768 ( .A(n69716), .B(n69715), .Y(n69368) );
  OR2X1 U42769 ( .A(n41252), .B(n68119), .Y(n68114) );
  AND2X1 U42770 ( .A(n67760), .B(n67759), .Y(n41252) );
  XOR2X1 U42771 ( .A(n72188), .B(n72164), .Y(n72167) );
  XOR2X1 U42772 ( .A(n41506), .B(n62409), .Y(n41253) );
  XOR2X1 U42773 ( .A(n71550), .B(n71551), .Y(n41254) );
  OR2X1 U42774 ( .A(n41255), .B(n41256), .Y(n66479) );
  AND2X1 U42775 ( .A(n66477), .B(n66476), .Y(n41255) );
  AND2X1 U42776 ( .A(n66478), .B(n44017), .Y(n41256) );
  OR2X1 U42777 ( .A(n59436), .B(n59364), .Y(n59365) );
  AND2X1 U42778 ( .A(n65858), .B(n66018), .Y(n41257) );
  AND2X1 U42779 ( .A(n64026), .B(n64027), .Y(n41258) );
  NOR2X1 U42780 ( .A(n41260), .B(n41261), .Y(n41259) );
  OR2X1 U42781 ( .A(n39769), .B(n62861), .Y(n41260) );
  AND2X1 U42782 ( .A(n62862), .B(n63141), .Y(n41261) );
  XOR2X1 U42783 ( .A(n59728), .B(n59724), .Y(n59277) );
  XOR2X1 U42784 ( .A(n41262), .B(n38684), .Y(n61120) );
  XOR2X1 U42785 ( .A(n61234), .B(n61233), .Y(n41262) );
  OR2X1 U42786 ( .A(n41263), .B(n41264), .Y(n59859) );
  AND2X1 U42787 ( .A(n59856), .B(n60061), .Y(n41263) );
  AND2X1 U42788 ( .A(n60057), .B(n59858), .Y(n41264) );
  AND2X1 U42789 ( .A(n63919), .B(n63453), .Y(n41265) );
  XOR2X1 U42790 ( .A(n61295), .B(n61104), .Y(n61116) );
  NOR2X1 U42791 ( .A(n41267), .B(n40481), .Y(n41266) );
  OR2X1 U42792 ( .A(n69917), .B(n43650), .Y(n41267) );
  XNOR2X1 U42793 ( .A(n66504), .B(n66505), .Y(n66507) );
  AND2X1 U42794 ( .A(n61289), .B(n61290), .Y(n61292) );
  NOR2X1 U42795 ( .A(n41269), .B(n41270), .Y(n41268) );
  AND2X1 U42796 ( .A(n62535), .B(n62536), .Y(n41269) );
  AND2X1 U42797 ( .A(n62539), .B(n62538), .Y(n41270) );
  XNOR2X1 U42798 ( .A(n61263), .B(n41271), .Y(n61267) );
  OR2X1 U42799 ( .A(n61262), .B(n61261), .Y(n41271) );
  OR2X1 U42800 ( .A(n59714), .B(n59713), .Y(n59718) );
  XOR2X1 U42801 ( .A(n65151), .B(n65667), .Y(n65478) );
  AND2X1 U42802 ( .A(n66205), .B(n66206), .Y(n41272) );
  NAND2X1 U42803 ( .A(n39044), .B(n59378), .Y(n59310) );
  AND2X1 U42804 ( .A(n71126), .B(n40456), .Y(n41273) );
  OR2X1 U42805 ( .A(n69244), .B(n41274), .Y(n69246) );
  INVX1 U42806 ( .A(n43529), .Y(n41274) );
  AND2X1 U42807 ( .A(n60915), .B(n60914), .Y(n41275) );
  AND2X1 U42808 ( .A(n66207), .B(n66205), .Y(n41276) );
  XNOR2X1 U42809 ( .A(n65479), .B(n41277), .Y(n65287) );
  XOR2X1 U42810 ( .A(n65152), .B(n65655), .Y(n41277) );
  AND2X1 U42811 ( .A(n60994), .B(n60993), .Y(n41278) );
  XNOR2X1 U42812 ( .A(n59705), .B(n41279), .Y(n59714) );
  OR2X1 U42813 ( .A(n59263), .B(n59262), .Y(n41279) );
  AND2X1 U42814 ( .A(n64356), .B(n41280), .Y(n64352) );
  INVX1 U42815 ( .A(n64351), .Y(n41280) );
  XOR2X1 U42816 ( .A(n64842), .B(n64844), .Y(n64484) );
  AND2X1 U42817 ( .A(n70491), .B(n70490), .Y(n41281) );
  XNOR2X1 U42818 ( .A(n60998), .B(n41282), .Y(n61003) );
  OR2X1 U42819 ( .A(n60657), .B(n60656), .Y(n41282) );
  AND2X1 U42820 ( .A(n37319), .B(n65481), .Y(n41283) );
  OR2X1 U42821 ( .A(n64321), .B(n64322), .Y(n64323) );
  XOR2X1 U42822 ( .A(n41284), .B(n63366), .Y(n63650) );
  OR2X1 U42823 ( .A(n63151), .B(n63150), .Y(n41284) );
  AND2X1 U42824 ( .A(n66604), .B(n41285), .Y(n66596) );
  AND2X1 U42825 ( .A(n66277), .B(n66600), .Y(n41285) );
  OR2X1 U42826 ( .A(n60260), .B(n41286), .Y(n61007) );
  AND2X1 U42827 ( .A(n63353), .B(n63356), .Y(n41287) );
  XNOR2X1 U42828 ( .A(n68198), .B(n41288), .Y(n68265) );
  XNOR2X1 U42829 ( .A(n68197), .B(n40317), .Y(n41288) );
  XNOR2X1 U42830 ( .A(n67856), .B(n41289), .Y(n67663) );
  XOR2X1 U42831 ( .A(n67855), .B(n43588), .Y(n41289) );
  AND2X1 U42832 ( .A(n64027), .B(n64028), .Y(n41290) );
  XOR2X1 U42833 ( .A(n65861), .B(n65860), .Y(n41291) );
  XNOR2X1 U42834 ( .A(n64638), .B(n41292), .Y(n64636) );
  XOR2X1 U42835 ( .A(n64504), .B(n64503), .Y(n41292) );
  OR2X1 U42836 ( .A(n61062), .B(n41293), .Y(n60703) );
  INVX1 U42837 ( .A(n61067), .Y(n41293) );
  OR2X1 U42838 ( .A(n41294), .B(n41295), .Y(n68560) );
  OR2X1 U42839 ( .A(n68253), .B(n68252), .Y(n41294) );
  AND2X1 U42840 ( .A(n39470), .B(n68254), .Y(n41295) );
  OR2X1 U42841 ( .A(n43632), .B(n67970), .Y(n41296) );
  AND2X1 U42842 ( .A(n66931), .B(n41297), .Y(n67268) );
  OR2X1 U42843 ( .A(n66935), .B(n43650), .Y(n41297) );
  AND2X1 U42844 ( .A(n64241), .B(n64319), .Y(n41298) );
  AND2X1 U42845 ( .A(n71165), .B(n71697), .Y(n41299) );
  XOR2X1 U42846 ( .A(n36525), .B(n65885), .Y(n66517) );
  XOR2X1 U42847 ( .A(n67276), .B(n67216), .Y(n41300) );
  AND2X1 U42848 ( .A(n38048), .B(n43682), .Y(n41301) );
  AND2X1 U42849 ( .A(n66008), .B(n41291), .Y(n41302) );
  XNOR2X1 U42850 ( .A(n41303), .B(n61003), .Y(n61032) );
  XOR2X1 U42851 ( .A(n61006), .B(n61002), .Y(n41303) );
  OR2X1 U42852 ( .A(n41304), .B(n41305), .Y(n67965) );
  AND2X1 U42853 ( .A(n67871), .B(n43635), .Y(n41304) );
  AND2X1 U42854 ( .A(n67879), .B(n67878), .Y(n41305) );
  AND2X1 U42855 ( .A(n64957), .B(n64958), .Y(n41306) );
  OR2X1 U42856 ( .A(n71116), .B(n38047), .Y(n71434) );
  OR2X1 U42857 ( .A(n38047), .B(n69543), .Y(n68864) );
  AND2X1 U42858 ( .A(n70484), .B(n43682), .Y(n41307) );
  AND2X1 U42859 ( .A(n63731), .B(n63991), .Y(n41308) );
  INVX1 U42860 ( .A(n64511), .Y(n41309) );
  XOR2X1 U42861 ( .A(n63486), .B(n63328), .Y(n63603) );
  XNOR2X1 U42862 ( .A(n63594), .B(n41310), .Y(n63498) );
  XNOR2X1 U42863 ( .A(n63593), .B(n63590), .Y(n41310) );
  XNOR2X1 U42864 ( .A(n63493), .B(n41311), .Y(n63491) );
  XOR2X1 U42865 ( .A(n63498), .B(n63497), .Y(n41311) );
  AND2X1 U42866 ( .A(n59915), .B(n41312), .Y(n59910) );
  OR2X1 U42867 ( .A(n40399), .B(n60216), .Y(n41312) );
  XNOR2X1 U42868 ( .A(n65637), .B(n65638), .Y(n41313) );
  OR2X1 U42869 ( .A(n41314), .B(n41315), .Y(n67222) );
  AND2X1 U42870 ( .A(n66265), .B(n43673), .Y(n41314) );
  AND2X1 U42871 ( .A(n66270), .B(n66269), .Y(n41315) );
  AND2X1 U42872 ( .A(n66935), .B(n43648), .Y(n41316) );
  AND2X1 U42873 ( .A(n41317), .B(n68809), .Y(n68807) );
  INVX1 U42874 ( .A(n43540), .Y(n41317) );
  AND2X1 U42875 ( .A(n38212), .B(n41318), .Y(n66947) );
  AND2X1 U42876 ( .A(n67546), .B(n43587), .Y(n41318) );
  OR2X1 U42877 ( .A(n67545), .B(n41321), .Y(n66946) );
  AND2X1 U42878 ( .A(n66871), .B(n66872), .Y(n41321) );
  AND2X1 U42879 ( .A(n65882), .B(n65981), .Y(n41322) );
  XNOR2X1 U42880 ( .A(n68198), .B(n41323), .Y(n67983) );
  XNOR2X1 U42881 ( .A(n68197), .B(n67857), .Y(n41323) );
  AND2X1 U42882 ( .A(n66874), .B(n66494), .Y(n41324) );
  AND2X1 U42883 ( .A(n63012), .B(n63011), .Y(n41325) );
  AND2X1 U42884 ( .A(n63037), .B(n38295), .Y(n41326) );
  XNOR2X1 U42885 ( .A(n63765), .B(n41327), .Y(n64205) );
  XNOR2X1 U42886 ( .A(n63762), .B(n63596), .Y(n41327) );
  XOR2X1 U42887 ( .A(n65154), .B(n65155), .Y(n65490) );
  OR2X1 U42888 ( .A(n62520), .B(n62522), .Y(n61279) );
  AND2X1 U42889 ( .A(n59767), .B(n59766), .Y(n41328) );
  OR2X1 U42890 ( .A(n39186), .B(n69933), .Y(n69935) );
  NAND2X1 U42891 ( .A(n60292), .B(n41329), .Y(n60295) );
  AND2X1 U42892 ( .A(n60294), .B(n60293), .Y(n41329) );
  OR2X1 U42893 ( .A(n62344), .B(n41330), .Y(n62348) );
  XOR2X1 U42894 ( .A(n62347), .B(n62346), .Y(n41330) );
  AND2X1 U42895 ( .A(n64588), .B(n64587), .Y(n41331) );
  XNOR2X1 U42896 ( .A(n59714), .B(n41332), .Y(n59725) );
  OR2X1 U42897 ( .A(n59276), .B(n59275), .Y(n41332) );
  AND2X1 U42898 ( .A(n65260), .B(n41333), .Y(n65259) );
  AND2X1 U42899 ( .A(n65257), .B(n44049), .Y(n41333) );
  XOR2X1 U42900 ( .A(n66887), .B(n66511), .Y(n41334) );
  AND2X1 U42901 ( .A(n66536), .B(n43649), .Y(n41335) );
  OR2X1 U42902 ( .A(n60081), .B(n41336), .Y(n60059) );
  XOR2X1 U42903 ( .A(n60058), .B(n60057), .Y(n41336) );
  AND2X1 U42904 ( .A(n60571), .B(n60573), .Y(n41337) );
  NAND2X1 U42905 ( .A(n60170), .B(n41338), .Y(n60056) );
  AND2X1 U42906 ( .A(n60055), .B(n60054), .Y(n41338) );
  NOR2X1 U42907 ( .A(n70181), .B(n41417), .Y(n41339) );
  AND2X1 U42908 ( .A(n71698), .B(n43656), .Y(n41340) );
  AND2X1 U42909 ( .A(n67536), .B(n39292), .Y(n66975) );
  XOR2X1 U42910 ( .A(n59451), .B(n59453), .Y(n59455) );
  XNOR2X1 U42911 ( .A(n67212), .B(n41341), .Y(n67218) );
  XNOR2X1 U42912 ( .A(n43551), .B(n67213), .Y(n41341) );
  AND2X1 U42913 ( .A(n65263), .B(n65262), .Y(n41342) );
  XOR2X1 U42914 ( .A(n65247), .B(n41342), .Y(n65249) );
  OR2X1 U42915 ( .A(n63763), .B(n41343), .Y(n63766) );
  INVX1 U42916 ( .A(n63764), .Y(n41343) );
  XNOR2X1 U42917 ( .A(n63512), .B(n63299), .Y(n63507) );
  XNOR2X1 U42918 ( .A(n66180), .B(n41344), .Y(n64982) );
  XOR2X1 U42919 ( .A(n65845), .B(n66179), .Y(n41344) );
  XNOR2X1 U42920 ( .A(n70845), .B(n41345), .Y(n70846) );
  XNOR2X1 U42921 ( .A(n70850), .B(n70844), .Y(n41345) );
  XOR2X1 U42922 ( .A(n63890), .B(n64221), .Y(n64039) );
  NOR2X1 U42923 ( .A(n65542), .B(n43667), .Y(n41346) );
  XNOR2X1 U42924 ( .A(n39715), .B(n41348), .Y(n41347) );
  XOR2X1 U42925 ( .A(n66967), .B(n66210), .Y(n41348) );
  AND2X1 U42926 ( .A(n64976), .B(n64975), .Y(n41349) );
  AND2X1 U42927 ( .A(n68571), .B(n41350), .Y(n68916) );
  OR2X1 U42928 ( .A(n68574), .B(n68573), .Y(n41350) );
  INVX1 U42929 ( .A(n41457), .Y(n41351) );
  AND2X1 U42930 ( .A(n63470), .B(n63472), .Y(n41353) );
  AND2X1 U42931 ( .A(n66990), .B(n41354), .Y(n66993) );
  INVX1 U42932 ( .A(n66991), .Y(n41354) );
  XOR2X1 U42933 ( .A(n68193), .B(n68279), .Y(n68276) );
  OR2X1 U42934 ( .A(n41355), .B(n41356), .Y(n68861) );
  OR2X1 U42935 ( .A(n41115), .B(n68217), .Y(n41355) );
  AND2X1 U42936 ( .A(n41094), .B(n68218), .Y(n41356) );
  AND2X1 U42937 ( .A(n70517), .B(n41357), .Y(n70519) );
  AND2X1 U42938 ( .A(n70516), .B(n43668), .Y(n41357) );
  AND2X1 U42939 ( .A(n69586), .B(n43646), .Y(n41358) );
  AND2X1 U42940 ( .A(n60665), .B(n41359), .Y(n60264) );
  AND2X1 U42941 ( .A(n38378), .B(n42708), .Y(n41359) );
  AND2X1 U42942 ( .A(n63995), .B(n64001), .Y(n41360) );
  XNOR2X1 U42943 ( .A(n41361), .B(n62886), .Y(n63306) );
  XOR2X1 U42944 ( .A(n63290), .B(n63291), .Y(n41361) );
  XOR2X1 U42945 ( .A(n69934), .B(n69924), .Y(n70452) );
  XNOR2X1 U42946 ( .A(n41363), .B(n65638), .Y(n41362) );
  XOR2X1 U42947 ( .A(n65637), .B(n65639), .Y(n41363) );
  AND2X1 U42948 ( .A(n64587), .B(n64588), .Y(n64590) );
  XOR2X1 U42949 ( .A(n65280), .B(n65170), .Y(n65524) );
  XOR2X1 U42950 ( .A(n63866), .B(n63588), .Y(n63762) );
  AND2X1 U42951 ( .A(n70771), .B(n41364), .Y(n70773) );
  AND2X1 U42952 ( .A(n70770), .B(n43658), .Y(n41364) );
  AND2X1 U42953 ( .A(n64533), .B(n64532), .Y(n41365) );
  XNOR2X1 U42954 ( .A(n39297), .B(n68013), .Y(n68014) );
  XNOR2X1 U42955 ( .A(n63474), .B(n41367), .Y(n63462) );
  XNOR2X1 U42956 ( .A(n63369), .B(n63368), .Y(n41367) );
  XOR2X1 U42957 ( .A(n67540), .B(n39378), .Y(n67849) );
  XNOR2X1 U42958 ( .A(n41369), .B(n67889), .Y(n68219) );
  AND2X1 U42959 ( .A(n67622), .B(n67926), .Y(n41369) );
  XNOR2X1 U42960 ( .A(n41370), .B(n63516), .Y(n63512) );
  XOR2X1 U42961 ( .A(n63514), .B(n63515), .Y(n41370) );
  XOR2X1 U42962 ( .A(n63869), .B(n64198), .Y(n64052) );
  AND2X1 U42963 ( .A(n64873), .B(n43668), .Y(n41371) );
  AND2X1 U42964 ( .A(n64051), .B(n41709), .Y(n41372) );
  XNOR2X1 U42965 ( .A(n66219), .B(n41373), .Y(n65917) );
  XOR2X1 U42966 ( .A(n43636), .B(n65911), .Y(n41373) );
  OR2X1 U42967 ( .A(n67891), .B(n41374), .Y(n68218) );
  INVX1 U42968 ( .A(n43684), .Y(n41374) );
  AND2X1 U42969 ( .A(n38556), .B(n66179), .Y(n41375) );
  AND2X1 U42970 ( .A(n67317), .B(n67676), .Y(n41377) );
  AND2X1 U42971 ( .A(n67306), .B(n67305), .Y(n41378) );
  OR2X1 U42972 ( .A(n65724), .B(n41379), .Y(n66084) );
  NOR2X1 U42973 ( .A(n36773), .B(n65727), .Y(n41379) );
  XOR2X1 U42974 ( .A(n68439), .B(n68618), .Y(n68726) );
  XNOR2X1 U42975 ( .A(n70111), .B(n41380), .Y(n70116) );
  XOR2X1 U42976 ( .A(n69944), .B(n69943), .Y(n41380) );
  XOR2X1 U42977 ( .A(n70237), .B(n36604), .Y(n70240) );
  XNOR2X1 U42978 ( .A(n70861), .B(n41381), .Y(n70865) );
  XNOR2X1 U42979 ( .A(n70860), .B(n70859), .Y(n41381) );
  XNOR2X1 U42980 ( .A(n67702), .B(n67698), .Y(n41382) );
  AND2X1 U42981 ( .A(n68077), .B(n68078), .Y(n41384) );
  XOR2X1 U42982 ( .A(n62480), .B(n41385), .Y(n62428) );
  XNOR2X1 U42983 ( .A(n62479), .B(n62481), .Y(n41385) );
  XNOR2X1 U42984 ( .A(n69860), .B(n41386), .Y(n69922) );
  XNOR2X1 U42985 ( .A(n69936), .B(n69859), .Y(n41386) );
  NAND2X1 U42986 ( .A(n63728), .B(n41387), .Y(n64247) );
  AND2X1 U42987 ( .A(n63726), .B(n63725), .Y(n41387) );
  XOR2X1 U42988 ( .A(n65852), .B(n66198), .Y(n66204) );
  OR2X1 U42989 ( .A(n62423), .B(n41388), .Y(n62426) );
  AND2X1 U42990 ( .A(n39899), .B(n62424), .Y(n41388) );
  XNOR2X1 U42991 ( .A(n64812), .B(n64997), .Y(n41389) );
  XNOR2X1 U42992 ( .A(n66161), .B(n41390), .Y(n66462) );
  XNOR2X1 U42993 ( .A(n66443), .B(n66160), .Y(n41390) );
  XOR2X1 U42994 ( .A(n64026), .B(n64019), .Y(n64025) );
  AND2X1 U42995 ( .A(n63502), .B(n63507), .Y(n41391) );
  AND2X1 U42996 ( .A(n71753), .B(n71754), .Y(n41392) );
  XNOR2X1 U42997 ( .A(n66937), .B(n41393), .Y(n67213) );
  XOR2X1 U42998 ( .A(n43628), .B(n66936), .Y(n41393) );
  XOR2X1 U42999 ( .A(n61110), .B(n60734), .Y(n60889) );
  XOR2X1 U43000 ( .A(n63301), .B(n62992), .Y(n41394) );
  XNOR2X1 U43001 ( .A(n65177), .B(n41395), .Y(n65182) );
  XOR2X1 U43002 ( .A(n43638), .B(n65178), .Y(n41395) );
  XNOR2X1 U43003 ( .A(n41396), .B(n70913), .Y(n70574) );
  XOR2X1 U43004 ( .A(n70912), .B(n43569), .Y(n41396) );
  XOR2X1 U43005 ( .A(n68597), .B(n68598), .Y(n68602) );
  XOR2X1 U43006 ( .A(n63441), .B(n41397), .Y(n63434) );
  XNOR2X1 U43007 ( .A(n63671), .B(n63384), .Y(n41397) );
  AND2X1 U43008 ( .A(n40971), .B(n43658), .Y(n41398) );
  AND2X1 U43009 ( .A(n66196), .B(n66195), .Y(n41399) );
  XOR2X1 U43010 ( .A(n63603), .B(n63599), .Y(n63476) );
  XNOR2X1 U43011 ( .A(n41400), .B(n62491), .Y(n62493) );
  XOR2X1 U43012 ( .A(n62488), .B(n62490), .Y(n41400) );
  XNOR2X1 U43013 ( .A(n69617), .B(n69846), .Y(n69854) );
  XNOR2X1 U43014 ( .A(n67017), .B(n41401), .Y(n67508) );
  XNOR2X1 U43015 ( .A(n67014), .B(n67016), .Y(n41401) );
  AND2X1 U43016 ( .A(n43567), .B(n68279), .Y(n41402) );
  AND2X1 U43017 ( .A(n67515), .B(n67834), .Y(n41403) );
  AND2X1 U43018 ( .A(n71752), .B(n43656), .Y(n41404) );
  XNOR2X1 U43019 ( .A(n67576), .B(n41405), .Y(n67276) );
  XOR2X1 U43020 ( .A(n43552), .B(n67575), .Y(n41405) );
  XNOR2X1 U43021 ( .A(n40307), .B(n41406), .Y(n67316) );
  XNOR2X1 U43022 ( .A(n67814), .B(n67314), .Y(n41406) );
  XNOR2X1 U43023 ( .A(n66445), .B(n67026), .Y(n41407) );
  XNOR2X1 U43024 ( .A(n66817), .B(n41408), .Y(n66829) );
  XNOR2X1 U43025 ( .A(n66816), .B(n66815), .Y(n41408) );
  OR2X1 U43026 ( .A(n64993), .B(n64992), .Y(n65353) );
  XOR2X1 U43027 ( .A(n63671), .B(n63439), .Y(n63450) );
  XNOR2X1 U43028 ( .A(n67323), .B(n41409), .Y(n67503) );
  XNOR2X1 U43029 ( .A(n67155), .B(n67154), .Y(n41409) );
  OR2X1 U43030 ( .A(n66087), .B(n41411), .Y(n66334) );
  AND2X1 U43031 ( .A(n66092), .B(n66091), .Y(n41411) );
  AND2X1 U43032 ( .A(n43567), .B(n68277), .Y(n41412) );
  AND2X1 U43033 ( .A(n66540), .B(n43531), .Y(n41413) );
  XNOR2X1 U43034 ( .A(n66035), .B(n66036), .Y(n66447) );
  XNOR2X1 U43035 ( .A(n66039), .B(n41414), .Y(n66171) );
  XNOR2X1 U43036 ( .A(n66036), .B(n65811), .Y(n41414) );
  AND2X1 U43037 ( .A(n68545), .B(n43697), .Y(n41415) );
  NOR2X1 U43038 ( .A(n67898), .B(n41417), .Y(n41416) );
  INVX1 U43039 ( .A(n43514), .Y(n41417) );
  XOR2X1 U43040 ( .A(n68306), .B(n68187), .Y(n68768) );
  XOR2X1 U43041 ( .A(n68961), .B(n68757), .Y(n69318) );
  XNOR2X1 U43042 ( .A(n68939), .B(n69305), .Y(n69498) );
  XOR2X1 U43043 ( .A(n67803), .B(n68738), .Y(n68310) );
  AND2X1 U43044 ( .A(n41729), .B(n68966), .Y(n41418) );
  AND2X1 U43045 ( .A(n70428), .B(n70429), .Y(n41419) );
  XNOR2X1 U43046 ( .A(n64460), .B(n41420), .Y(n64716) );
  XOR2X1 U43047 ( .A(n64455), .B(n64459), .Y(n41420) );
  XNOR2X1 U43048 ( .A(n64463), .B(n41421), .Y(n64473) );
  XNOR2X1 U43049 ( .A(n64462), .B(n64716), .Y(n41421) );
  XNOR2X1 U43050 ( .A(n64472), .B(n41422), .Y(n64477) );
  XOR2X1 U43051 ( .A(n64473), .B(n64703), .Y(n41422) );
  XOR2X1 U43052 ( .A(n64184), .B(n64183), .Y(n41423) );
  AND2X1 U43053 ( .A(n66099), .B(n66338), .Y(n41424) );
  XNOR2X1 U43054 ( .A(n40261), .B(n41425), .Y(n65708) );
  XNOR2X1 U43055 ( .A(n65359), .B(n65360), .Y(n41425) );
  AND2X1 U43056 ( .A(n69287), .B(n69286), .Y(n41426) );
  XOR2X1 U43057 ( .A(n65988), .B(n65987), .Y(n41427) );
  XOR2X1 U43058 ( .A(n64676), .B(n64675), .Y(n41428) );
  XOR2X1 U43059 ( .A(n69947), .B(n41638), .Y(n70270) );
  AND2X1 U43060 ( .A(n66069), .B(n41429), .Y(n66050) );
  AND2X1 U43061 ( .A(n66066), .B(n66070), .Y(n41429) );
  OR2X1 U43062 ( .A(n70115), .B(n41430), .Y(n70117) );
  OR2X1 U43063 ( .A(n39983), .B(n43587), .Y(n41430) );
  NOR2X1 U43064 ( .A(n68838), .B(n41417), .Y(n41431) );
  XNOR2X1 U43065 ( .A(n68078), .B(n41432), .Y(n68179) );
  XNOR2X1 U43066 ( .A(n67787), .B(n67786), .Y(n41432) );
  OR2X1 U43067 ( .A(n41433), .B(n64473), .Y(n64707) );
  AND2X1 U43068 ( .A(n64378), .B(n64377), .Y(n41433) );
  XOR2X1 U43069 ( .A(n64816), .B(n64817), .Y(n64819) );
  XNOR2X1 U43070 ( .A(n66681), .B(n41434), .Y(n67344) );
  XNOR2X1 U43071 ( .A(n66788), .B(n66434), .Y(n41434) );
  XOR2X1 U43072 ( .A(n69647), .B(n69952), .Y(n70087) );
  XNOR2X1 U43073 ( .A(n65453), .B(n65118), .Y(n65304) );
  XNOR2X1 U43074 ( .A(n60442), .B(n60441), .Y(n41436) );
  XNOR2X1 U43075 ( .A(n63866), .B(n41437), .Y(n64191) );
  XNOR2X1 U43076 ( .A(n63865), .B(n63864), .Y(n41437) );
  OR2X1 U43077 ( .A(n68442), .B(n41438), .Y(n68720) );
  AND2X1 U43078 ( .A(n68444), .B(n68443), .Y(n41438) );
  AND2X1 U43079 ( .A(n68077), .B(n68079), .Y(n41439) );
  OR2X1 U43080 ( .A(n68045), .B(n41440), .Y(n68048) );
  OR2X1 U43081 ( .A(n68047), .B(n68046), .Y(n41440) );
  XOR2X1 U43082 ( .A(n68169), .B(n68429), .Y(n68436) );
  AND2X1 U43083 ( .A(n63533), .B(n63532), .Y(n63252) );
  AND2X1 U43084 ( .A(n67811), .B(n67810), .Y(n41441) );
  XOR2X1 U43085 ( .A(n68718), .B(n68996), .Y(n69450) );
  XNOR2X1 U43086 ( .A(n69468), .B(n41443), .Y(n41442) );
  XOR2X1 U43087 ( .A(n69444), .B(n69142), .Y(n41443) );
  OR2X1 U43088 ( .A(n64884), .B(n41444), .Y(n65234) );
  AND2X1 U43089 ( .A(n64885), .B(n43532), .Y(n41444) );
  AND2X1 U43090 ( .A(n41445), .B(n41446), .Y(n67363) );
  NOR2X1 U43091 ( .A(n67341), .B(n67147), .Y(n41445) );
  NOR2X1 U43092 ( .A(n67145), .B(n67144), .Y(n41446) );
  OR2X1 U43093 ( .A(n68699), .B(n41447), .Y(n69005) );
  AND2X1 U43094 ( .A(n68703), .B(n68702), .Y(n41447) );
  XOR2X1 U43095 ( .A(n69464), .B(n41726), .Y(n41448) );
  OR2X1 U43096 ( .A(n71660), .B(n41449), .Y(n71672) );
  AND2X1 U43097 ( .A(n71670), .B(n43549), .Y(n41449) );
  AND2X1 U43098 ( .A(n41450), .B(n39746), .Y(n69504) );
  AND2X1 U43099 ( .A(n43592), .B(n38962), .Y(n41450) );
  XOR2X1 U43100 ( .A(n66446), .B(n40122), .Y(n66457) );
  XOR2X1 U43101 ( .A(n69810), .B(n69965), .Y(n69675) );
  AND2X1 U43102 ( .A(n71078), .B(n71080), .Y(n41451) );
  XOR2X1 U43103 ( .A(n71239), .B(n41452), .Y(n71386) );
  XNOR2X1 U43104 ( .A(n71606), .B(n71085), .Y(n41452) );
  XOR2X1 U43105 ( .A(n41657), .B(n70725), .Y(n41453) );
  OR2X1 U43106 ( .A(n67918), .B(n41454), .Y(n68540) );
  INVX1 U43107 ( .A(n43698), .Y(n41454) );
  XNOR2X1 U43108 ( .A(n67806), .B(n41455), .Y(n67826) );
  XNOR2X1 U43109 ( .A(n39972), .B(n67816), .Y(n41455) );
  AND2X1 U43110 ( .A(n41689), .B(n63794), .Y(n41456) );
  AND2X1 U43111 ( .A(n63472), .B(n63473), .Y(n41457) );
  OR2X1 U43112 ( .A(n41458), .B(n41459), .Y(n71083) );
  NOR2X1 U43113 ( .A(n72353), .B(n71374), .Y(n41458) );
  NOR2X1 U43114 ( .A(n71082), .B(n71081), .Y(n41459) );
  XOR2X1 U43115 ( .A(n72058), .B(n72059), .Y(n72060) );
  XNOR2X1 U43116 ( .A(n72159), .B(n72069), .Y(n72070) );
  AND2X1 U43117 ( .A(n71373), .B(n41460), .Y(n71076) );
  AND2X1 U43118 ( .A(n71080), .B(n71078), .Y(n41460) );
  AND2X1 U43119 ( .A(n70708), .B(n70924), .Y(n41461) );
  AND2X1 U43120 ( .A(n70904), .B(n70903), .Y(n41462) );
  XNOR2X1 U43121 ( .A(n64439), .B(n64440), .Y(n64739) );
  XNOR2X1 U43122 ( .A(n70716), .B(n70717), .Y(n70719) );
  XNOR2X1 U43123 ( .A(n64119), .B(n41463), .Y(n64139) );
  XOR2X1 U43124 ( .A(n64134), .B(n64133), .Y(n41463) );
  XOR2X1 U43125 ( .A(n70728), .B(n70731), .Y(n70734) );
  AND2X1 U43126 ( .A(n68681), .B(n41464), .Y(n68686) );
  AND2X1 U43127 ( .A(n68688), .B(n43983), .Y(n41464) );
  NOR2X1 U43128 ( .A(n41466), .B(n66548), .Y(n41465) );
  INVX1 U43129 ( .A(n43699), .Y(n41466) );
  XNOR2X1 U43130 ( .A(n69685), .B(n41467), .Y(n69805) );
  XNOR2X1 U43131 ( .A(n69684), .B(n69681), .Y(n41467) );
  XNOR2X1 U43132 ( .A(n70681), .B(n41469), .Y(n41468) );
  XOR2X1 U43133 ( .A(n70368), .B(n70064), .Y(n41469) );
  XOR2X1 U43134 ( .A(n70698), .B(n70940), .Y(n70935) );
  AND2X1 U43135 ( .A(n65225), .B(n65224), .Y(n41470) );
  XNOR2X1 U43136 ( .A(n71622), .B(n41471), .Y(n71625) );
  AND2X1 U43137 ( .A(n71624), .B(n71623), .Y(n41471) );
  NAND2X1 U43138 ( .A(n70055), .B(n41472), .Y(n70059) );
  AND2X1 U43139 ( .A(n70058), .B(n70057), .Y(n41472) );
  XNOR2X1 U43140 ( .A(n70055), .B(n41473), .Y(n70065) );
  XNOR2X1 U43141 ( .A(n70054), .B(n70052), .Y(n41473) );
  XNOR2X1 U43142 ( .A(n64146), .B(n41474), .Y(n64448) );
  XNOR2X1 U43143 ( .A(n64119), .B(n64060), .Y(n41474) );
  XNOR2X1 U43144 ( .A(n63843), .B(n41475), .Y(n64147) );
  XNOR2X1 U43145 ( .A(n64060), .B(n64062), .Y(n41475) );
  XOR2X1 U43146 ( .A(n67376), .B(n67075), .Y(n67442) );
  XNOR2X1 U43147 ( .A(n65416), .B(n64806), .Y(n65087) );
  XOR2X1 U43148 ( .A(n66703), .B(n41476), .Y(n66330) );
  XNOR2X1 U43149 ( .A(n66362), .B(n66154), .Y(n41476) );
  XOR2X1 U43150 ( .A(n70616), .B(n70617), .Y(n70367) );
  OR2X1 U43151 ( .A(n41477), .B(n41478), .Y(n71383) );
  NOR2X1 U43152 ( .A(n43594), .B(n71377), .Y(n41477) );
  NOR2X1 U43153 ( .A(n71608), .B(n71376), .Y(n41478) );
  AND2X1 U43154 ( .A(n65399), .B(n41479), .Y(n65403) );
  OR2X1 U43155 ( .A(n65401), .B(n65400), .Y(n41479) );
  XOR2X1 U43156 ( .A(n65747), .B(n65748), .Y(n65767) );
  XOR2X1 U43157 ( .A(n66409), .B(n67109), .Y(n67122) );
  AND2X1 U43158 ( .A(n66147), .B(n66148), .Y(n66150) );
  AND2X1 U43159 ( .A(n64274), .B(n43514), .Y(n41480) );
  AND2X1 U43160 ( .A(n72155), .B(n72154), .Y(n41481) );
  XOR2X1 U43161 ( .A(n63421), .B(n63393), .Y(n63414) );
  AND2X1 U43162 ( .A(n65389), .B(n41482), .Y(n65397) );
  AND2X1 U43163 ( .A(n65396), .B(n43861), .Y(n41482) );
  AND2X1 U43164 ( .A(n43840), .B(n42640), .Y(n41483) );
  AND2X1 U43165 ( .A(n63412), .B(n63411), .Y(n41484) );
  XOR2X1 U43166 ( .A(n41239), .B(n69688), .Y(n41485) );
  XOR2X1 U43167 ( .A(n66401), .B(n66745), .Y(n66752) );
  XNOR2X1 U43168 ( .A(n65754), .B(n41486), .Y(n65373) );
  XOR2X1 U43169 ( .A(n65761), .B(n65792), .Y(n41486) );
  AND2X1 U43170 ( .A(n62810), .B(n62809), .Y(n41487) );
  OR2X1 U43171 ( .A(n70354), .B(n70355), .Y(n70361) );
  XNOR2X1 U43172 ( .A(n70613), .B(n41488), .Y(n70617) );
  OR2X1 U43173 ( .A(n70366), .B(n70365), .Y(n41488) );
  AND2X1 U43174 ( .A(n43631), .B(n72595), .Y(n41489) );
  AND2X1 U43175 ( .A(n43850), .B(n43607), .Y(n41490) );
  XOR2X1 U43176 ( .A(n71350), .B(n71351), .Y(n71357) );
  OR2X1 U43177 ( .A(n72146), .B(n41491), .Y(n72147) );
  AND2X1 U43178 ( .A(n43535), .B(n72177), .Y(n41491) );
  XNOR2X1 U43179 ( .A(n70030), .B(n70031), .Y(n41492) );
  XNOR2X1 U43180 ( .A(n71811), .B(n72021), .Y(n71813) );
  OR2X1 U43181 ( .A(n70614), .B(n41493), .Y(n70611) );
  XOR2X1 U43182 ( .A(n70662), .B(n70610), .Y(n41493) );
  XOR2X1 U43183 ( .A(n66749), .B(n67098), .Y(n67385) );
  AND2X1 U43184 ( .A(n63083), .B(n63082), .Y(n41494) );
  XOR2X1 U43185 ( .A(n71596), .B(n71597), .Y(n71598) );
  XOR2X1 U43186 ( .A(n41531), .B(n71998), .Y(n71820) );
  AND2X1 U43187 ( .A(n44035), .B(n42633), .Y(n41495) );
  OR2X1 U43188 ( .A(n69127), .B(n41496), .Y(n68645) );
  AND2X1 U43189 ( .A(n69126), .B(n69128), .Y(n41496) );
  AND2X1 U43190 ( .A(n62799), .B(n62798), .Y(n41497) );
  AND2X1 U43191 ( .A(n43962), .B(n39653), .Y(n41498) );
  AND2X1 U43192 ( .A(n42657), .B(n43852), .Y(n41499) );
  XNOR2X1 U43193 ( .A(n69715), .B(n41500), .Y(n69385) );
  XOR2X1 U43194 ( .A(n69367), .B(n69716), .Y(n41500) );
  XNOR2X1 U43195 ( .A(n41501), .B(n67416), .Y(n67762) );
  XOR2X1 U43196 ( .A(n67415), .B(n67752), .Y(n41501) );
  XNOR2X1 U43197 ( .A(n68648), .B(n41502), .Y(n69093) );
  XNOR2X1 U43198 ( .A(n68646), .B(n68647), .Y(n41502) );
  XOR2X1 U43199 ( .A(n70337), .B(n70336), .Y(n70340) );
  AND2X1 U43200 ( .A(n41705), .B(n67756), .Y(n41503) );
  XNOR2X1 U43201 ( .A(n69094), .B(n41504), .Y(n68644) );
  XNOR2X1 U43202 ( .A(n69093), .B(n69096), .Y(n41504) );
  XOR2X1 U43203 ( .A(n71503), .B(n71570), .Y(n71505) );
  XOR2X1 U43204 ( .A(n71994), .B(n72521), .Y(n72545) );
  AND2X1 U43205 ( .A(n43952), .B(n43518), .Y(n41505) );
  AND2X1 U43206 ( .A(n42660), .B(n43954), .Y(n41506) );
  XNOR2X1 U43207 ( .A(n69082), .B(n68660), .Y(n69076) );
  XNOR2X1 U43208 ( .A(n69080), .B(n69108), .Y(n69117) );
  AND2X1 U43209 ( .A(n43952), .B(n43496), .Y(n41507) );
  XOR2X1 U43210 ( .A(n69723), .B(n69727), .Y(n69752) );
  XOR2X1 U43211 ( .A(n70015), .B(n70296), .Y(n70331) );
  AND2X1 U43212 ( .A(n43492), .B(n43953), .Y(n41508) );
  XOR2X1 U43213 ( .A(n69767), .B(n69768), .Y(n69773) );
  AND2X1 U43214 ( .A(n43889), .B(n43608), .Y(n41509) );
  XOR2X1 U43215 ( .A(n71320), .B(n71025), .Y(n71329) );
  XOR2X1 U43216 ( .A(n67079), .B(n41711), .Y(n66770) );
  AND2X1 U43217 ( .A(n43918), .B(n39653), .Y(n41510) );
  XNOR2X1 U43218 ( .A(n41700), .B(n71885), .Y(n41511) );
  XNOR2X1 U43219 ( .A(n41696), .B(n71881), .Y(n41512) );
  AND2X1 U43220 ( .A(n43927), .B(n42632), .Y(n41513) );
  XOR2X1 U43221 ( .A(n71909), .B(n71910), .Y(n71922) );
  AND2X1 U43222 ( .A(n43927), .B(n43497), .Y(n41514) );
  AND2X1 U43223 ( .A(n43928), .B(n39961), .Y(n41515) );
  XOR2X1 U43224 ( .A(n41703), .B(n41511), .Y(n41516) );
  AND2X1 U43225 ( .A(n43942), .B(n43607), .Y(n41517) );
  AND2X1 U43226 ( .A(n42711), .B(n43973), .Y(n41518) );
  AND2X1 U43227 ( .A(n43942), .B(n43486), .Y(n41519) );
  XOR2X1 U43228 ( .A(n41685), .B(n72374), .Y(n72384) );
  XOR2X1 U43229 ( .A(n41684), .B(n72311), .Y(n41520) );
  AND2X1 U43230 ( .A(n43491), .B(n43972), .Y(n41521) );
  AND2X1 U43231 ( .A(n67683), .B(n67478), .Y(n41522) );
  AND2X1 U43232 ( .A(n43982), .B(n38311), .Y(n41523) );
  XNOR2X1 U43233 ( .A(n72473), .B(n41524), .Y(n72481) );
  XOR2X1 U43234 ( .A(n72475), .B(n72474), .Y(n41524) );
  XOR2X1 U43235 ( .A(n68167), .B(n68421), .Y(n68075) );
  XNOR2X1 U43236 ( .A(n41525), .B(n72730), .Y(n72731) );
  XOR2X1 U43237 ( .A(n43708), .B(n72729), .Y(n41525) );
  AND2X1 U43238 ( .A(n43972), .B(n43517), .Y(n41526) );
  AND2X1 U43239 ( .A(n42711), .B(n44017), .Y(n41527) );
  AND2X1 U43240 ( .A(n43999), .B(n39844), .Y(n41528) );
  AND2X1 U43241 ( .A(n43491), .B(n44016), .Y(n41529) );
  XOR2X1 U43242 ( .A(n43558), .B(n43537), .Y(n70752) );
  AND2X1 U43243 ( .A(n44016), .B(n43517), .Y(n41530) );
  XOR2X1 U43244 ( .A(n43616), .B(n43601), .Y(n41531) );
  AND2X1 U43245 ( .A(n57680), .B(n57717), .Y(n41532) );
  OR2X1 U43246 ( .A(n42711), .B(n59075), .Y(n59081) );
  OR2X1 U43247 ( .A(n41533), .B(n41534), .Y(n65290) );
  AND2X1 U43248 ( .A(n64949), .B(n64948), .Y(n41533) );
  AND2X1 U43249 ( .A(n42005), .B(n65154), .Y(n41534) );
  AND2X1 U43250 ( .A(n62515), .B(n41536), .Y(n62513) );
  INVX1 U43251 ( .A(n62511), .Y(n41536) );
  AND2X1 U43252 ( .A(n63744), .B(n41967), .Y(n41537) );
  AND2X1 U43253 ( .A(n66964), .B(n66850), .Y(n66639) );
  OR2X1 U43254 ( .A(n41538), .B(n59444), .Y(n59383) );
  NOR2X1 U43255 ( .A(n59443), .B(n39090), .Y(n41538) );
  NAND2X1 U43256 ( .A(n38791), .B(n59419), .Y(n59348) );
  OR2X1 U43257 ( .A(n59951), .B(n41539), .Y(n60274) );
  AND2X1 U43258 ( .A(n40586), .B(n59952), .Y(n41539) );
  AND2X1 U43259 ( .A(n41540), .B(n41541), .Y(n42840) );
  NAND2X1 U43260 ( .A(n59204), .B(n59205), .Y(n41540) );
  NAND2X1 U43261 ( .A(n59207), .B(n59206), .Y(n41541) );
  NAND2X1 U43262 ( .A(n41542), .B(n59307), .Y(n59206) );
  INVX1 U43263 ( .A(n59205), .Y(n41542) );
  AND2X1 U43264 ( .A(n63141), .B(n62860), .Y(n62861) );
  OR2X1 U43265 ( .A(n41543), .B(n41544), .Y(n60727) );
  AND2X1 U43266 ( .A(n60299), .B(n60298), .Y(n41543) );
  AND2X1 U43267 ( .A(n41944), .B(n60302), .Y(n41544) );
  OR2X1 U43268 ( .A(n41545), .B(n41546), .Y(n60299) );
  AND2X1 U43269 ( .A(n59860), .B(n59859), .Y(n41545) );
  AND2X1 U43270 ( .A(n59862), .B(n59861), .Y(n41546) );
  OR2X1 U43271 ( .A(n41547), .B(n41548), .Y(n59856) );
  AND2X1 U43272 ( .A(n59848), .B(n59849), .Y(n41547) );
  AND2X1 U43273 ( .A(n59851), .B(n59850), .Y(n41548) );
  OR2X1 U43274 ( .A(n60900), .B(n41549), .Y(n61289) );
  AND2X1 U43275 ( .A(n39750), .B(n60901), .Y(n41549) );
  OR2X1 U43276 ( .A(n63372), .B(n41550), .Y(n63030) );
  AND2X1 U43277 ( .A(n38851), .B(n63028), .Y(n41550) );
  OR2X1 U43278 ( .A(n59607), .B(n59606), .Y(n59608) );
  AND2X1 U43279 ( .A(n64640), .B(n41551), .Y(n64656) );
  AND2X1 U43280 ( .A(n42047), .B(n64641), .Y(n41551) );
  AND2X1 U43281 ( .A(n64338), .B(n64686), .Y(n41552) );
  AND2X1 U43282 ( .A(n62378), .B(n41553), .Y(n62377) );
  INVX1 U43283 ( .A(n62376), .Y(n41553) );
  OR2X1 U43284 ( .A(n60193), .B(n41554), .Y(n60914) );
  NOR2X1 U43285 ( .A(n38253), .B(n60196), .Y(n41554) );
  XNOR2X1 U43286 ( .A(n66646), .B(n41555), .Y(n66977) );
  XOR2X1 U43287 ( .A(n66482), .B(n66645), .Y(n41555) );
  AND2X1 U43288 ( .A(n64487), .B(n41556), .Y(n64489) );
  INVX1 U43289 ( .A(n64488), .Y(n41556) );
  AND2X1 U43290 ( .A(n64980), .B(n40439), .Y(n41557) );
  NAND2X1 U43291 ( .A(n65268), .B(n41558), .Y(n65267) );
  OR2X1 U43292 ( .A(n64931), .B(n65270), .Y(n41558) );
  XNOR2X1 U43293 ( .A(n38515), .B(n41560), .Y(n41559) );
  XOR2X1 U43294 ( .A(n65256), .B(n65255), .Y(n41560) );
  OR2X1 U43295 ( .A(n60683), .B(n42835), .Y(n61049) );
  XNOR2X1 U43296 ( .A(n62515), .B(n62511), .Y(n41561) );
  AND2X1 U43297 ( .A(n41999), .B(n38377), .Y(n41562) );
  XOR2X1 U43298 ( .A(n39926), .B(n63027), .Y(n63455) );
  OR2X1 U43299 ( .A(n59791), .B(n59792), .Y(n59793) );
  XNOR2X1 U43300 ( .A(n65479), .B(n41563), .Y(n65481) );
  XOR2X1 U43301 ( .A(n65478), .B(n65656), .Y(n41563) );
  AND2X1 U43302 ( .A(n42020), .B(n64238), .Y(n41564) );
  XNOR2X1 U43303 ( .A(n61205), .B(n41565), .Y(n61216) );
  OR2X1 U43304 ( .A(n60981), .B(n60980), .Y(n41565) );
  OR2X1 U43305 ( .A(n59994), .B(n59995), .Y(n59996) );
  AND2X1 U43306 ( .A(n63750), .B(n64031), .Y(n41566) );
  AND2X1 U43307 ( .A(n65644), .B(n65639), .Y(n65643) );
  OR2X1 U43308 ( .A(n41567), .B(n41568), .Y(n66519) );
  AND2X1 U43309 ( .A(n64921), .B(n65177), .Y(n41567) );
  AND2X1 U43310 ( .A(n64923), .B(n64922), .Y(n41568) );
  XNOR2X1 U43311 ( .A(n59443), .B(n59446), .Y(n59448) );
  XNOR2X1 U43312 ( .A(n64978), .B(n41569), .Y(n65475) );
  XNOR2X1 U43313 ( .A(n64966), .B(n64977), .Y(n41569) );
  OR2X1 U43314 ( .A(n41570), .B(n41571), .Y(n59853) );
  AND2X1 U43315 ( .A(n59844), .B(n59660), .Y(n41570) );
  AND2X1 U43316 ( .A(n59663), .B(n59662), .Y(n41571) );
  AND2X1 U43317 ( .A(n41973), .B(n40361), .Y(n41572) );
  AND2X1 U43318 ( .A(n66303), .B(n66302), .Y(n41573) );
  XNOR2X1 U43319 ( .A(n60934), .B(n41574), .Y(n60974) );
  OR2X1 U43320 ( .A(n60628), .B(n60627), .Y(n41574) );
  OR2X1 U43321 ( .A(n59675), .B(n59674), .Y(n60227) );
  AND2X1 U43322 ( .A(n41967), .B(n63743), .Y(n41575) );
  AND2X1 U43323 ( .A(n64976), .B(n64977), .Y(n41576) );
  XNOR2X1 U43324 ( .A(n59330), .B(n41577), .Y(n59318) );
  XOR2X1 U43325 ( .A(n39114), .B(n59278), .Y(n41577) );
  XOR2X1 U43326 ( .A(n41578), .B(n64869), .Y(n65251) );
  OR2X1 U43327 ( .A(n39259), .B(n65271), .Y(n41578) );
  AND2X1 U43328 ( .A(n41973), .B(n64953), .Y(n41579) );
  OR2X1 U43329 ( .A(n59968), .B(n41580), .Y(n60294) );
  AND2X1 U43330 ( .A(n39313), .B(n59969), .Y(n41580) );
  XOR2X1 U43331 ( .A(n63917), .B(n63665), .Y(n63991) );
  XNOR2X1 U43332 ( .A(n59193), .B(n41581), .Y(n59215) );
  XNOR2X1 U43333 ( .A(n59192), .B(n59191), .Y(n41581) );
  OR2X1 U43334 ( .A(n41582), .B(n41583), .Y(n63019) );
  AND2X1 U43335 ( .A(n62381), .B(n62380), .Y(n41582) );
  AND2X1 U43336 ( .A(n62390), .B(n62389), .Y(n41583) );
  AND2X1 U43337 ( .A(n65496), .B(n65495), .Y(n41584) );
  XNOR2X1 U43338 ( .A(n68006), .B(n67996), .Y(n67997) );
  OR2X1 U43339 ( .A(n41585), .B(n41586), .Y(n60283) );
  AND2X1 U43340 ( .A(n59961), .B(n59960), .Y(n41585) );
  AND2X1 U43341 ( .A(n59965), .B(n59964), .Y(n41586) );
  OR2X1 U43342 ( .A(n59591), .B(n41587), .Y(n59767) );
  OR2X1 U43343 ( .A(n61074), .B(n41588), .Y(n61269) );
  AND2X1 U43344 ( .A(n36686), .B(n61075), .Y(n41588) );
  XOR2X1 U43345 ( .A(n41589), .B(n39537), .Y(n62538) );
  XOR2X1 U43346 ( .A(n62527), .B(n62526), .Y(n41589) );
  XNOR2X1 U43347 ( .A(n40530), .B(n41590), .Y(n66968) );
  XNOR2X1 U43348 ( .A(n66482), .B(n66481), .Y(n41590) );
  OR2X1 U43349 ( .A(n60723), .B(n41591), .Y(n60902) );
  AND2X1 U43350 ( .A(n39695), .B(n38289), .Y(n41591) );
  XNOR2X1 U43351 ( .A(n60904), .B(n60725), .Y(n60726) );
  OR2X1 U43352 ( .A(n63112), .B(n41592), .Y(n63114) );
  AND2X1 U43353 ( .A(n39987), .B(n63113), .Y(n41592) );
  OR2X1 U43354 ( .A(n60110), .B(n60111), .Y(n60112) );
  AND2X1 U43355 ( .A(n65485), .B(n65511), .Y(n41593) );
  NAND2X1 U43356 ( .A(n41594), .B(n41595), .Y(n61283) );
  OR2X1 U43357 ( .A(n60905), .B(n60904), .Y(n41594) );
  OR2X1 U43358 ( .A(n60909), .B(n60908), .Y(n41595) );
  OR2X1 U43359 ( .A(n63989), .B(n41596), .Y(n64508) );
  AND2X1 U43360 ( .A(n63994), .B(n63993), .Y(n41596) );
  XOR2X1 U43361 ( .A(n64496), .B(n64341), .Y(n64683) );
  OR2X1 U43362 ( .A(n60083), .B(n41597), .Y(n60055) );
  AND2X1 U43363 ( .A(n60084), .B(n60082), .Y(n41597) );
  XNOR2X1 U43364 ( .A(n61052), .B(n41598), .Y(n61063) );
  OR2X1 U43365 ( .A(n60693), .B(n60692), .Y(n41598) );
  XOR2X1 U43366 ( .A(n63358), .B(n63362), .Y(n63614) );
  AND2X1 U43367 ( .A(n41983), .B(n63132), .Y(n41599) );
  OR2X1 U43368 ( .A(n63442), .B(n41600), .Y(n63719) );
  AND2X1 U43369 ( .A(n63451), .B(n63450), .Y(n41600) );
  OR2X1 U43370 ( .A(n63032), .B(n41601), .Y(n63039) );
  XNOR2X1 U43371 ( .A(n64510), .B(n64245), .Y(n64607) );
  AND2X1 U43372 ( .A(n64862), .B(n64861), .Y(n41602) );
  INVX1 U43373 ( .A(n41998), .Y(n41603) );
  NOR2X1 U43374 ( .A(n63900), .B(n63899), .Y(n41604) );
  XNOR2X1 U43375 ( .A(n41605), .B(n59454), .Y(n59528) );
  XOR2X1 U43376 ( .A(n59521), .B(n59520), .Y(n41605) );
  AND2X1 U43377 ( .A(n42020), .B(n64240), .Y(n41606) );
  AND2X1 U43378 ( .A(n65486), .B(n41607), .Y(n65487) );
  AND2X1 U43379 ( .A(n44004), .B(n65159), .Y(n41607) );
  XOR2X1 U43380 ( .A(n63132), .B(n63026), .Y(n63130) );
  AND2X1 U43381 ( .A(n64980), .B(n64982), .Y(n41608) );
  OR2X1 U43382 ( .A(n60340), .B(n60341), .Y(n60342) );
  XOR2X1 U43383 ( .A(n66995), .B(n66847), .Y(n66848) );
  XOR2X1 U43384 ( .A(n63901), .B(n63913), .Y(n63664) );
  XNOR2X1 U43385 ( .A(n41610), .B(n59763), .Y(n59665) );
  XOR2X1 U43386 ( .A(n59764), .B(n59762), .Y(n41610) );
  XNOR2X1 U43387 ( .A(n36627), .B(n41611), .Y(n66488) );
  XNOR2X1 U43388 ( .A(n66646), .B(n66209), .Y(n41611) );
  OR2X1 U43389 ( .A(n64674), .B(n64673), .Y(n41612) );
  OR2X1 U43390 ( .A(n61101), .B(n41613), .Y(n63035) );
  XNOR2X1 U43391 ( .A(n62494), .B(n41614), .Y(n62500) );
  XNOR2X1 U43392 ( .A(n62492), .B(n62493), .Y(n41614) );
  XNOR2X1 U43393 ( .A(n63991), .B(n41615), .Y(n63728) );
  XNOR2X1 U43394 ( .A(n63731), .B(n63736), .Y(n41615) );
  XOR2X1 U43395 ( .A(n63978), .B(n63927), .Y(n64252) );
  XNOR2X1 U43396 ( .A(n63119), .B(n63127), .Y(n41616) );
  XNOR2X1 U43397 ( .A(n63361), .B(n63017), .Y(n63018) );
  OR2X1 U43398 ( .A(n64008), .B(n41617), .Y(n64329) );
  AND2X1 U43399 ( .A(n64015), .B(n64014), .Y(n41617) );
  OR2X1 U43400 ( .A(n60461), .B(n60462), .Y(n60463) );
  AND2X1 U43401 ( .A(n66202), .B(n66203), .Y(n41618) );
  OR2X1 U43402 ( .A(n67183), .B(n41619), .Y(n66295) );
  AND2X1 U43403 ( .A(n66627), .B(n66626), .Y(n41619) );
  XOR2X1 U43404 ( .A(n67315), .B(n67173), .Y(n67531) );
  XOR2X1 U43405 ( .A(n68482), .B(n68483), .Y(n41620) );
  XNOR2X1 U43406 ( .A(n64946), .B(n41621), .Y(n65155) );
  XNOR2X1 U43407 ( .A(n65475), .B(n64855), .Y(n41621) );
  OR2X1 U43408 ( .A(n60804), .B(n60805), .Y(n60806) );
  XNOR2X1 U43409 ( .A(n60446), .B(n60449), .Y(n60509) );
  AND2X1 U43410 ( .A(n68477), .B(n42992), .Y(n41622) );
  OR2X1 U43411 ( .A(n60566), .B(n41623), .Y(n61085) );
  AND2X1 U43412 ( .A(n60568), .B(n60567), .Y(n41623) );
  OR2X1 U43413 ( .A(n60932), .B(n41624), .Y(n61142) );
  AND2X1 U43414 ( .A(n38274), .B(n60934), .Y(n41624) );
  NAND2X1 U43415 ( .A(n61140), .B(n41625), .Y(n61143) );
  AND2X1 U43416 ( .A(n61142), .B(n61141), .Y(n41625) );
  OR2X1 U43417 ( .A(n64024), .B(n64025), .Y(n64333) );
  XNOR2X1 U43418 ( .A(n64993), .B(n41626), .Y(n64989) );
  XOR2X1 U43419 ( .A(n65352), .B(n64992), .Y(n41626) );
  XOR2X1 U43420 ( .A(n70242), .B(n41766), .Y(n70248) );
  XNOR2X1 U43421 ( .A(n40280), .B(n62352), .Y(n62353) );
  XNOR2X1 U43422 ( .A(n64181), .B(n41627), .Y(n63863) );
  XNOR2X1 U43423 ( .A(n64054), .B(n63862), .Y(n41627) );
  XNOR2X1 U43424 ( .A(n41628), .B(n61272), .Y(n61286) );
  XOR2X1 U43425 ( .A(n61275), .B(n61071), .Y(n41628) );
  XNOR2X1 U43426 ( .A(n41629), .B(n69300), .Y(n69293) );
  XOR2X1 U43427 ( .A(n69157), .B(n69156), .Y(n41629) );
  XOR2X1 U43428 ( .A(n60735), .B(n60305), .Y(n60564) );
  XNOR2X1 U43429 ( .A(n63728), .B(n41630), .Y(n63722) );
  XNOR2X1 U43430 ( .A(n63730), .B(n63724), .Y(n41630) );
  XNOR2X1 U43431 ( .A(n60169), .B(n41631), .Y(n60172) );
  XOR2X1 U43432 ( .A(n60170), .B(n41923), .Y(n41631) );
  XNOR2X1 U43433 ( .A(n61080), .B(n41632), .Y(n60884) );
  XNOR2X1 U43434 ( .A(n61081), .B(n61084), .Y(n41632) );
  XOR2X1 U43435 ( .A(n69842), .B(n69843), .Y(n69847) );
  XNOR2X1 U43436 ( .A(n63721), .B(n63677), .Y(n63980) );
  XNOR2X1 U43437 ( .A(n60511), .B(n41634), .Y(n60514) );
  XNOR2X1 U43438 ( .A(n60513), .B(n60512), .Y(n41634) );
  XNOR2X1 U43439 ( .A(n60524), .B(n60523), .Y(n41635) );
  XNOR2X1 U43440 ( .A(n41636), .B(n60192), .Y(n60284) );
  XOR2X1 U43441 ( .A(n60193), .B(n38253), .Y(n41636) );
  AND2X1 U43442 ( .A(n41983), .B(n63133), .Y(n41639) );
  XOR2X1 U43443 ( .A(n63986), .B(n42083), .Y(n41640) );
  XNOR2X1 U43444 ( .A(n64496), .B(n41641), .Y(n64332) );
  XNOR2X1 U43445 ( .A(n64497), .B(n64230), .Y(n41641) );
  XNOR2X1 U43446 ( .A(n65154), .B(n41642), .Y(n65168) );
  XNOR2X1 U43447 ( .A(n65163), .B(n65155), .Y(n41642) );
  OR2X1 U43448 ( .A(n61352), .B(n61353), .Y(n61354) );
  XNOR2X1 U43449 ( .A(n62344), .B(n41643), .Y(n62559) );
  XNOR2X1 U43450 ( .A(n62343), .B(n62342), .Y(n41643) );
  AND2X1 U43451 ( .A(n66202), .B(n66204), .Y(n41645) );
  XNOR2X1 U43452 ( .A(n59530), .B(n41646), .Y(n59590) );
  XNOR2X1 U43453 ( .A(n59529), .B(n59528), .Y(n41646) );
  OR2X1 U43454 ( .A(n61497), .B(n61498), .Y(n61499) );
  AND2X1 U43455 ( .A(n69679), .B(n69678), .Y(n41647) );
  XNOR2X1 U43456 ( .A(n60081), .B(n41648), .Y(n60175) );
  XNOR2X1 U43457 ( .A(n60080), .B(n60079), .Y(n41648) );
  OR2X1 U43458 ( .A(n61649), .B(n61650), .Y(n61651) );
  XNOR2X1 U43459 ( .A(n38676), .B(n41649), .Y(n62850) );
  XOR2X1 U43460 ( .A(n62378), .B(n62376), .Y(n41649) );
  NAND2X1 U43461 ( .A(n64375), .B(n41650), .Y(n64699) );
  AND2X1 U43462 ( .A(n64180), .B(n64179), .Y(n41650) );
  XNOR2X1 U43463 ( .A(n64317), .B(n41651), .Y(n64313) );
  XNOR2X1 U43464 ( .A(n64936), .B(n64234), .Y(n41651) );
  OR2X1 U43465 ( .A(n70110), .B(n72152), .Y(n69833) );
  XNOR2X1 U43466 ( .A(n64863), .B(n41652), .Y(n64675) );
  XNOR2X1 U43467 ( .A(n64864), .B(n64501), .Y(n41652) );
  XNOR2X1 U43468 ( .A(n61439), .B(n41653), .Y(n61589) );
  XOR2X1 U43469 ( .A(n61440), .B(n42053), .Y(n41653) );
  XNOR2X1 U43470 ( .A(n65280), .B(n41654), .Y(n64930) );
  XNOR2X1 U43471 ( .A(n65278), .B(n64867), .Y(n41654) );
  XNOR2X1 U43472 ( .A(n63709), .B(n63679), .Y(n63704) );
  XNOR2X1 U43473 ( .A(n63928), .B(n41655), .Y(n64263) );
  XNOR2X1 U43474 ( .A(n64253), .B(n64252), .Y(n41655) );
  AND2X1 U43475 ( .A(n70749), .B(n70748), .Y(n41656) );
  AND2X1 U43476 ( .A(n70586), .B(n70585), .Y(n41657) );
  OR2X1 U43477 ( .A(n61824), .B(n61825), .Y(n61826) );
  AND2X1 U43478 ( .A(n70567), .B(n41658), .Y(n70263) );
  OR2X1 U43479 ( .A(n70421), .B(n70262), .Y(n41658) );
  XNOR2X1 U43480 ( .A(n41659), .B(n71235), .Y(n71606) );
  XOR2X1 U43481 ( .A(n71068), .B(n71067), .Y(n41659) );
  XOR2X1 U43482 ( .A(n71066), .B(n71368), .Y(n71067) );
  XNOR2X1 U43483 ( .A(n63544), .B(n41660), .Y(n63531) );
  XNOR2X1 U43484 ( .A(n63543), .B(n63541), .Y(n41660) );
  XOR2X1 U43485 ( .A(n71385), .B(n41661), .Y(n71622) );
  XNOR2X1 U43486 ( .A(n71475), .B(n71384), .Y(n41661) );
  AND2X1 U43487 ( .A(n69447), .B(n41662), .Y(n69456) );
  OR2X1 U43488 ( .A(n69454), .B(n69453), .Y(n41662) );
  OR2X1 U43489 ( .A(n69973), .B(n41663), .Y(n69976) );
  AND2X1 U43490 ( .A(n72510), .B(n69974), .Y(n41663) );
  XOR2X1 U43491 ( .A(n41801), .B(n64102), .Y(n63549) );
  AND2X1 U43492 ( .A(n71611), .B(n71610), .Y(n41664) );
  OR2X1 U43493 ( .A(n69804), .B(n41665), .Y(n70068) );
  AND2X1 U43494 ( .A(n69806), .B(n69805), .Y(n41665) );
  OR2X1 U43495 ( .A(n41666), .B(n70068), .Y(n70073) );
  OR2X1 U43496 ( .A(n72200), .B(n70395), .Y(n41666) );
  AND2X1 U43497 ( .A(n71258), .B(n71257), .Y(n41667) );
  AND2X1 U43498 ( .A(n72510), .B(n70931), .Y(n41668) );
  OR2X1 U43499 ( .A(n64797), .B(n41669), .Y(n64799) );
  AND2X1 U43500 ( .A(n64798), .B(n65067), .Y(n41669) );
  AND2X1 U43501 ( .A(n71238), .B(n71237), .Y(n41670) );
  XOR2X1 U43502 ( .A(n66124), .B(n41490), .Y(n41671) );
  XOR2X1 U43503 ( .A(n64772), .B(n65385), .Y(n64399) );
  AND2X1 U43504 ( .A(n71262), .B(n41672), .Y(n70928) );
  AND2X1 U43505 ( .A(n70927), .B(n43001), .Y(n41672) );
  AND2X1 U43506 ( .A(n70604), .B(n70603), .Y(n41673) );
  OR2X1 U43507 ( .A(n62010), .B(n62011), .Y(n62012) );
  AND2X1 U43508 ( .A(n62816), .B(n62815), .Y(n41674) );
  XOR2X1 U43509 ( .A(n65780), .B(n41675), .Y(n65787) );
  XOR2X1 U43510 ( .A(n71265), .B(n71280), .Y(n71271) );
  XNOR2X1 U43511 ( .A(n71277), .B(n71359), .Y(n71278) );
  OR2X1 U43512 ( .A(n62207), .B(n62208), .Y(n62209) );
  XOR2X1 U43513 ( .A(n65776), .B(n41498), .Y(n41675) );
  XOR2X1 U43514 ( .A(n72200), .B(n71578), .Y(n41676) );
  XNOR2X1 U43515 ( .A(n71996), .B(n41677), .Y(n71990) );
  XNOR2X1 U43516 ( .A(n71997), .B(n71995), .Y(n41677) );
  OR2X1 U43517 ( .A(n62656), .B(n62655), .Y(n62657) );
  AND2X1 U43518 ( .A(n43798), .B(n43862), .Y(n41678) );
  AND2X1 U43519 ( .A(n70984), .B(n70983), .Y(n41679) );
  XOR2X1 U43520 ( .A(n71998), .B(n41680), .Y(n71999) );
  XNOR2X1 U43521 ( .A(n71997), .B(n71996), .Y(n41680) );
  AND2X1 U43522 ( .A(n41681), .B(n41682), .Y(n71853) );
  NOR2X1 U43523 ( .A(n67749), .B(n67748), .Y(n41681) );
  NOR2X1 U43524 ( .A(n67754), .B(n67753), .Y(n41682) );
  XNOR2X1 U43525 ( .A(n69076), .B(n69062), .Y(n41683) );
  AND2X1 U43526 ( .A(n67430), .B(n67429), .Y(n41684) );
  XOR2X1 U43527 ( .A(n72370), .B(n72371), .Y(n41685) );
  XOR2X1 U43528 ( .A(n41862), .B(n68651), .Y(n68647) );
  XOR2X1 U43529 ( .A(n68650), .B(n72397), .Y(n41686) );
  XOR2X1 U43530 ( .A(n71573), .B(n71941), .Y(n71955) );
  XOR2X1 U43531 ( .A(n72318), .B(n71954), .Y(n41687) );
  AND2X1 U43532 ( .A(n43963), .B(n43483), .Y(n41688) );
  AND2X1 U43533 ( .A(n43952), .B(n43478), .Y(n41689) );
  XOR2X1 U43534 ( .A(n71986), .B(n72204), .Y(n72520) );
  XOR2X1 U43535 ( .A(n71833), .B(n71982), .Y(n71839) );
  XOR2X1 U43536 ( .A(n72291), .B(n69358), .Y(n41690) );
  XOR2X1 U43537 ( .A(n69775), .B(n41691), .Y(n69723) );
  XNOR2X1 U43538 ( .A(n69767), .B(n69355), .Y(n41691) );
  XNOR2X1 U43539 ( .A(n71978), .B(n71979), .Y(n71980) );
  XOR2X1 U43540 ( .A(n69760), .B(n71872), .Y(n69992) );
  XOR2X1 U43541 ( .A(n72326), .B(n70299), .Y(n41692) );
  XNOR2X1 U43542 ( .A(n41693), .B(n71013), .Y(n70646) );
  XOR2X1 U43543 ( .A(n71014), .B(n42061), .Y(n41693) );
  XNOR2X1 U43544 ( .A(n72326), .B(n71877), .Y(n41694) );
  XOR2X1 U43545 ( .A(n72355), .B(n70303), .Y(n41695) );
  XNOR2X1 U43546 ( .A(n72355), .B(n71882), .Y(n41696) );
  XOR2X1 U43547 ( .A(n72263), .B(n70995), .Y(n41697) );
  XNOR2X1 U43548 ( .A(n72509), .B(n41698), .Y(n72514) );
  XOR2X1 U43549 ( .A(n72520), .B(n72510), .Y(n41698) );
  AND2X1 U43550 ( .A(n71959), .B(n71958), .Y(n41699) );
  XOR2X1 U43551 ( .A(n71299), .B(n71300), .Y(n71009) );
  XOR2X1 U43552 ( .A(n71538), .B(n71539), .Y(n71326) );
  XNOR2X1 U43553 ( .A(n72422), .B(n71886), .Y(n41700) );
  XNOR2X1 U43554 ( .A(n72263), .B(n71889), .Y(n41701) );
  XOR2X1 U43555 ( .A(n72422), .B(n70998), .Y(n41702) );
  AND2X1 U43556 ( .A(n71893), .B(n71894), .Y(n41703) );
  XNOR2X1 U43557 ( .A(n71532), .B(n41704), .Y(n71538) );
  XNOR2X1 U43558 ( .A(n71530), .B(n71531), .Y(n41704) );
  AND2X1 U43559 ( .A(n43903), .B(n43607), .Y(n41705) );
  XOR2X1 U43560 ( .A(n71930), .B(n72486), .Y(n41706) );
  XNOR2X1 U43561 ( .A(n72221), .B(n41707), .Y(n72210) );
  XOR2X1 U43562 ( .A(n72218), .B(n72217), .Y(n41707) );
  AND2X1 U43563 ( .A(n43896), .B(n43517), .Y(n41708) );
  AND2X1 U43564 ( .A(n43896), .B(n42712), .Y(n41709) );
  AND2X1 U43565 ( .A(n71535), .B(n71534), .Y(n41710) );
  AND2X1 U43566 ( .A(n43909), .B(n43497), .Y(n41711) );
  AND2X1 U43567 ( .A(n71934), .B(n71933), .Y(n41712) );
  AND2X1 U43568 ( .A(n43909), .B(n43517), .Y(n41713) );
  AND2X1 U43569 ( .A(n43918), .B(n43501), .Y(n41714) );
  XOR2X1 U43570 ( .A(n71865), .B(n71524), .Y(n71871) );
  OR2X1 U43571 ( .A(n71899), .B(n41715), .Y(n71897) );
  OR2X1 U43572 ( .A(n72439), .B(n41516), .Y(n41715) );
  AND2X1 U43573 ( .A(n43933), .B(n43500), .Y(n41716) );
  AND2X1 U43574 ( .A(n71907), .B(n71906), .Y(n41717) );
  XOR2X1 U43575 ( .A(n71896), .B(n72436), .Y(n72448) );
  AND2X1 U43576 ( .A(n43477), .B(n43973), .Y(n41718) );
  AND2X1 U43577 ( .A(n43942), .B(n43482), .Y(n41719) );
  XOR2X1 U43578 ( .A(n71859), .B(n72298), .Y(n72289) );
  XOR2X1 U43579 ( .A(n71880), .B(n72270), .Y(n72261) );
  AND2X1 U43580 ( .A(n71863), .B(n71862), .Y(n41720) );
  AND2X1 U43581 ( .A(n71874), .B(n71873), .Y(n41721) );
  XNOR2X1 U43582 ( .A(n41722), .B(n72384), .Y(n72308) );
  XOR2X1 U43583 ( .A(n72382), .B(n72387), .Y(n41722) );
  AND2X1 U43584 ( .A(n71883), .B(n70625), .Y(n41723) );
  AND2X1 U43585 ( .A(n43477), .B(n44017), .Y(n41724) );
  XNOR2X1 U43586 ( .A(n72421), .B(n41725), .Y(n72429) );
  XOR2X1 U43587 ( .A(n72423), .B(n72422), .Y(n41725) );
  AND2X1 U43588 ( .A(n43477), .B(n44025), .Y(n41726) );
  AND2X1 U43589 ( .A(n43796), .B(n44055), .Y(n41727) );
  AND2X1 U43590 ( .A(n43799), .B(n44055), .Y(n41728) );
  AND2X1 U43591 ( .A(n42711), .B(n44055), .Y(n41729) );
  AND2X1 U43592 ( .A(n43483), .B(n44055), .Y(n41730) );
  AND2X1 U43593 ( .A(n43477), .B(n44055), .Y(n41731) );
  AND2X1 U43594 ( .A(n57673), .B(n57672), .Y(n41732) );
  AND2X1 U43595 ( .A(n38311), .B(n44055), .Y(n41733) );
  XOR2X1 U43596 ( .A(n72510), .B(n72200), .Y(n41734) );
  AND2X1 U43597 ( .A(n43500), .B(n44047), .Y(n41735) );
  AND2X1 U43598 ( .A(n57801), .B(n57809), .Y(n57802) );
  AND2X1 U43599 ( .A(n43496), .B(n44054), .Y(n41736) );
  AND2X1 U43600 ( .A(n43518), .B(n44054), .Y(n41737) );
  AND2X1 U43601 ( .A(n73172), .B(n73503), .Y(n41738) );
  XOR2X1 U43602 ( .A(n60201), .B(n39900), .Y(n41739) );
  AND2X1 U43603 ( .A(n38604), .B(n46906), .Y(n41740) );
  AND2X1 U43604 ( .A(n40499), .B(n40035), .Y(n41741) );
  AND2X1 U43605 ( .A(n40499), .B(n46979), .Y(n41742) );
  OR2X1 U43606 ( .A(n59394), .B(n59395), .Y(n59396) );
  OR2X1 U43607 ( .A(n59173), .B(n59174), .Y(n59175) );
  OR2X1 U43608 ( .A(n59199), .B(n59198), .Y(n59200) );
  OR2X1 U43609 ( .A(n59209), .B(n41743), .Y(n59183) );
  AND2X1 U43610 ( .A(n39051), .B(n59181), .Y(n41743) );
  OR2X1 U43611 ( .A(n41744), .B(n41745), .Y(n63481) );
  AND2X1 U43612 ( .A(n63344), .B(n63343), .Y(n41744) );
  AND2X1 U43613 ( .A(n42182), .B(n63351), .Y(n41745) );
  AND2X1 U43614 ( .A(n63876), .B(n41746), .Y(n63874) );
  INVX1 U43615 ( .A(n63872), .Y(n41746) );
  AND2X1 U43616 ( .A(n41747), .B(n41748), .Y(n42829) );
  NAND2X1 U43617 ( .A(n40288), .B(n59332), .Y(n41747) );
  NAND2X1 U43618 ( .A(n59317), .B(n59316), .Y(n41748) );
  AND2X1 U43619 ( .A(n60240), .B(n63824), .Y(n41749) );
  OR2X1 U43620 ( .A(n60231), .B(n60232), .Y(n60937) );
  XNOR2X1 U43621 ( .A(n41750), .B(n59265), .Y(n59330) );
  XOR2X1 U43622 ( .A(n59270), .B(n59266), .Y(n41750) );
  XOR2X1 U43623 ( .A(n62404), .B(n62393), .Y(n61238) );
  AND2X1 U43624 ( .A(n43456), .B(n42709), .Y(n41751) );
  XNOR2X1 U43625 ( .A(n60637), .B(n41752), .Y(n60648) );
  XNOR2X1 U43626 ( .A(n60631), .B(n60250), .Y(n41752) );
  NAND2X1 U43627 ( .A(n62659), .B(n72811), .Y(n59245) );
  OR2X1 U43628 ( .A(n60598), .B(n60599), .Y(n60935) );
  XNOR2X1 U43629 ( .A(n61137), .B(n41753), .Y(n61205) );
  XNOR2X1 U43630 ( .A(n61136), .B(n60973), .Y(n41753) );
  XNOR2X1 U43631 ( .A(n64487), .B(n41754), .Y(n64346) );
  XNOR2X1 U43632 ( .A(n64486), .B(n64488), .Y(n41754) );
  OR2X1 U43633 ( .A(n41755), .B(n41756), .Y(n66203) );
  AND2X1 U43634 ( .A(n65664), .B(n65663), .Y(n41755) );
  AND2X1 U43635 ( .A(n65674), .B(n65673), .Y(n41756) );
  XNOR2X1 U43636 ( .A(n66203), .B(n41757), .Y(n66023) );
  XNOR2X1 U43637 ( .A(n66201), .B(n66204), .Y(n41757) );
  AND2X1 U43638 ( .A(n41758), .B(n66001), .Y(n66004) );
  OR2X1 U43639 ( .A(n65999), .B(n66000), .Y(n41758) );
  AND2X1 U43640 ( .A(n40471), .B(n43456), .Y(n41759) );
  AND2X1 U43641 ( .A(n43456), .B(n40482), .Y(n41760) );
  XOR2X1 U43642 ( .A(n40614), .B(n60631), .Y(n60638) );
  AND2X1 U43643 ( .A(n43458), .B(n40462), .Y(n41761) );
  AND2X1 U43644 ( .A(n66668), .B(n41762), .Y(n66307) );
  INVX1 U43645 ( .A(n66659), .Y(n41762) );
  AND2X1 U43646 ( .A(n66310), .B(n66665), .Y(n41763) );
  XNOR2X1 U43647 ( .A(n41764), .B(n66308), .Y(n66646) );
  XOR2X1 U43648 ( .A(n66659), .B(n66309), .Y(n41764) );
  XNOR2X1 U43649 ( .A(n40218), .B(n41765), .Y(n63888) );
  XNOR2X1 U43650 ( .A(n63875), .B(n63872), .Y(n41765) );
  AND2X1 U43651 ( .A(n40152), .B(n46019), .Y(n45453) );
  XOR2X1 U43652 ( .A(n38098), .B(n61136), .Y(n61140) );
  NOR2X1 U43653 ( .A(n41767), .B(n41768), .Y(n41766) );
  AND2X1 U43654 ( .A(n70108), .B(n40670), .Y(n41767) );
  AND2X1 U43655 ( .A(n70255), .B(n70254), .Y(n41768) );
  AND2X1 U43656 ( .A(n43458), .B(n72820), .Y(n41769) );
  AND2X1 U43657 ( .A(n43464), .B(n43502), .Y(n41770) );
  XNOR2X1 U43658 ( .A(n67508), .B(n41771), .Y(n66997) );
  XOR2X1 U43659 ( .A(n67506), .B(n66846), .Y(n41771) );
  AND2X1 U43660 ( .A(n43819), .B(n43456), .Y(n41772) );
  AND2X1 U43661 ( .A(n40392), .B(n43787), .Y(n41773) );
  AND2X1 U43662 ( .A(n43472), .B(n40484), .Y(n41774) );
  AND2X1 U43663 ( .A(n43458), .B(n43757), .Y(n41775) );
  AND2X1 U43664 ( .A(n43458), .B(n72760), .Y(n41776) );
  AND2X1 U43665 ( .A(n69634), .B(n41777), .Y(n69489) );
  AND2X1 U43666 ( .A(n69633), .B(n40683), .Y(n41777) );
  AND2X1 U43667 ( .A(n40472), .B(n40392), .Y(n41778) );
  AND2X1 U43668 ( .A(n43465), .B(n43795), .Y(n41779) );
  AND2X1 U43669 ( .A(n40393), .B(n40465), .Y(n41780) );
  AND2X1 U43670 ( .A(n43458), .B(n39164), .Y(n41781) );
  XNOR2X1 U43671 ( .A(n66832), .B(n66470), .Y(n66640) );
  XOR2X1 U43672 ( .A(n42183), .B(n67313), .Y(n67163) );
  XOR2X1 U43673 ( .A(n62949), .B(n63236), .Y(n63249) );
  AND2X1 U43674 ( .A(n39810), .B(n43017), .Y(n41782) );
  AND2X1 U43675 ( .A(n38364), .B(n43017), .Y(n41783) );
  AND2X1 U43676 ( .A(n71371), .B(n71370), .Y(n41784) );
  AND2X1 U43677 ( .A(n40392), .B(n43810), .Y(n41785) );
  XOR2X1 U43678 ( .A(n63234), .B(n63812), .Y(n63544) );
  NOR2X1 U43679 ( .A(n41787), .B(n42672), .Y(n41786) );
  INVX1 U43680 ( .A(n39810), .Y(n41787) );
  AND2X1 U43681 ( .A(n63229), .B(n41788), .Y(n63233) );
  OR2X1 U43682 ( .A(n38514), .B(n63230), .Y(n41788) );
  AND2X1 U43683 ( .A(n43456), .B(n43743), .Y(n41789) );
  AND2X1 U43684 ( .A(n43456), .B(n72810), .Y(n41790) );
  AND2X1 U43685 ( .A(n39810), .B(n42756), .Y(n41791) );
  AND2X1 U43686 ( .A(n43820), .B(n43471), .Y(n41792) );
  AND2X1 U43687 ( .A(n40392), .B(n43759), .Y(n41793) );
  AND2X1 U43688 ( .A(n40473), .B(n43465), .Y(n41794) );
  AND2X1 U43689 ( .A(n43465), .B(n43787), .Y(n41795) );
  AND2X1 U43690 ( .A(n40393), .B(n43737), .Y(n41796) );
  AND2X1 U43691 ( .A(n43465), .B(n40485), .Y(n41797) );
  AND2X1 U43692 ( .A(n43464), .B(n40463), .Y(n41798) );
  AND2X1 U43693 ( .A(n40393), .B(n39163), .Y(n41799) );
  AND2X1 U43694 ( .A(n71242), .B(n71241), .Y(n41800) );
  AND2X1 U43695 ( .A(n63218), .B(n63217), .Y(n41801) );
  XOR2X1 U43696 ( .A(n63811), .B(n63574), .Y(n63809) );
  AND2X1 U43697 ( .A(n64098), .B(n64097), .Y(n41802) );
  AND2X1 U43698 ( .A(n39082), .B(n64079), .Y(n41803) );
  AND2X1 U43699 ( .A(n43456), .B(n39525), .Y(n41804) );
  XNOR2X1 U43700 ( .A(n64106), .B(n64777), .Y(n41805) );
  AND2X1 U43701 ( .A(n43471), .B(n43791), .Y(n41806) );
  AND2X1 U43702 ( .A(n43464), .B(n72820), .Y(n41807) );
  AND2X1 U43703 ( .A(n39937), .B(n43787), .Y(n41808) );
  AND2X1 U43704 ( .A(n40473), .B(n39943), .Y(n41809) );
  AND2X1 U43705 ( .A(n43472), .B(n43743), .Y(n41810) );
  AND2X1 U43706 ( .A(n43820), .B(n43466), .Y(n41811) );
  AND2X1 U43707 ( .A(n39942), .B(n40486), .Y(n41812) );
  AND2X1 U43708 ( .A(n43464), .B(n43759), .Y(n41813) );
  AND2X1 U43709 ( .A(n43464), .B(n43737), .Y(n41814) );
  AND2X1 U43710 ( .A(n39938), .B(n40464), .Y(n41815) );
  AND2X1 U43711 ( .A(n43464), .B(n43781), .Y(n41816) );
  AND2X1 U43712 ( .A(n43471), .B(n39525), .Y(n41817) );
  AND2X1 U43713 ( .A(n43464), .B(n43791), .Y(n41818) );
  XOR2X1 U43714 ( .A(n65077), .B(n65078), .Y(n65385) );
  AND2X1 U43715 ( .A(n39940), .B(n43810), .Y(n41819) );
  AND2X1 U43716 ( .A(n43802), .B(n43458), .Y(n41820) );
  AND2X1 U43717 ( .A(n71276), .B(n71275), .Y(n41821) );
  AND2X1 U43718 ( .A(n43464), .B(n43743), .Y(n41822) );
  AND2X1 U43719 ( .A(n71283), .B(n71282), .Y(n41823) );
  AND2X1 U43720 ( .A(n43820), .B(n39939), .Y(n41824) );
  AND2X1 U43721 ( .A(n39941), .B(n43759), .Y(n41825) );
  XNOR2X1 U43722 ( .A(n71359), .B(n41826), .Y(n71265) );
  XOR2X1 U43723 ( .A(n72202), .B(n71277), .Y(n41826) );
  AND2X1 U43724 ( .A(n43840), .B(n40487), .Y(n41827) );
  AND2X1 U43725 ( .A(n40474), .B(n43842), .Y(n41828) );
  AND2X1 U43726 ( .A(n39937), .B(n43737), .Y(n41829) );
  AND2X1 U43727 ( .A(n43840), .B(n40464), .Y(n41830) );
  AND2X1 U43728 ( .A(n39943), .B(n43780), .Y(n41831) );
  XNOR2X1 U43729 ( .A(n65774), .B(n65386), .Y(n65776) );
  AND2X1 U43730 ( .A(n71362), .B(n71361), .Y(n41832) );
  AND2X1 U43731 ( .A(n71355), .B(n71354), .Y(n41833) );
  AND2X1 U43732 ( .A(n43791), .B(n39942), .Y(n41834) );
  AND2X1 U43733 ( .A(n43840), .B(n72820), .Y(n41835) );
  AND2X1 U43734 ( .A(n43802), .B(n40393), .Y(n41836) );
  AND2X1 U43735 ( .A(n43742), .B(n39943), .Y(n41837) );
  AND2X1 U43736 ( .A(n43820), .B(n43842), .Y(n41838) );
  AND2X1 U43737 ( .A(n40475), .B(n38382), .Y(n41839) );
  AND2X1 U43738 ( .A(n43841), .B(n43758), .Y(n41840) );
  AND2X1 U43739 ( .A(n43841), .B(n43737), .Y(n41841) );
  AND2X1 U43740 ( .A(n38383), .B(n40488), .Y(n41842) );
  AND2X1 U43741 ( .A(n38381), .B(n40465), .Y(n41843) );
  AND2X1 U43742 ( .A(n43841), .B(n39164), .Y(n41844) );
  AND2X1 U43743 ( .A(n43764), .B(n39938), .Y(n41845) );
  AND2X1 U43744 ( .A(n43750), .B(n43456), .Y(n41846) );
  AND2X1 U43745 ( .A(n38379), .B(n43810), .Y(n41847) );
  AND2X1 U43746 ( .A(n40392), .B(n43814), .Y(n41848) );
  AND2X1 U43747 ( .A(n40476), .B(n44038), .Y(n41849) );
  AND2X1 U43748 ( .A(n38582), .B(n43466), .Y(n41850) );
  AND2X1 U43749 ( .A(n43821), .B(n38384), .Y(n41851) );
  AND2X1 U43750 ( .A(n43841), .B(n43742), .Y(n41852) );
  AND2X1 U43751 ( .A(n71844), .B(n72366), .Y(n41853) );
  AND2X1 U43752 ( .A(n44035), .B(n40489), .Y(n41854) );
  AND2X1 U43753 ( .A(n38381), .B(n43758), .Y(n41855) );
  AND2X1 U43754 ( .A(n43736), .B(n38382), .Y(n41856) );
  AND2X1 U43755 ( .A(n43779), .B(n38380), .Y(n41857) );
  AND2X1 U43756 ( .A(n44036), .B(n40466), .Y(n41858) );
  XNOR2X1 U43757 ( .A(n71504), .B(n41859), .Y(n71494) );
  XOR2X1 U43758 ( .A(n72225), .B(n71503), .Y(n41859) );
  AND2X1 U43759 ( .A(n43472), .B(n43752), .Y(n41860) );
  AND2X1 U43760 ( .A(n43764), .B(n43842), .Y(n41861) );
  XOR2X1 U43761 ( .A(n68376), .B(n68649), .Y(n41862) );
  AND2X1 U43762 ( .A(n43792), .B(n38383), .Y(n41863) );
  AND2X1 U43763 ( .A(n43815), .B(n43466), .Y(n41864) );
  AND2X1 U43764 ( .A(n38582), .B(n39939), .Y(n41865) );
  AND2X1 U43765 ( .A(n43731), .B(n43458), .Y(n41866) );
  AND2X1 U43766 ( .A(n43742), .B(n38384), .Y(n41867) );
  AND2X1 U43767 ( .A(n44035), .B(n43758), .Y(n41868) );
  AND2X1 U43768 ( .A(n43850), .B(n40467), .Y(n41869) );
  AND2X1 U43769 ( .A(n44035), .B(n39163), .Y(n41870) );
  AND2X1 U43770 ( .A(n43764), .B(n38378), .Y(n41871) );
  AND2X1 U43771 ( .A(n43750), .B(n43466), .Y(n41872) );
  AND2X1 U43772 ( .A(n43792), .B(n44037), .Y(n41873) );
  AND2X1 U43773 ( .A(n43816), .B(n39940), .Y(n41874) );
  AND2X1 U43774 ( .A(n38582), .B(n43842), .Y(n41875) );
  AND2X1 U43775 ( .A(n43471), .B(n43731), .Y(n41876) );
  AND2X1 U43776 ( .A(n43742), .B(n44037), .Y(n41877) );
  AND2X1 U43777 ( .A(n43850), .B(n43758), .Y(n41878) );
  AND2X1 U43778 ( .A(n43736), .B(n43852), .Y(n41879) );
  AND2X1 U43779 ( .A(n71843), .B(n72372), .Y(n41880) );
  AND2X1 U43780 ( .A(n43781), .B(n43852), .Y(n41881) );
  AND2X1 U43781 ( .A(n43764), .B(n44037), .Y(n41882) );
  AND2X1 U43782 ( .A(n43750), .B(n39941), .Y(n41883) );
  AND2X1 U43783 ( .A(n43792), .B(n43852), .Y(n41884) );
  AND2X1 U43784 ( .A(n43816), .B(n43842), .Y(n41885) );
  AND2X1 U43785 ( .A(n43803), .B(n38379), .Y(n41886) );
  AND2X1 U43786 ( .A(n43730), .B(n43466), .Y(n41887) );
  AND2X1 U43787 ( .A(n43742), .B(n43852), .Y(n41888) );
  AND2X1 U43788 ( .A(n43859), .B(n43736), .Y(n41889) );
  AND2X1 U43789 ( .A(n43860), .B(n39164), .Y(n41890) );
  AND2X1 U43790 ( .A(n43764), .B(n43852), .Y(n41891) );
  AND2X1 U43791 ( .A(n43750), .B(n43842), .Y(n41892) );
  AND2X1 U43792 ( .A(n43859), .B(n43792), .Y(n41893) );
  AND2X1 U43793 ( .A(n43821), .B(n43964), .Y(n41894) );
  AND2X1 U43794 ( .A(n43809), .B(n43965), .Y(n41895) );
  AND2X1 U43795 ( .A(n43816), .B(n38380), .Y(n41896) );
  AND2X1 U43796 ( .A(n43803), .B(n44037), .Y(n41897) );
  AND2X1 U43797 ( .A(n43730), .B(n39942), .Y(n41898) );
  AND2X1 U43798 ( .A(n43860), .B(n38611), .Y(n41899) );
  AND2X1 U43799 ( .A(n72387), .B(n72310), .Y(n41900) );
  AND2X1 U43800 ( .A(n43736), .B(n43964), .Y(n41901) );
  XOR2X1 U43801 ( .A(n71305), .B(n70999), .Y(n71314) );
  XOR2X1 U43802 ( .A(n71004), .B(n71315), .Y(n71300) );
  AND2X1 U43803 ( .A(n39163), .B(n43964), .Y(n41902) );
  AND2X1 U43804 ( .A(n43860), .B(n39525), .Y(n41903) );
  AND2X1 U43805 ( .A(n43750), .B(n38381), .Y(n41904) );
  AND2X1 U43806 ( .A(n43792), .B(n43964), .Y(n41905) );
  AND2X1 U43807 ( .A(n43816), .B(n44037), .Y(n41906) );
  AND2X1 U43808 ( .A(n43803), .B(n43852), .Y(n41907) );
  AND2X1 U43809 ( .A(n43730), .B(n43841), .Y(n41908) );
  XOR2X1 U43810 ( .A(n71516), .B(n71313), .Y(n71511) );
  XOR2X1 U43811 ( .A(n71318), .B(n71512), .Y(n71531) );
  AND2X1 U43812 ( .A(n43742), .B(n43964), .Y(n41909) );
  AND2X1 U43813 ( .A(n43821), .B(n43954), .Y(n41910) );
  AND2X1 U43814 ( .A(n43758), .B(n43954), .Y(n41911) );
  AND2X1 U43815 ( .A(n43736), .B(n43954), .Y(n41912) );
  AND2X1 U43816 ( .A(n43781), .B(n43954), .Y(n41913) );
  AND2X1 U43817 ( .A(n43764), .B(n43964), .Y(n41914) );
  AND2X1 U43818 ( .A(n43750), .B(n44037), .Y(n41915) );
  AND2X1 U43819 ( .A(n43792), .B(n43954), .Y(n41916) );
  AND2X1 U43820 ( .A(n43816), .B(n43852), .Y(n41917) );
  AND2X1 U43821 ( .A(n43730), .B(n38382), .Y(n41918) );
  AND2X1 U43822 ( .A(n43860), .B(n43804), .Y(n41919) );
  AND2X1 U43823 ( .A(n43742), .B(n43954), .Y(n41920) );
  AND2X1 U43824 ( .A(n43869), .B(n43780), .Y(n41921) );
  AND2X1 U43825 ( .A(n43909), .B(n43724), .Y(n41922) );
  AND2X1 U43826 ( .A(n72820), .B(n43881), .Y(n41923) );
  AND2X1 U43827 ( .A(n43764), .B(n43954), .Y(n41924) );
  AND2X1 U43828 ( .A(n43750), .B(n43852), .Y(n41925) );
  AND2X1 U43829 ( .A(n43870), .B(n43792), .Y(n41926) );
  AND2X1 U43830 ( .A(n43860), .B(n43816), .Y(n41927) );
  AND2X1 U43831 ( .A(n43730), .B(n44037), .Y(n41928) );
  AND2X1 U43832 ( .A(n43803), .B(n43964), .Y(n41929) );
  AND2X1 U43833 ( .A(n43897), .B(n43788), .Y(n41930) );
  AND2X1 U43834 ( .A(n43870), .B(n43742), .Y(n41931) );
  AND2X1 U43835 ( .A(n39164), .B(n43881), .Y(n41932) );
  AND2X1 U43836 ( .A(n43870), .B(n39525), .Y(n41933) );
  AND2X1 U43837 ( .A(n43860), .B(n43752), .Y(n41934) );
  XOR2X1 U43838 ( .A(n41935), .B(n71529), .Y(n71904) );
  NOR2X1 U43839 ( .A(n71519), .B(n71518), .Y(n41935) );
  AND2X1 U43840 ( .A(n43792), .B(n43881), .Y(n41936) );
  AND2X1 U43841 ( .A(n43816), .B(n43963), .Y(n41937) );
  AND2X1 U43842 ( .A(n43758), .B(n43891), .Y(n41938) );
  AND2X1 U43843 ( .A(n43803), .B(n43954), .Y(n41939) );
  AND2X1 U43844 ( .A(n43730), .B(n43851), .Y(n41940) );
  AND2X1 U43845 ( .A(n43742), .B(n43881), .Y(n41941) );
  AND2X1 U43846 ( .A(n43736), .B(n43891), .Y(n41942) );
  AND2X1 U43847 ( .A(n39163), .B(n43891), .Y(n41943) );
  AND2X1 U43848 ( .A(n43898), .B(n40463), .Y(n41944) );
  AND2X1 U43849 ( .A(n43764), .B(n43881), .Y(n41945) );
  AND2X1 U43850 ( .A(n43751), .B(n43963), .Y(n41946) );
  AND2X1 U43851 ( .A(n43897), .B(n43758), .Y(n41947) );
  AND2X1 U43852 ( .A(n43792), .B(n43891), .Y(n41948) );
  AND2X1 U43853 ( .A(n43816), .B(n43954), .Y(n41949) );
  AND2X1 U43854 ( .A(n43860), .B(n43731), .Y(n41950) );
  AND2X1 U43855 ( .A(n43870), .B(n43804), .Y(n41951) );
  AND2X1 U43856 ( .A(n43741), .B(n43891), .Y(n41952) );
  AND2X1 U43857 ( .A(n43897), .B(n43781), .Y(n41953) );
  AND2X1 U43858 ( .A(n43764), .B(n43891), .Y(n41954) );
  AND2X1 U43859 ( .A(n43750), .B(n43953), .Y(n41955) );
  XOR2X1 U43860 ( .A(n71871), .B(n71525), .Y(n71876) );
  AND2X1 U43861 ( .A(n43897), .B(n43792), .Y(n41956) );
  AND2X1 U43862 ( .A(n43821), .B(n43905), .Y(n41957) );
  AND2X1 U43863 ( .A(n43870), .B(n43816), .Y(n41958) );
  AND2X1 U43864 ( .A(n43730), .B(n43963), .Y(n41959) );
  AND2X1 U43865 ( .A(n43803), .B(n43881), .Y(n41960) );
  AND2X1 U43866 ( .A(n43897), .B(n43742), .Y(n41961) );
  AND2X1 U43867 ( .A(n43780), .B(n43905), .Y(n41962) );
  AND2X1 U43868 ( .A(n43897), .B(n39525), .Y(n41963) );
  AND2X1 U43869 ( .A(n43870), .B(n43752), .Y(n41964) );
  AND2X1 U43870 ( .A(n43792), .B(n43905), .Y(n41965) );
  AND2X1 U43871 ( .A(n43919), .B(n40482), .Y(n41966) );
  AND2X1 U43872 ( .A(n43788), .B(n43934), .Y(n41967) );
  AND2X1 U43873 ( .A(n43816), .B(n43881), .Y(n41968) );
  AND2X1 U43874 ( .A(n43730), .B(n43953), .Y(n41969) );
  AND2X1 U43875 ( .A(n43803), .B(n43891), .Y(n41970) );
  AND2X1 U43876 ( .A(n43741), .B(n43905), .Y(n41971) );
  AND2X1 U43877 ( .A(n43910), .B(n39164), .Y(n41972) );
  AND2X1 U43878 ( .A(n43724), .B(n43973), .Y(n41973) );
  AND2X1 U43879 ( .A(n43763), .B(n43905), .Y(n41974) );
  AND2X1 U43880 ( .A(n43751), .B(n43880), .Y(n41975) );
  AND2X1 U43881 ( .A(n43910), .B(n43792), .Y(n41976) );
  AND2X1 U43882 ( .A(n43920), .B(n43821), .Y(n41977) );
  AND2X1 U43883 ( .A(n43816), .B(n43891), .Y(n41978) );
  AND2X1 U43884 ( .A(n43871), .B(n43731), .Y(n41979) );
  AND2X1 U43885 ( .A(n43897), .B(n43804), .Y(n41980) );
  AND2X1 U43886 ( .A(n43910), .B(n38611), .Y(n41981) );
  AND2X1 U43887 ( .A(n43920), .B(n39163), .Y(n41982) );
  AND2X1 U43888 ( .A(n40470), .B(n43935), .Y(n41983) );
  AND2X1 U43889 ( .A(n43910), .B(n39525), .Y(n41984) );
  AND2X1 U43890 ( .A(n43751), .B(n43891), .Y(n41985) );
  AND2X1 U43891 ( .A(n43919), .B(n43792), .Y(n41986) );
  AND2X1 U43892 ( .A(n43897), .B(n43816), .Y(n41987) );
  AND2X1 U43893 ( .A(n43730), .B(n43880), .Y(n41988) );
  AND2X1 U43894 ( .A(n43803), .B(n43905), .Y(n41989) );
  AND2X1 U43895 ( .A(n43919), .B(n38611), .Y(n41990) );
  AND2X1 U43896 ( .A(n43926), .B(n43737), .Y(n41991) );
  AND2X1 U43897 ( .A(n40473), .B(n43943), .Y(n41992) );
  AND2X1 U43898 ( .A(n43926), .B(n39163), .Y(n41993) );
  AND2X1 U43899 ( .A(n40468), .B(n43944), .Y(n41994) );
  AND2X1 U43900 ( .A(n43919), .B(n39525), .Y(n41995) );
  AND2X1 U43901 ( .A(n43897), .B(n43752), .Y(n41996) );
  AND2X1 U43902 ( .A(n43926), .B(n43792), .Y(n41997) );
  AND2X1 U43903 ( .A(n40474), .B(n43974), .Y(n41998) );
  AND2X1 U43904 ( .A(n43788), .B(n43983), .Y(n41999) );
  AND2X1 U43905 ( .A(n43816), .B(n43904), .Y(n42000) );
  AND2X1 U43906 ( .A(n43730), .B(n43890), .Y(n42001) );
  AND2X1 U43907 ( .A(n43910), .B(n43804), .Y(n42002) );
  AND2X1 U43908 ( .A(n43927), .B(n38611), .Y(n42003) );
  AND2X1 U43909 ( .A(n40488), .B(n43984), .Y(n42004) );
  AND2X1 U43910 ( .A(n43788), .B(n43992), .Y(n42005) );
  AND2X1 U43911 ( .A(n43735), .B(n43936), .Y(n42006) );
  AND2X1 U43912 ( .A(n43779), .B(n43935), .Y(n42007) );
  AND2X1 U43913 ( .A(n43926), .B(n39525), .Y(n42008) );
  AND2X1 U43914 ( .A(n43751), .B(n43904), .Y(n42009) );
  AND2X1 U43915 ( .A(n43792), .B(n43935), .Y(n42010) );
  AND2X1 U43916 ( .A(n43910), .B(n43816), .Y(n42011) );
  AND2X1 U43917 ( .A(n43896), .B(n43731), .Y(n42012) );
  AND2X1 U43918 ( .A(n43919), .B(n43804), .Y(n42013) );
  AND2X1 U43919 ( .A(n43741), .B(n43935), .Y(n42014) );
  AND2X1 U43920 ( .A(n43735), .B(n43945), .Y(n42015) );
  AND2X1 U43921 ( .A(n43779), .B(n43944), .Y(n42016) );
  AND2X1 U43922 ( .A(n43910), .B(n43752), .Y(n42017) );
  AND2X1 U43923 ( .A(n43763), .B(n43935), .Y(n42018) );
  AND2X1 U43924 ( .A(n43792), .B(n43944), .Y(n42019) );
  AND2X1 U43925 ( .A(n40461), .B(n43993), .Y(n42020) );
  AND2X1 U43926 ( .A(n43919), .B(n43816), .Y(n42021) );
  AND2X1 U43927 ( .A(n43730), .B(n43904), .Y(n42022) );
  AND2X1 U43928 ( .A(n43927), .B(n43804), .Y(n42023) );
  AND2X1 U43929 ( .A(n43741), .B(n43944), .Y(n42024) );
  AND2X1 U43930 ( .A(n43735), .B(n43975), .Y(n42025) );
  AND2X1 U43931 ( .A(n43477), .B(n44008), .Y(n42026) );
  AND2X1 U43932 ( .A(n43779), .B(n43975), .Y(n42027) );
  AND2X1 U43933 ( .A(n43758), .B(n43984), .Y(n42028) );
  AND2X1 U43934 ( .A(n43919), .B(n43752), .Y(n42029) );
  AND2X1 U43935 ( .A(n43763), .B(n43944), .Y(n42030) );
  AND2X1 U43936 ( .A(n43792), .B(n43974), .Y(n42031) );
  AND2X1 U43937 ( .A(n43821), .B(n43993), .Y(n42032) );
  AND2X1 U43938 ( .A(n44007), .B(n43496), .Y(n42033) );
  AND2X1 U43939 ( .A(n43774), .B(n44008), .Y(n42034) );
  AND2X1 U43940 ( .A(n43927), .B(n43816), .Y(n42035) );
  AND2X1 U43941 ( .A(n43910), .B(n43731), .Y(n42036) );
  AND2X1 U43942 ( .A(n43804), .B(n43935), .Y(n42037) );
  AND2X1 U43943 ( .A(n43741), .B(n43974), .Y(n42038) );
  AND2X1 U43944 ( .A(n43779), .B(n43985), .Y(n42039) );
  AND2X1 U43945 ( .A(n43809), .B(n44009), .Y(n42040) );
  AND2X1 U43946 ( .A(n43926), .B(n43752), .Y(n42041) );
  AND2X1 U43947 ( .A(n43763), .B(n43974), .Y(n42042) );
  AND2X1 U43948 ( .A(n43792), .B(n43985), .Y(n42043) );
  AND2X1 U43949 ( .A(n40461), .B(n44009), .Y(n42044) );
  OR2X1 U43950 ( .A(n49805), .B(n43494), .Y(n49873) );
  OR2X1 U43951 ( .A(n42045), .B(n31152), .Y(n49802) );
  AND2X1 U43952 ( .A(n49800), .B(n49799), .Y(n42045) );
  AND2X1 U43953 ( .A(n42186), .B(n57632), .Y(n42046) );
  AND2X1 U43954 ( .A(n43809), .B(n44018), .Y(n42047) );
  AND2X1 U43955 ( .A(n43816), .B(n43935), .Y(n42048) );
  AND2X1 U43956 ( .A(n43919), .B(n43731), .Y(n42049) );
  AND2X1 U43957 ( .A(n43804), .B(n43944), .Y(n42050) );
  AND2X1 U43958 ( .A(n43741), .B(n43985), .Y(n42051) );
  AND2X1 U43959 ( .A(n43779), .B(n43994), .Y(n42052) );
  AND2X1 U43960 ( .A(n43792), .B(n43994), .Y(n42053) );
  AND2X1 U43961 ( .A(n43763), .B(n43984), .Y(n42054) );
  AND2X1 U43962 ( .A(n43751), .B(n43935), .Y(n42055) );
  AND2X1 U43963 ( .A(n44007), .B(n43607), .Y(n42056) );
  AND2X1 U43964 ( .A(n40465), .B(n44056), .Y(n42057) );
  AND2X1 U43965 ( .A(n43816), .B(n43944), .Y(n42058) );
  AND2X1 U43966 ( .A(n43926), .B(n43731), .Y(n42059) );
  AND2X1 U43967 ( .A(n43803), .B(n43974), .Y(n42060) );
  AND2X1 U43968 ( .A(n44007), .B(n43518), .Y(n42061) );
  AND2X1 U43969 ( .A(n43779), .B(n44001), .Y(n42062) );
  AND2X1 U43970 ( .A(n43741), .B(n43994), .Y(n42063) );
  AND2X1 U43971 ( .A(n43792), .B(n44002), .Y(n42064) );
  AND2X1 U43972 ( .A(n43763), .B(n43994), .Y(n42065) );
  AND2X1 U43973 ( .A(n43751), .B(n43944), .Y(n42066) );
  AND2X1 U43974 ( .A(n43809), .B(n44049), .Y(n42067) );
  AND2X1 U43975 ( .A(n57640), .B(n48689), .Y(n42068) );
  AND2X1 U43976 ( .A(n48827), .B(n48826), .Y(n42069) );
  AND2X1 U43977 ( .A(n43729), .B(n43935), .Y(n42070) );
  AND2X1 U43978 ( .A(n43816), .B(n43974), .Y(n42071) );
  AND2X1 U43979 ( .A(n43803), .B(n43984), .Y(n42072) );
  AND2X1 U43980 ( .A(n43779), .B(n44009), .Y(n42073) );
  AND2X1 U43981 ( .A(n43741), .B(n44002), .Y(n42074) );
  AND2X1 U43982 ( .A(n43792), .B(n44009), .Y(n42075) );
  AND2X1 U43983 ( .A(n43763), .B(n44002), .Y(n42076) );
  AND2X1 U43984 ( .A(n43751), .B(n43974), .Y(n42077) );
  AND2X1 U43985 ( .A(n43779), .B(n44018), .Y(n42078) );
  AND2X1 U43986 ( .A(n43729), .B(n43944), .Y(n42079) );
  AND2X1 U43987 ( .A(n43816), .B(n43984), .Y(n42080) );
  AND2X1 U43988 ( .A(n43803), .B(n43994), .Y(n42081) );
  AND2X1 U43989 ( .A(n43742), .B(n44010), .Y(n42082) );
  AND2X1 U43990 ( .A(n43735), .B(n44026), .Y(n42083) );
  AND2X1 U43991 ( .A(n49234), .B(n49233), .Y(n42084) );
  AND2X1 U43992 ( .A(n43792), .B(n44018), .Y(n42085) );
  AND2X1 U43993 ( .A(n43763), .B(n44010), .Y(n42086) );
  AND2X1 U43994 ( .A(n43750), .B(n43984), .Y(n42087) );
  AND2X1 U43995 ( .A(n43779), .B(n44049), .Y(n42088) );
  AND2X1 U43996 ( .A(n43729), .B(n43974), .Y(n42089) );
  AND2X1 U43997 ( .A(n43816), .B(n43994), .Y(n42090) );
  AND2X1 U43998 ( .A(n57766), .B(n42091), .Y(n57767) );
  OR2X1 U43999 ( .A(n39944), .B(n43744), .Y(n42091) );
  AND2X1 U44000 ( .A(n43803), .B(n44002), .Y(n42092) );
  AND2X1 U44001 ( .A(n43741), .B(n44019), .Y(n42093) );
  AND2X1 U44002 ( .A(n43792), .B(n44026), .Y(n42094) );
  AND2X1 U44003 ( .A(n43764), .B(n44019), .Y(n42095) );
  AND2X1 U44004 ( .A(n43751), .B(n43993), .Y(n42096) );
  AND2X1 U44005 ( .A(n43729), .B(n43984), .Y(n42097) );
  AND2X1 U44006 ( .A(n43816), .B(n44002), .Y(n42098) );
  AND2X1 U44007 ( .A(n38582), .B(n44010), .Y(n42099) );
  AND2X1 U44008 ( .A(n43741), .B(n44026), .Y(n42100) );
  AND2X1 U44009 ( .A(n43763), .B(n44027), .Y(n42101) );
  AND2X1 U44010 ( .A(n43751), .B(n44002), .Y(n42102) );
  AND2X1 U44011 ( .A(n43729), .B(n43993), .Y(n42103) );
  AND2X1 U44012 ( .A(n43816), .B(n44009), .Y(n42104) );
  AND2X1 U44013 ( .A(n38582), .B(n44019), .Y(n42105) );
  AND2X1 U44014 ( .A(n43741), .B(n44049), .Y(n42106) );
  XOR2X1 U44015 ( .A(n72354), .B(n72357), .Y(n72359) );
  AND2X1 U44016 ( .A(n43763), .B(n44050), .Y(n42107) );
  AND2X1 U44017 ( .A(n43751), .B(n44009), .Y(n42108) );
  AND2X1 U44018 ( .A(n43730), .B(n44001), .Y(n42109) );
  AND2X1 U44019 ( .A(n43816), .B(n44019), .Y(n42110) );
  AND2X1 U44020 ( .A(n43741), .B(n44056), .Y(n42111) );
  AND2X1 U44021 ( .A(n38582), .B(n44027), .Y(n42112) );
  AND2X1 U44022 ( .A(n43763), .B(n44056), .Y(n42113) );
  AND2X1 U44023 ( .A(n43751), .B(n44019), .Y(n42114) );
  AND2X1 U44024 ( .A(n43729), .B(n44009), .Y(n42115) );
  AND2X1 U44025 ( .A(n43816), .B(n44027), .Y(n42116) );
  AND2X1 U44026 ( .A(n38582), .B(n44050), .Y(n42117) );
  AND2X1 U44027 ( .A(n43751), .B(n44027), .Y(n42118) );
  AND2X1 U44028 ( .A(n43816), .B(n44050), .Y(n42119) );
  AND2X1 U44029 ( .A(n38582), .B(n44056), .Y(n42120) );
  AND2X1 U44030 ( .A(n44815), .B(n31408), .Y(n31148) );
  OR2X1 U44031 ( .A(n42121), .B(n42122), .Y(n50040) );
  OR2X1 U44032 ( .A(n31460), .B(n31461), .Y(n42121) );
  OR2X1 U44033 ( .A(n32471), .B(n32472), .Y(n42122) );
  AND2X1 U44034 ( .A(n56623), .B(n56622), .Y(n42123) );
  AND2X1 U44035 ( .A(n43750), .B(n44050), .Y(n42124) );
  AND2X1 U44036 ( .A(n43729), .B(n44027), .Y(n42125) );
  AND2X1 U44037 ( .A(n43816), .B(n44057), .Y(n42126) );
  AND2X1 U44038 ( .A(n43504), .B(n44027), .Y(n42127) );
  AND2X1 U44039 ( .A(n43750), .B(n44057), .Y(n42128) );
  AND2X1 U44040 ( .A(n43729), .B(n44050), .Y(n42129) );
  AND2X1 U44041 ( .A(n43729), .B(n44057), .Y(n42130) );
  AND2X1 U44042 ( .A(n57247), .B(n73503), .Y(n42131) );
  OR2X1 U44043 ( .A(n25786), .B(n72835), .Y(n42132) );
  NAND2X1 U44044 ( .A(n26115), .B(n26116), .Y(n42133) );
  NAND2X1 U44045 ( .A(n26855), .B(n26856), .Y(n42134) );
  AND2X1 U44046 ( .A(n55061), .B(n73503), .Y(n42135) );
  AND2X1 U44047 ( .A(n57247), .B(n73173), .Y(n42136) );
  AND2X1 U44048 ( .A(n55061), .B(n73173), .Y(n42137) );
  AND2X1 U44049 ( .A(n58283), .B(n73173), .Y(n42138) );
  AND2X1 U44050 ( .A(n73173), .B(n73172), .Y(n42139) );
  AND2X1 U44051 ( .A(n72834), .B(n73173), .Y(n42140) );
  AND2X1 U44052 ( .A(n73167), .B(n73173), .Y(n42141) );
  AND2X1 U44053 ( .A(n58232), .B(n38383), .Y(n42142) );
  AND2X1 U44054 ( .A(n58229), .B(n73173), .Y(n42143) );
  AND2X1 U44055 ( .A(n58266), .B(n42962), .Y(n42144) );
  AND2X1 U44056 ( .A(n58478), .B(n73503), .Y(n42145) );
  OR2X1 U44057 ( .A(n59340), .B(n59341), .Y(n59342) );
  OR2X1 U44058 ( .A(n59122), .B(n59121), .Y(n59231) );
  OR2X1 U44059 ( .A(n59543), .B(n59544), .Y(n59545) );
  AND2X1 U44060 ( .A(n46019), .B(n45176), .Y(n42146) );
  XOR2X1 U44061 ( .A(n59891), .B(n60228), .Y(n59892) );
  AND2X1 U44062 ( .A(n42697), .B(n40512), .Y(n42147) );
  AND2X1 U44063 ( .A(n72811), .B(n42148), .Y(n59167) );
  AND2X1 U44064 ( .A(n40391), .B(n40228), .Y(n42148) );
  AND2X1 U44065 ( .A(n40398), .B(n45610), .Y(n42149) );
  NOR2X1 U44066 ( .A(n43726), .B(n40589), .Y(n42150) );
  XOR2X1 U44067 ( .A(n63221), .B(n62468), .Y(n42151) );
  XNOR2X1 U44068 ( .A(n42152), .B(n60966), .Y(n60967) );
  AND2X1 U44069 ( .A(n71546), .B(n62659), .Y(n42152) );
  AND2X1 U44070 ( .A(n61190), .B(n61189), .Y(n42153) );
  AND2X1 U44071 ( .A(n39669), .B(n48370), .Y(n42154) );
  NOR2X1 U44072 ( .A(n43727), .B(n43470), .Y(n42155) );
  XNOR2X1 U44073 ( .A(n42156), .B(n62937), .Y(n63241) );
  XOR2X1 U44074 ( .A(n63816), .B(n63231), .Y(n42156) );
  AND2X1 U44075 ( .A(n68620), .B(n42157), .Y(n68626) );
  OR2X1 U44076 ( .A(n44012), .B(n68623), .Y(n42157) );
  AND2X1 U44077 ( .A(n47674), .B(n43017), .Y(n42158) );
  AND2X1 U44078 ( .A(n39810), .B(n48372), .Y(n42159) );
  NOR2X1 U44079 ( .A(n43728), .B(n39944), .Y(n42160) );
  AND2X1 U44080 ( .A(n63568), .B(n63567), .Y(n42161) );
  NOR2X1 U44081 ( .A(n63552), .B(n39082), .Y(n42162) );
  XOR2X1 U44082 ( .A(n64079), .B(n42237), .Y(n64777) );
  XNOR2X1 U44083 ( .A(n64101), .B(n42163), .Y(n63818) );
  OR2X1 U44084 ( .A(n64102), .B(n63572), .Y(n42163) );
  AND2X1 U44085 ( .A(n47674), .B(n39669), .Y(n42164) );
  AND2X1 U44086 ( .A(n47674), .B(n48015), .Y(n42165) );
  AND2X1 U44087 ( .A(n38305), .B(n63817), .Y(n42166) );
  XOR2X1 U44088 ( .A(n65080), .B(n65772), .Y(n65379) );
  OR2X1 U44089 ( .A(n42167), .B(n42168), .Y(n50471) );
  AND2X1 U44090 ( .A(n50115), .B(n50117), .Y(n42167) );
  AND2X1 U44091 ( .A(n50010), .B(n50114), .Y(n42168) );
  OR2X1 U44092 ( .A(n42169), .B(n42170), .Y(n49999) );
  AND2X1 U44093 ( .A(n50411), .B(n49995), .Y(n42169) );
  AND2X1 U44094 ( .A(n49998), .B(n50410), .Y(n42170) );
  OR2X1 U44095 ( .A(n42171), .B(n42172), .Y(n49995) );
  AND2X1 U44096 ( .A(n50397), .B(n49991), .Y(n42171) );
  AND2X1 U44097 ( .A(n49994), .B(n50396), .Y(n42172) );
  OR2X1 U44098 ( .A(n42173), .B(n42174), .Y(n50199) );
  AND2X1 U44099 ( .A(n50469), .B(n50471), .Y(n42173) );
  AND2X1 U44100 ( .A(n50014), .B(n50468), .Y(n42174) );
  OR2X1 U44101 ( .A(n42175), .B(n42176), .Y(n50253) );
  AND2X1 U44102 ( .A(n50197), .B(n50199), .Y(n42175) );
  AND2X1 U44103 ( .A(n50019), .B(n50196), .Y(n42176) );
  OR2X1 U44104 ( .A(n42177), .B(n42178), .Y(n50117) );
  AND2X1 U44105 ( .A(n50213), .B(n50003), .Y(n42177) );
  AND2X1 U44106 ( .A(n50006), .B(n50212), .Y(n42178) );
  OR2X1 U44107 ( .A(n42179), .B(n42180), .Y(n50003) );
  AND2X1 U44108 ( .A(n50131), .B(n49999), .Y(n42179) );
  AND2X1 U44109 ( .A(n50002), .B(n50130), .Y(n42180) );
  AND2X1 U44110 ( .A(n40260), .B(n43862), .Y(n42181) );
  AND2X1 U44111 ( .A(n40260), .B(n43898), .Y(n42182) );
  XOR2X1 U44112 ( .A(n50213), .B(n50212), .Y(n50214) );
  XOR2X1 U44113 ( .A(n50131), .B(n50130), .Y(n50132) );
  XOR2X1 U44114 ( .A(n50411), .B(n50410), .Y(n50412) );
  XOR2X1 U44115 ( .A(n50397), .B(n50396), .Y(n50398) );
  AND2X1 U44116 ( .A(n40260), .B(n44025), .Y(n42183) );
  AND2X1 U44117 ( .A(n43613), .B(n42641), .Y(n42184) );
  XOR2X1 U44118 ( .A(n50268), .B(n50267), .Y(n50269) );
  AND2X1 U44119 ( .A(n43613), .B(n43724), .Y(n42185) );
  AND2X1 U44120 ( .A(n48226), .B(n48225), .Y(n42186) );
  AND2X1 U44121 ( .A(n43613), .B(n42661), .Y(n42187) );
  AND2X1 U44122 ( .A(n43613), .B(n42711), .Y(n42188) );
  AND2X1 U44123 ( .A(n58752), .B(n58751), .Y(n42189) );
  XOR2X1 U44124 ( .A(n50425), .B(n50424), .Y(n50426) );
  AND2X1 U44125 ( .A(n43613), .B(n43799), .Y(n42190) );
  AND2X1 U44126 ( .A(n43613), .B(n40474), .Y(n42191) );
  AND2X1 U44127 ( .A(n40627), .B(n43816), .Y(n42192) );
  AND2X1 U44128 ( .A(n58737), .B(n58736), .Y(n42193) );
  AND2X1 U44129 ( .A(n43740), .B(n44036), .Y(n42194) );
  AND2X1 U44130 ( .A(n43761), .B(n43851), .Y(n42195) );
  AND2X1 U44131 ( .A(n43822), .B(n43862), .Y(n42196) );
  AND2X1 U44132 ( .A(n58664), .B(n58663), .Y(n42197) );
  AND2X1 U44133 ( .A(n58653), .B(n58652), .Y(n42198) );
  AND2X1 U44134 ( .A(n58645), .B(n58644), .Y(n42199) );
  AND2X1 U44135 ( .A(n42859), .B(n45347), .Y(n42200) );
  AND2X1 U44136 ( .A(n58637), .B(n58636), .Y(n42201) );
  AND2X1 U44137 ( .A(n58616), .B(n58615), .Y(n42202) );
  AND2X1 U44138 ( .A(n58613), .B(n58612), .Y(n42203) );
  AND2X1 U44139 ( .A(n58602), .B(n58601), .Y(n42204) );
  AND2X1 U44140 ( .A(n42323), .B(n73503), .Y(n42205) );
  NAND2X1 U44141 ( .A(n27095), .B(n27096), .Y(n42206) );
  NAND2X1 U44142 ( .A(n27305), .B(n26242), .Y(n42207) );
  NOR2X1 U44143 ( .A(n42208), .B(n72833), .Y(n26162) );
  OR2X1 U44144 ( .A(n25792), .B(n72834), .Y(n42208) );
  AND2X1 U44145 ( .A(n42962), .B(n42327), .Y(n42209) );
  AND2X1 U44146 ( .A(n44078), .B(n44083), .Y(n42210) );
  AND2X1 U44147 ( .A(n58810), .B(n58809), .Y(n42211) );
  AND2X1 U44148 ( .A(n42327), .B(n73173), .Y(n42212) );
  NAND2X1 U44149 ( .A(n27201), .B(n27202), .Y(n42213) );
  AND2X1 U44150 ( .A(n42323), .B(n73173), .Y(n42214) );
  AND2X1 U44151 ( .A(n27326), .B(n73576), .Y(n42215) );
  OR2X1 U44152 ( .A(n24877), .B(n73575), .Y(n42216) );
  AND2X1 U44153 ( .A(n58279), .B(n58278), .Y(n42217) );
  AND2X1 U44154 ( .A(n16774), .B(n42218), .Y(n17160) );
  OR2X1 U44155 ( .A(n73464), .B(n43417), .Y(n42218) );
  AND2X1 U44156 ( .A(n44833), .B(n43375), .Y(n42219) );
  OR2X1 U44157 ( .A(n46894), .B(n46915), .Y(n59201) );
  XNOR2X1 U44158 ( .A(n39714), .B(n42220), .Y(n42817) );
  XNOR2X1 U44159 ( .A(n59153), .B(n59232), .Y(n42220) );
  AND2X1 U44160 ( .A(n59886), .B(n59887), .Y(n42221) );
  AND2X1 U44161 ( .A(n38848), .B(n36759), .Y(n42222) );
  AND2X1 U44162 ( .A(n38825), .B(n36707), .Y(n42223) );
  OR2X1 U44163 ( .A(n46389), .B(n46364), .Y(n70051) );
  AND2X1 U44164 ( .A(n40593), .B(n42486), .Y(n42224) );
  OR2X1 U44165 ( .A(n60960), .B(n60961), .Y(n71546) );
  AND2X1 U44166 ( .A(n61188), .B(n61187), .Y(n42225) );
  AND2X1 U44167 ( .A(n63835), .B(n63550), .Y(n42226) );
  AND2X1 U44168 ( .A(n45290), .B(n45289), .Y(n42227) );
  AND2X1 U44169 ( .A(n64083), .B(n48624), .Y(n42228) );
  XNOR2X1 U44170 ( .A(n63556), .B(n42229), .Y(n63221) );
  XOR2X1 U44171 ( .A(n62464), .B(n62463), .Y(n42229) );
  AND2X1 U44172 ( .A(n42360), .B(n45446), .Y(n42230) );
  NOR2X1 U44173 ( .A(n42232), .B(n42233), .Y(n42231) );
  OR2X1 U44174 ( .A(n45165), .B(n45164), .Y(n42232) );
  OR2X1 U44175 ( .A(n38663), .B(n37392), .Y(n42233) );
  AND2X1 U44176 ( .A(n61180), .B(n61179), .Y(n42234) );
  AND2X1 U44177 ( .A(n48762), .B(n48761), .Y(n42235) );
  AND2X1 U44178 ( .A(n62914), .B(n62913), .Y(n42236) );
  AND2X1 U44179 ( .A(n63839), .B(n39653), .Y(n42237) );
  AND2X1 U44180 ( .A(n48899), .B(n48898), .Y(n42238) );
  AND2X1 U44181 ( .A(n47552), .B(n47551), .Y(n42239) );
  XOR2X1 U44182 ( .A(n56617), .B(n56616), .Y(u_fetch_N79) );
  AND2X1 U44183 ( .A(n49306), .B(n49305), .Y(n42240) );
  AND2X1 U44184 ( .A(n49034), .B(n49033), .Y(n42241) );
  AND2X1 U44185 ( .A(n49168), .B(n49167), .Y(n42242) );
  NOR2X1 U44186 ( .A(n42244), .B(n42245), .Y(n42243) );
  OR2X1 U44187 ( .A(n49429), .B(n49428), .Y(n42244) );
  AND2X1 U44188 ( .A(n42802), .B(n49490), .Y(n42245) );
  XOR2X1 U44189 ( .A(n42409), .B(n55992), .Y(u_fetch_N74) );
  NOR2X1 U44190 ( .A(n42247), .B(n42248), .Y(n42246) );
  OR2X1 U44191 ( .A(n47360), .B(n47359), .Y(n42247) );
  AND2X1 U44192 ( .A(n42803), .B(n47421), .Y(n42248) );
  XOR2X1 U44193 ( .A(n55623), .B(n55670), .Y(u_fetch_N70) );
  NOR2X1 U44194 ( .A(n42250), .B(n42251), .Y(n42249) );
  OR2X1 U44195 ( .A(n47182), .B(n47181), .Y(n42250) );
  AND2X1 U44196 ( .A(n42804), .B(n47243), .Y(n42251) );
  XOR2X1 U44197 ( .A(n55416), .B(n55467), .Y(u_fetch_N66) );
  AND2X1 U44198 ( .A(n43380), .B(n56767), .Y(n42252) );
  NOR2X1 U44199 ( .A(n40687), .B(n57397), .Y(n42253) );
  XOR2X1 U44200 ( .A(n42406), .B(n55251), .Y(u_fetch_N62) );
  AND2X1 U44201 ( .A(n51999), .B(n54435), .Y(n42254) );
  XOR2X1 U44202 ( .A(n54958), .B(n55023), .Y(u_fetch_N58) );
  NOR2X1 U44203 ( .A(n42256), .B(n42257), .Y(n42255) );
  OR2X1 U44204 ( .A(n49725), .B(n49724), .Y(n42256) );
  AND2X1 U44205 ( .A(n42801), .B(n49786), .Y(n42257) );
  AND2X1 U44206 ( .A(n50500), .B(n38001), .Y(n42258) );
  NOR2X1 U44207 ( .A(n42260), .B(n42261), .Y(n42259) );
  OR2X1 U44208 ( .A(n46789), .B(n46788), .Y(n42260) );
  AND2X1 U44209 ( .A(n42803), .B(n46850), .Y(n42261) );
  XOR2X1 U44210 ( .A(n54710), .B(n54769), .Y(u_fetch_N54) );
  AND2X1 U44211 ( .A(n43318), .B(n50496), .Y(n42262) );
  AND2X1 U44212 ( .A(n54372), .B(n43406), .Y(n42263) );
  AND2X1 U44213 ( .A(n51973), .B(n72840), .Y(n51943) );
  OR2X1 U44214 ( .A(n42264), .B(n51967), .Y(n57240) );
  OR2X1 U44215 ( .A(n51936), .B(n51965), .Y(n42264) );
  NOR2X1 U44216 ( .A(n42266), .B(n42267), .Y(n42265) );
  OR2X1 U44217 ( .A(n46462), .B(n46461), .Y(n42266) );
  AND2X1 U44218 ( .A(n42805), .B(n46523), .Y(n42267) );
  OR2X1 U44219 ( .A(n51968), .B(n51967), .Y(n42268) );
  NOR2X1 U44220 ( .A(n42270), .B(n42271), .Y(n42269) );
  OR2X1 U44221 ( .A(n46589), .B(n46588), .Y(n42270) );
  AND2X1 U44222 ( .A(n42806), .B(n46651), .Y(n42271) );
  NOR2X1 U44223 ( .A(n42273), .B(n42274), .Y(n42272) );
  OR2X1 U44224 ( .A(n46247), .B(n46246), .Y(n42273) );
  AND2X1 U44225 ( .A(n42801), .B(n46308), .Y(n42274) );
  NOR2X1 U44226 ( .A(n42276), .B(n42277), .Y(n42275) );
  OR2X1 U44227 ( .A(n46096), .B(n46095), .Y(n42276) );
  AND2X1 U44228 ( .A(n42802), .B(n46157), .Y(n42277) );
  XOR2X1 U44229 ( .A(n44637), .B(n43888), .Y(n50328) );
  NOR2X1 U44230 ( .A(n42279), .B(n42280), .Y(n42278) );
  OR2X1 U44231 ( .A(n45942), .B(n45941), .Y(n42279) );
  AND2X1 U44232 ( .A(n42803), .B(n46004), .Y(n42280) );
  XOR2X1 U44233 ( .A(n44637), .B(n73224), .Y(n49966) );
  NOR2X1 U44234 ( .A(n42282), .B(n42283), .Y(n42281) );
  OR2X1 U44235 ( .A(n45795), .B(n45794), .Y(n42282) );
  AND2X1 U44236 ( .A(n42804), .B(n45856), .Y(n42283) );
  NOR2X1 U44237 ( .A(n42285), .B(n42286), .Y(n42284) );
  OR2X1 U44238 ( .A(n45384), .B(n45383), .Y(n42285) );
  AND2X1 U44239 ( .A(n42806), .B(n45445), .Y(n42286) );
  OR2X1 U44240 ( .A(n42287), .B(n42288), .Y(n73379) );
  OR2X1 U44241 ( .A(n45309), .B(n45308), .Y(n42287) );
  AND2X1 U44242 ( .A(n42801), .B(n45380), .Y(n42288) );
  XOR2X1 U44243 ( .A(n44637), .B(n43917), .Y(n50449) );
  NOR2X1 U44244 ( .A(n42290), .B(n42291), .Y(n42289) );
  OR2X1 U44245 ( .A(n45546), .B(n45545), .Y(n42290) );
  AND2X1 U44246 ( .A(n42802), .B(n45607), .Y(n42291) );
  AND2X1 U44247 ( .A(n43013), .B(n44635), .Y(n42292) );
  XOR2X1 U44248 ( .A(n50078), .B(n50079), .Y(n50081) );
  XOR2X1 U44249 ( .A(n44638), .B(n44002), .Y(n50213) );
  XNOR2X1 U44250 ( .A(n58760), .B(n42293), .Y(n57318) );
  OR2X1 U44251 ( .A(n57088), .B(n57087), .Y(n42293) );
  OR2X1 U44252 ( .A(n42294), .B(n42295), .Y(n50045) );
  NAND2X1 U44253 ( .A(n45002), .B(n45001), .Y(n42294) );
  OR2X1 U44254 ( .A(n45154), .B(n45153), .Y(n42295) );
  NOR2X1 U44255 ( .A(n50615), .B(n39625), .Y(n42296) );
  XNOR2X1 U44256 ( .A(n42297), .B(n44023), .Y(n50197) );
  INVX1 U44257 ( .A(n44638), .Y(n42297) );
  AND2X1 U44258 ( .A(n42922), .B(n49902), .Y(n42298) );
  AND2X1 U44259 ( .A(n58629), .B(n58628), .Y(n42299) );
  AND2X1 U44260 ( .A(n58591), .B(n58590), .Y(n42300) );
  AND2X1 U44261 ( .A(n58583), .B(n58582), .Y(n42301) );
  INVX1 U44262 ( .A(n72829), .Y(n42302) );
  AND2X1 U44263 ( .A(n58575), .B(n58574), .Y(n42303) );
  AND2X1 U44264 ( .A(n73539), .B(n73173), .Y(n42304) );
  AND2X1 U44265 ( .A(n58800), .B(n58799), .Y(n42305) );
  AND2X1 U44266 ( .A(n58453), .B(n38824), .Y(n42306) );
  AND2X1 U44267 ( .A(n58279), .B(n58276), .Y(n42307) );
  AND2X1 U44268 ( .A(n72840), .B(n73517), .Y(n42308) );
  AND2X1 U44269 ( .A(n16562), .B(n42309), .Y(n17328) );
  AND2X1 U44270 ( .A(n17331), .B(n16815), .Y(n42309) );
  AND2X1 U44271 ( .A(n51411), .B(n73525), .Y(n42310) );
  AND2X1 U44272 ( .A(n42948), .B(n15846), .Y(n42311) );
  AND2X1 U44273 ( .A(n42949), .B(n16449), .Y(n42312) );
  AND2X1 U44274 ( .A(n42948), .B(n15801), .Y(n42313) );
  AND2X1 U44275 ( .A(n42949), .B(n16048), .Y(n42314) );
  AND2X1 U44276 ( .A(n51411), .B(n15742), .Y(n42315) );
  AND2X1 U44277 ( .A(n57331), .B(n73523), .Y(n42316) );
  AND2X1 U44278 ( .A(n42947), .B(n16181), .Y(n42317) );
  AND2X1 U44279 ( .A(n57359), .B(n73430), .Y(n42318) );
  AND2X1 U44280 ( .A(n43415), .B(n15805), .Y(n42319) );
  AND2X1 U44281 ( .A(n43415), .B(n16181), .Y(n42320) );
  AND2X1 U44282 ( .A(n43415), .B(n15846), .Y(n42321) );
  AND2X1 U44283 ( .A(n43415), .B(n16042), .Y(n42322) );
  AND2X1 U44284 ( .A(n58254), .B(n58233), .Y(n42323) );
  AND2X1 U44285 ( .A(n42451), .B(n15977), .Y(n42324) );
  OR2X1 U44286 ( .A(n73374), .B(n42325), .Y(n58521) );
  AND2X1 U44287 ( .A(n24365), .B(n42439), .Y(n42325) );
  AND2X1 U44288 ( .A(n43419), .B(n15977), .Y(n42326) );
  AND2X1 U44289 ( .A(n73506), .B(n38501), .Y(n42327) );
  OR2X1 U44290 ( .A(n42329), .B(n42328), .Y(n45619) );
  INVX1 U44291 ( .A(n45534), .Y(n42328) );
  OR2X1 U44292 ( .A(n40579), .B(n38637), .Y(n42329) );
  NOR2X1 U44293 ( .A(n42330), .B(n42331), .Y(n42838) );
  OR2X1 U44294 ( .A(n46530), .B(n46529), .Y(n42330) );
  AND2X1 U44295 ( .A(n40490), .B(n46568), .Y(n42331) );
  OR2X1 U44296 ( .A(n42332), .B(n42333), .Y(n72741) );
  OR2X1 U44297 ( .A(n47346), .B(n47345), .Y(n42332) );
  OR2X1 U44298 ( .A(n47358), .B(n47357), .Y(n42333) );
  OR2X1 U44299 ( .A(n49624), .B(n37148), .Y(n42334) );
  OR2X1 U44300 ( .A(n46749), .B(n46748), .Y(n42335) );
  AND2X1 U44301 ( .A(n40490), .B(n46785), .Y(n42336) );
  OR2X1 U44302 ( .A(n42337), .B(n42338), .Y(n72807) );
  OR2X1 U44303 ( .A(n47302), .B(n47301), .Y(n42338) );
  NOR2X1 U44304 ( .A(n42340), .B(n42341), .Y(n42339) );
  OR2X1 U44305 ( .A(n49654), .B(n49653), .Y(n42340) );
  OR2X1 U44306 ( .A(n49704), .B(n49703), .Y(n42341) );
  OR2X1 U44307 ( .A(n42342), .B(n42343), .Y(n72766) );
  OR2X1 U44308 ( .A(n49413), .B(n49412), .Y(n42342) );
  OR2X1 U44309 ( .A(n49427), .B(n49426), .Y(n42343) );
  NOR2X1 U44310 ( .A(n42345), .B(n42346), .Y(n42344) );
  OR2X1 U44311 ( .A(n49714), .B(n49713), .Y(n42345) );
  OR2X1 U44312 ( .A(n49723), .B(n49722), .Y(n42346) );
  AND2X1 U44313 ( .A(n46243), .B(n46242), .Y(n42347) );
  OR2X1 U44314 ( .A(n47177), .B(n47176), .Y(n42349) );
  NOR2X1 U44315 ( .A(n42351), .B(n42352), .Y(n42350) );
  OR2X1 U44316 ( .A(n46582), .B(n46581), .Y(n42351) );
  OR2X1 U44317 ( .A(n46973), .B(n46972), .Y(n42353) );
  OR2X1 U44318 ( .A(n46985), .B(n46984), .Y(n42354) );
  OR2X1 U44319 ( .A(n42355), .B(n42356), .Y(n72787) );
  OR2X1 U44320 ( .A(n49357), .B(n49356), .Y(n42355) );
  OR2X1 U44321 ( .A(n49369), .B(n49368), .Y(n42356) );
  NAND2X1 U44322 ( .A(n42357), .B(n42358), .Y(n46782) );
  NOR2X1 U44323 ( .A(n46769), .B(n46768), .Y(n42357) );
  NOR2X1 U44324 ( .A(n46771), .B(n46770), .Y(n42358) );
  OR2X1 U44325 ( .A(n49699), .B(n42359), .Y(n46067) );
  AND2X1 U44326 ( .A(n46044), .B(n46043), .Y(n42359) );
  AND2X1 U44327 ( .A(n45276), .B(n45533), .Y(n42360) );
  AND2X1 U44328 ( .A(n45173), .B(n42361), .Y(n45520) );
  AND2X1 U44329 ( .A(n45175), .B(n45174), .Y(n42361) );
  NOR2X1 U44330 ( .A(n42364), .B(n42363), .Y(n42362) );
  INVX1 U44331 ( .A(n42724), .Y(n42363) );
  OR2X1 U44332 ( .A(n42686), .B(n42728), .Y(n42364) );
  OR2X1 U44333 ( .A(n42365), .B(n53762), .Y(n46585) );
  OR2X1 U44334 ( .A(n46583), .B(n40152), .Y(n42365) );
  OR2X1 U44335 ( .A(n45537), .B(n45536), .Y(n42366) );
  NOR2X1 U44336 ( .A(n42368), .B(n42369), .Y(n42367) );
  OR2X1 U44337 ( .A(n45695), .B(n45694), .Y(n42368) );
  OR2X1 U44338 ( .A(n45701), .B(n45700), .Y(n42369) );
  OR2X1 U44339 ( .A(n42365), .B(n55947), .Y(n45930) );
  AND2X1 U44340 ( .A(n44983), .B(n42685), .Y(n42370) );
  OR2X1 U44341 ( .A(n42371), .B(n42372), .Y(n72780) );
  OR2X1 U44342 ( .A(n47473), .B(n47472), .Y(n42371) );
  OR2X1 U44343 ( .A(n47487), .B(n47486), .Y(n42372) );
  AND2X1 U44344 ( .A(n45534), .B(n45533), .Y(n42373) );
  OR2X1 U44345 ( .A(n59148), .B(n59149), .Y(n59150) );
  OR2X1 U44346 ( .A(n42365), .B(n53889), .Y(n46401) );
  OR2X1 U44347 ( .A(n42374), .B(n56124), .Y(n45785) );
  OR2X1 U44348 ( .A(n46583), .B(n38441), .Y(n42374) );
  AND2X1 U44349 ( .A(n44994), .B(n42687), .Y(n42375) );
  AND2X1 U44350 ( .A(n62902), .B(n47930), .Y(n42376) );
  AND2X1 U44351 ( .A(n45313), .B(n45312), .Y(n42377) );
  AND2X1 U44352 ( .A(n48174), .B(n42685), .Y(n42378) );
  AND2X1 U44353 ( .A(n48398), .B(n48397), .Y(n42379) );
  OR2X1 U44354 ( .A(n42380), .B(n48186), .Y(n48172) );
  OR2X1 U44355 ( .A(n36810), .B(n48109), .Y(n42380) );
  OR2X1 U44356 ( .A(n42381), .B(n42382), .Y(n72806) );
  OR2X1 U44357 ( .A(n48813), .B(n48812), .Y(n42381) );
  OR2X1 U44358 ( .A(n48825), .B(n48824), .Y(n42382) );
  NOR2X1 U44359 ( .A(n42384), .B(n42385), .Y(n42383) );
  AND2X1 U44360 ( .A(n45256), .B(n45615), .Y(n42384) );
  AND2X1 U44361 ( .A(n45261), .B(n45260), .Y(n42385) );
  OR2X1 U44362 ( .A(n42386), .B(n42387), .Y(n72810) );
  OR2X1 U44363 ( .A(n48675), .B(n48674), .Y(n42386) );
  OR2X1 U44364 ( .A(n48688), .B(n48687), .Y(n42387) );
  OR2X1 U44365 ( .A(n42388), .B(n42389), .Y(n72765) );
  OR2X1 U44366 ( .A(n48515), .B(n48514), .Y(n42388) );
  OR2X1 U44367 ( .A(n48528), .B(n48527), .Y(n42389) );
  OR2X1 U44368 ( .A(n42390), .B(n42391), .Y(n72786) );
  OR2X1 U44369 ( .A(n48451), .B(n48450), .Y(n42390) );
  OR2X1 U44370 ( .A(n48464), .B(n48463), .Y(n42391) );
  AND2X1 U44371 ( .A(n61176), .B(n62907), .Y(n42392) );
  OR2X1 U44372 ( .A(n42393), .B(n42394), .Y(n72819) );
  OR2X1 U44373 ( .A(n47603), .B(n47602), .Y(n42393) );
  OR2X1 U44374 ( .A(n47617), .B(n47616), .Y(n42394) );
  OR2X1 U44375 ( .A(n42395), .B(n42396), .Y(n72759) );
  OR2X1 U44376 ( .A(n48088), .B(n48087), .Y(n42395) );
  OR2X1 U44377 ( .A(n48102), .B(n48101), .Y(n42396) );
  NOR2X1 U44378 ( .A(n42398), .B(n55416), .Y(n42397) );
  NOR2X1 U44379 ( .A(n42400), .B(n54958), .Y(n42399) );
  AND2X1 U44380 ( .A(mem_i_pc_o[2]), .B(mem_i_pc_o[3]), .Y(n42401) );
  AND2X1 U44381 ( .A(n42405), .B(n22), .Y(n42402) );
  NOR2X1 U44382 ( .A(n42404), .B(n55623), .Y(n42403) );
  NOR2X1 U44383 ( .A(n42407), .B(n42406), .Y(n42405) );
  INVX1 U44384 ( .A(n9), .Y(n42406) );
  NOR2X1 U44385 ( .A(n42410), .B(n42409), .Y(n42408) );
  INVX1 U44386 ( .A(n23), .Y(n42409) );
  AND2X1 U44387 ( .A(n42408), .B(n19), .Y(n42411) );
  AND2X1 U44388 ( .A(n42397), .B(n20), .Y(n42412) );
  AND2X1 U44389 ( .A(n42411), .B(n18), .Y(n42414) );
  AND2X1 U44390 ( .A(n42399), .B(mem_i_pc_o[11]), .Y(n42415) );
  AND2X1 U44391 ( .A(n42417), .B(mem_i_pc_o[7]), .Y(n42416) );
  AND2X1 U44392 ( .A(n54771), .B(mem_i_pc_o[5]), .Y(n42417) );
  OR2X1 U44393 ( .A(n42418), .B(n42419), .Y(n72779) );
  OR2X1 U44394 ( .A(n47912), .B(n47911), .Y(n42418) );
  OR2X1 U44395 ( .A(n47926), .B(n47925), .Y(n42419) );
  XOR2X1 U44396 ( .A(n19), .B(n42408), .Y(u_fetch_N76) );
  XOR2X1 U44397 ( .A(n11), .B(n42413), .Y(u_fetch_N73) );
  XOR2X1 U44398 ( .A(n22), .B(n42405), .Y(u_fetch_N64) );
  AND2X1 U44399 ( .A(n56710), .B(n56709), .Y(n42420) );
  AND2X1 U44400 ( .A(n56555), .B(n56554), .Y(n42421) );
  AND2X1 U44401 ( .A(n56369), .B(n56368), .Y(n42422) );
  AND2X1 U44402 ( .A(n56629), .B(n56628), .Y(n42423) );
  OR2X1 U44403 ( .A(n55306), .B(n29013), .Y(n51998) );
  XOR2X1 U44404 ( .A(n21), .B(n42415), .Y(u_fetch_N61) );
  XOR2X1 U44405 ( .A(mem_i_pc_o[11]), .B(n42399), .Y(u_fetch_N60) );
  XOR2X1 U44406 ( .A(mem_i_pc_o[8]), .B(n42416), .Y(u_fetch_N57) );
  XOR2X1 U44407 ( .A(mem_i_pc_o[7]), .B(n42417), .Y(u_fetch_N56) );
  AND2X1 U44408 ( .A(n57593), .B(n57579), .Y(n42424) );
  AND2X1 U44409 ( .A(n57593), .B(n50633), .Y(n42425) );
  AND2X1 U44410 ( .A(n54375), .B(n54374), .Y(n42426) );
  AND2X1 U44411 ( .A(n54359), .B(n57559), .Y(n42427) );
  XOR2X1 U44412 ( .A(mem_i_pc_o[4]), .B(n42401), .Y(u_fetch_N53) );
  XOR2X1 U44413 ( .A(mem_i_pc_o[2]), .B(mem_i_pc_o[3]), .Y(u_fetch_N52) );
  AND2X1 U44414 ( .A(n24429), .B(n42428), .Y(u_decode_N757) );
  AND2X1 U44415 ( .A(n50655), .B(n57593), .Y(n42428) );
  OR2X1 U44416 ( .A(n54381), .B(n42429), .Y(n54446) );
  AND2X1 U44417 ( .A(n54384), .B(n54383), .Y(n42429) );
  AND2X1 U44418 ( .A(n42430), .B(opcode_instr_w_25), .Y(n49889) );
  OR2X1 U44419 ( .A(n49888), .B(n49887), .Y(n42430) );
  AND2X1 U44420 ( .A(n42431), .B(n42432), .Y(n45703) );
  AND2X1 U44421 ( .A(n49896), .B(n57677), .Y(n42431) );
  AND2X1 U44422 ( .A(n58159), .B(n50028), .Y(n42432) );
  NOR2X1 U44423 ( .A(n50693), .B(n50692), .Y(n42433) );
  AND2X1 U44424 ( .A(n50658), .B(n58541), .Y(n42434) );
  AND2X1 U44425 ( .A(n57316), .B(n16593), .Y(n42435) );
  XOR2X1 U44426 ( .A(n54899), .B(n54898), .Y(n54900) );
  XOR2X1 U44427 ( .A(n54781), .B(n54780), .Y(n54782) );
  XOR2X1 U44428 ( .A(n54823), .B(n54822), .Y(n54824) );
  XOR2X1 U44429 ( .A(n54721), .B(n54720), .Y(n54722) );
  XOR2X1 U44430 ( .A(n54658), .B(n54657), .Y(n54659) );
  OR2X1 U44431 ( .A(n57473), .B(n42436), .Y(n45147) );
  AND2X1 U44432 ( .A(n42629), .B(n45350), .Y(n42436) );
  AND2X1 U44433 ( .A(n30493), .B(n50257), .Y(n42437) );
  AND2X1 U44434 ( .A(n57628), .B(n42438), .Y(n35945) );
  INVX1 U44435 ( .A(n37436), .Y(n42438) );
  AND2X1 U44436 ( .A(n57351), .B(n28934), .Y(n42439) );
  XNOR2X1 U44437 ( .A(n54395), .B(n42440), .Y(n54396) );
  XNOR2X1 U44438 ( .A(n54394), .B(n54393), .Y(n42440) );
  AND2X1 U44439 ( .A(n58278), .B(n45159), .Y(n42441) );
  AND2X1 U44440 ( .A(n42962), .B(n27964), .Y(n42442) );
  NAND2X1 U44441 ( .A(n27560), .B(n27960), .Y(n42443) );
  OR2X1 U44442 ( .A(n24877), .B(n27964), .Y(n42444) );
  AND2X1 U44443 ( .A(n73367), .B(n58256), .Y(n42445) );
  AND2X1 U44444 ( .A(n42588), .B(n39766), .Y(n42446) );
  AND2X1 U44445 ( .A(n28510), .B(n51990), .Y(n42447) );
  AND2X1 U44446 ( .A(n42947), .B(n15845), .Y(n42448) );
  AND2X1 U44447 ( .A(n42947), .B(n15414), .Y(n42449) );
  AND2X1 U44448 ( .A(n42947), .B(n15441), .Y(n42450) );
  AND2X1 U44449 ( .A(n57331), .B(n16593), .Y(n42451) );
  AND2X1 U44450 ( .A(n42949), .B(n16290), .Y(n42452) );
  AND2X1 U44451 ( .A(n58822), .B(n73428), .Y(n42453) );
  AND2X1 U44452 ( .A(n58599), .B(n58598), .Y(n42454) );
  AND2X1 U44453 ( .A(n50866), .B(n58544), .Y(n42455) );
  AND2X1 U44454 ( .A(n43415), .B(n15728), .Y(n42456) );
  AND2X1 U44455 ( .A(n43424), .B(n15845), .Y(n42457) );
  AND2X1 U44456 ( .A(n43424), .B(n15443), .Y(n42458) );
  AND2X1 U44457 ( .A(n42451), .B(n15845), .Y(n42459) );
  AND2X1 U44458 ( .A(n57430), .B(n58521), .Y(n42460) );
  AND2X1 U44459 ( .A(n42559), .B(n58223), .Y(n42461) );
  AND2X1 U44460 ( .A(n55202), .B(n58312), .Y(n42462) );
  AND2X1 U44461 ( .A(n55146), .B(n58305), .Y(n42463) );
  AND2X1 U44462 ( .A(n58167), .B(n58216), .Y(n42464) );
  AND2X1 U44463 ( .A(n55038), .B(n58291), .Y(n42465) );
  OR2X1 U44464 ( .A(n46903), .B(n42466), .Y(n46410) );
  NOR2X1 U44465 ( .A(n42469), .B(n42763), .Y(n42467) );
  INVX1 U44466 ( .A(n40453), .Y(n42468) );
  OR2X1 U44467 ( .A(opcode_opcode_w[20]), .B(opcode_opcode_w[22]), .Y(n42469)
         );
  OR2X1 U44468 ( .A(opcode_opcode_w[22]), .B(n42470), .Y(n45168) );
  OR2X1 U44469 ( .A(n42763), .B(n42739), .Y(n42470) );
  OR2X1 U44470 ( .A(n42471), .B(n49610), .Y(n47270) );
  OR2X1 U44471 ( .A(n49400), .B(n36856), .Y(n42472) );
  OR2X1 U44472 ( .A(n40497), .B(n36861), .Y(n42473) );
  OR2X1 U44473 ( .A(n42474), .B(n49710), .Y(n49711) );
  NAND2X1 U44474 ( .A(n2497), .B(n40514), .Y(n42475) );
  OR2X1 U44475 ( .A(n42476), .B(n46312), .Y(n46313) );
  OR2X1 U44476 ( .A(n42477), .B(n46382), .Y(n46384) );
  AND2X1 U44477 ( .A(n42478), .B(n42479), .Y(n49626) );
  OR2X1 U44478 ( .A(n49624), .B(n37135), .Y(n42478) );
  OR2X1 U44479 ( .A(n42908), .B(n37132), .Y(n42479) );
  OR2X1 U44480 ( .A(n42480), .B(n42891), .Y(n46028) );
  NOR2X1 U44481 ( .A(n42702), .B(n46326), .Y(n42481) );
  OR2X1 U44482 ( .A(n42482), .B(n46231), .Y(n46020) );
  OR2X1 U44483 ( .A(n42483), .B(n46007), .Y(n46008) );
  AND2X1 U44484 ( .A(n42484), .B(n42485), .Y(n49627) );
  OR2X1 U44485 ( .A(n40517), .B(n37134), .Y(n42484) );
  OR2X1 U44486 ( .A(n40277), .B(n37131), .Y(n42485) );
  AND2X1 U44487 ( .A(opcode_opcode_w[24]), .B(n42761), .Y(n42486) );
  AND2X1 U44488 ( .A(n44959), .B(n38115), .Y(n42487) );
  OR2X1 U44489 ( .A(n42739), .B(n42489), .Y(n58469) );
  OR2X1 U44490 ( .A(n40453), .B(opcode_opcode_w[22]), .Y(n42489) );
  AND2X1 U44491 ( .A(n42779), .B(n2561), .Y(n46762) );
  NOR2X1 U44492 ( .A(n40604), .B(n42740), .Y(n42490) );
  OR2X1 U44493 ( .A(n42491), .B(n40497), .Y(n46169) );
  AND2X1 U44494 ( .A(n42492), .B(n42493), .Y(n45313) );
  XNOR2X1 U44495 ( .A(writeback_exec_idx_w[0]), .B(n42729), .Y(n42492) );
  XNOR2X1 U44496 ( .A(writeback_exec_idx_w[3]), .B(n42669), .Y(n42493) );
  AND2X1 U44497 ( .A(n38739), .B(n42494), .Y(n48012) );
  AND2X1 U44498 ( .A(n48008), .B(n1971), .Y(n42494) );
  NOR2X1 U44499 ( .A(n42496), .B(n42497), .Y(n42495) );
  OR2X1 U44500 ( .A(n48607), .B(n42854), .Y(n42497) );
  AND2X1 U44501 ( .A(writeback_exec_idx_w[4]), .B(n42747), .Y(n42498) );
  AND2X1 U44502 ( .A(n42499), .B(n42500), .Y(n47350) );
  OR2X1 U44503 ( .A(n40407), .B(n37178), .Y(n42499) );
  OR2X1 U44504 ( .A(n43142), .B(n42899), .Y(n42500) );
  OR2X1 U44505 ( .A(n42501), .B(n57609), .Y(n48339) );
  AND2X1 U44506 ( .A(n42502), .B(n42503), .Y(n45312) );
  XNOR2X1 U44507 ( .A(writeback_exec_idx_w[1]), .B(n42724), .Y(n42502) );
  XNOR2X1 U44508 ( .A(writeback_exec_idx_w[2]), .B(n42685), .Y(n42503) );
  AND2X1 U44509 ( .A(n44970), .B(opcode_opcode_w[17]), .Y(n42504) );
  OR2X1 U44510 ( .A(n42505), .B(n46007), .Y(n45620) );
  OR2X1 U44511 ( .A(n42506), .B(n39654), .Y(n46162) );
  OR2X1 U44512 ( .A(n42507), .B(n46236), .Y(n45608) );
  OR2X1 U44513 ( .A(n42508), .B(n49604), .Y(n46159) );
  OR2X1 U44514 ( .A(n42509), .B(n48116), .Y(n48027) );
  OR2X1 U44515 ( .A(n42510), .B(n46207), .Y(n45616) );
  OR2X1 U44516 ( .A(n42511), .B(n57608), .Y(n45611) );
  OR2X1 U44517 ( .A(n42512), .B(n38712), .Y(n49057) );
  OR2X1 U44518 ( .A(n42513), .B(n38711), .Y(n47445) );
  OR2X1 U44519 ( .A(n42514), .B(n38712), .Y(n48922) );
  AND2X1 U44520 ( .A(n2921), .B(n39449), .Y(n45209) );
  AND2X1 U44521 ( .A(n2918), .B(n36759), .Y(n45210) );
  AND2X1 U44522 ( .A(n45534), .B(n42517), .Y(n45261) );
  AND2X1 U44523 ( .A(writeback_exec_value_w[31]), .B(n45533), .Y(n42517) );
  OR2X1 U44524 ( .A(n42518), .B(n51965), .Y(n50042) );
  INVX1 U44525 ( .A(n42439), .Y(n42518) );
  AND2X1 U44526 ( .A(n42519), .B(n42520), .Y(n50033) );
  OR2X1 U44527 ( .A(opcode_instr_w_25), .B(n49895), .Y(n42519) );
  OR2X1 U44528 ( .A(n58158), .B(n50032), .Y(n42520) );
  AND2X1 U44529 ( .A(u_fetch_branch_valid_q), .B(n38001), .Y(n42521) );
  OR2X1 U44530 ( .A(n42522), .B(n42523), .Y(n21) );
  OR2X1 U44531 ( .A(n50324), .B(n55088), .Y(n42522) );
  NOR2X1 U44532 ( .A(n1770), .B(n43314), .Y(n42523) );
  NAND2X1 U44533 ( .A(n42524), .B(n58126), .Y(n50493) );
  INVX1 U44534 ( .A(mem_i_accept_i), .Y(n42524) );
  MX2X1 U44535 ( .A(challenge[7]), .B(n43380), .S0(n44860), .Y(n17215) );
  OR2X1 U44536 ( .A(n57960), .B(n42525), .Y(n8559) );
  AND2X1 U44537 ( .A(n57398), .B(n58183), .Y(n42525) );
  OR2X1 U44538 ( .A(n42526), .B(n43353), .Y(n49734) );
  OR2X1 U44539 ( .A(n42527), .B(n47637), .Y(n49775) );
  OR2X1 U44540 ( .A(n42528), .B(n57609), .Y(n49825) );
  OR2X1 U44541 ( .A(n42529), .B(n45350), .Y(n49843) );
  OR2X1 U44542 ( .A(n42530), .B(n45347), .Y(n49839) );
  OR2X1 U44543 ( .A(n42531), .B(n43046), .Y(n49840) );
  OR2X1 U44544 ( .A(n42532), .B(n45317), .Y(n49811) );
  AND2X1 U44545 ( .A(n42533), .B(n42534), .Y(n49890) );
  OR2X1 U44546 ( .A(n58158), .B(n45703), .Y(n42533) );
  AND2X1 U44547 ( .A(opcode_instr_w_28), .B(n45705), .Y(n42534) );
  AND2X1 U44548 ( .A(n56831), .B(n36599), .Y(n56825) );
  OR2X1 U44549 ( .A(n42535), .B(n42536), .Y(n58216) );
  OR2X1 U44550 ( .A(n44953), .B(n58189), .Y(n42535) );
  NOR2X1 U44551 ( .A(n35956), .B(n37433), .Y(n42536) );
  OR2X1 U44552 ( .A(n73367), .B(n58560), .Y(n17534) );
  OR2X1 U44553 ( .A(n42537), .B(n42538), .Y(n44907) );
  XNOR2X1 U44554 ( .A(n2817), .B(u_mmu_dtlb_va_addr_q[25]), .Y(n42537) );
  XNOR2X1 U44555 ( .A(n2785), .B(u_mmu_dtlb_va_addr_q[27]), .Y(n42538) );
  OR2X1 U44556 ( .A(n42539), .B(n42540), .Y(n44889) );
  XNOR2X1 U44557 ( .A(n8296), .B(u_mmu_dtlb_va_addr_q[12]), .Y(n42539) );
  XNOR2X1 U44558 ( .A(n8328), .B(u_mmu_dtlb_va_addr_q[27]), .Y(n42540) );
  OR2X1 U44559 ( .A(n42541), .B(n42542), .Y(n44923) );
  XNOR2X1 U44560 ( .A(n1869), .B(u_mmu_dtlb_va_addr_q[15]), .Y(n42541) );
  XNOR2X1 U44561 ( .A(n2882), .B(u_mmu_dtlb_va_addr_q[17]), .Y(n42542) );
  OR2X1 U44562 ( .A(n42543), .B(n42544), .Y(n58179) );
  AND2X1 U44563 ( .A(u_csr_N3161), .B(u_csr_N3162), .Y(n42544) );
  OR2X1 U44564 ( .A(n58338), .B(n42545), .Y(n30711) );
  NOR2X1 U44565 ( .A(n44838), .B(n57890), .Y(n42545) );
  OR2X1 U44566 ( .A(n42546), .B(n59119), .Y(n72732) );
  OR2X1 U44567 ( .A(n42547), .B(n42548), .Y(n29470) );
  NOR2X1 U44568 ( .A(n29472), .B(n37445), .Y(n42548) );
  OR2X1 U44569 ( .A(n42549), .B(n42550), .Y(n29454) );
  NOR2X1 U44570 ( .A(n29456), .B(n37461), .Y(n42550) );
  OR2X1 U44571 ( .A(n42551), .B(n42552), .Y(n29438) );
  NOR2X1 U44572 ( .A(n29440), .B(n1471), .Y(n42552) );
  OR2X1 U44573 ( .A(n42553), .B(n42554), .Y(n29422) );
  NOR2X1 U44574 ( .A(n29424), .B(n1511), .Y(n42554) );
  OR2X1 U44575 ( .A(n42555), .B(n42556), .Y(n29486) );
  NOR2X1 U44576 ( .A(n29488), .B(n37437), .Y(n42556) );
  NOR2X1 U44577 ( .A(n42557), .B(n42558), .Y(n45160) );
  NAND2X1 U44578 ( .A(n8647), .B(n8954), .Y(n42557) );
  AND2X1 U44579 ( .A(n1887), .B(n8810), .Y(n42559) );
  AND2X1 U44580 ( .A(n45704), .B(n36761), .Y(n49898) );
  XOR2X1 U44581 ( .A(n50442), .B(n42560), .Y(n50353) );
  XNOR2X1 U44582 ( .A(opcode_pc_w[18]), .B(n44836), .Y(n42560) );
  XOR2X1 U44583 ( .A(n50288), .B(n42561), .Y(n50289) );
  XNOR2X1 U44584 ( .A(opcode_pc_w[14]), .B(n44836), .Y(n42561) );
  XOR2X1 U44585 ( .A(n50325), .B(n42562), .Y(n50326) );
  XNOR2X1 U44586 ( .A(opcode_pc_w[15]), .B(n44836), .Y(n42562) );
  MX2X1 U44587 ( .A(n59092), .B(n59093), .S0(n38313), .Y(n14243) );
  XOR2X1 U44588 ( .A(n50148), .B(n42563), .Y(n50149) );
  XNOR2X1 U44589 ( .A(opcode_pc_w[16]), .B(n42851), .Y(n42563) );
  AND2X1 U44590 ( .A(u_csr_csr_mepc_q[13]), .B(n42131), .Y(n42564) );
  AND2X1 U44591 ( .A(u_csr_csr_mepc_q[20]), .B(n42131), .Y(n42565) );
  AND2X1 U44592 ( .A(u_csr_csr_mepc_q[18]), .B(n42131), .Y(n42566) );
  XOR2X1 U44593 ( .A(n50076), .B(n50349), .Y(n50077) );
  OR2X1 U44594 ( .A(n54609), .B(n58426), .Y(n54668) );
  OR2X1 U44595 ( .A(n54668), .B(n58431), .Y(n54669) );
  AND2X1 U44596 ( .A(n54832), .B(opcode_pc_w[8]), .Y(n42567) );
  AND2X1 U44597 ( .A(n54908), .B(opcode_pc_w[10]), .Y(n42568) );
  AND2X1 U44598 ( .A(u_csr_csr_sepc_q[13]), .B(n73501), .Y(n42569) );
  AND2X1 U44599 ( .A(u_csr_csr_sepc_q[21]), .B(n73501), .Y(n42570) );
  AND2X1 U44600 ( .A(u_csr_csr_sepc_q[19]), .B(n73501), .Y(n42571) );
  AND2X1 U44601 ( .A(u_csr_csr_sepc_q[17]), .B(n73501), .Y(n42572) );
  AND2X1 U44602 ( .A(u_csr_csr_sepc_q[16]), .B(n73501), .Y(n42573) );
  XOR2X1 U44603 ( .A(n50308), .B(n42574), .Y(n50309) );
  XNOR2X1 U44604 ( .A(opcode_pc_w[12]), .B(n44836), .Y(n42574) );
  XOR2X1 U44605 ( .A(n54968), .B(n42575), .Y(n54969) );
  XNOR2X1 U44606 ( .A(opcode_pc_w[11]), .B(opcode_opcode_w[7]), .Y(n42575) );
  XOR2X1 U44607 ( .A(n50372), .B(n42576), .Y(n50373) );
  XNOR2X1 U44608 ( .A(opcode_pc_w[13]), .B(n44836), .Y(n42576) );
  MX2X1 U44609 ( .A(n59085), .B(n59086), .S0(n72803), .Y(n14258) );
  OR2X1 U44610 ( .A(n42577), .B(n28526), .Y(n26931) );
  OR2X1 U44611 ( .A(u_csr_N3162), .B(n51398), .Y(n42577) );
  XOR2X1 U44612 ( .A(n54587), .B(n42578), .Y(n54456) );
  XNOR2X1 U44613 ( .A(opcode_pc_w[4]), .B(opcode_opcode_w[11]), .Y(n42578) );
  XOR2X1 U44614 ( .A(n54511), .B(n42580), .Y(n54512) );
  XNOR2X1 U44615 ( .A(opcode_pc_w[3]), .B(opcode_opcode_w[10]), .Y(n42580) );
  MX2X1 U44616 ( .A(n59076), .B(n59077), .S0(n42712), .Y(n14275) );
  XOR2X1 U44617 ( .A(n43849), .B(n58120), .Y(u_lsu_mem_addr_r[9]) );
  MX2X1 U44618 ( .A(n59072), .B(n59073), .S0(n42652), .Y(n14282) );
  XOR2X1 U44619 ( .A(n44034), .B(n58116), .Y(u_lsu_mem_addr_r[8]) );
  MX2X1 U44620 ( .A(n59065), .B(n59066), .S0(n43798), .Y(n14291) );
  AND2X1 U44621 ( .A(opcode_opcode_w[29]), .B(n58256), .Y(n42581) );
  AND2X1 U44622 ( .A(n50753), .B(writeback_exec_idx_w[0]), .Y(n42582) );
  NOR2X1 U44623 ( .A(opcode_opcode_w[29]), .B(n51991), .Y(n42583) );
  AND2X1 U44624 ( .A(writeback_exec_idx_w[2]), .B(n50720), .Y(n42584) );
  AND2X1 U44625 ( .A(n42584), .B(n50824), .Y(n42585) );
  NOR2X1 U44626 ( .A(n42587), .B(writeback_exec_idx_w[4]), .Y(n42586) );
  OR2X1 U44627 ( .A(writeback_exec_idx_w[0]), .B(n50837), .Y(n42587) );
  AND2X1 U44628 ( .A(writeback_exec_idx_w[0]), .B(n50838), .Y(n42588) );
  AND2X1 U44629 ( .A(writeback_exec_idx_w[3]), .B(writeback_exec_idx_w[4]), 
        .Y(n42589) );
  AND2X1 U44630 ( .A(n42589), .B(writeback_exec_idx_w[0]), .Y(n42590) );
  AND2X1 U44631 ( .A(writeback_exec_idx_w[3]), .B(n42588), .Y(n42591) );
  AND2X1 U44632 ( .A(n42593), .B(writeback_exec_idx_w[2]), .Y(n42592) );
  AND2X1 U44633 ( .A(writeback_exec_idx_w[1]), .B(n50824), .Y(n42593) );
  AND2X1 U44634 ( .A(n42593), .B(n50802), .Y(n42594) );
  NAND2X1 U44635 ( .A(n42596), .B(n42597), .Y(n42595) );
  NOR2X1 U44636 ( .A(n28179), .B(n57427), .Y(n42597) );
  AND2X1 U44637 ( .A(u_muldiv_div_busy_q), .B(n44631), .Y(n42598) );
  AND2X1 U44638 ( .A(n50793), .B(n50824), .Y(n42599) );
  AND2X1 U44639 ( .A(writeback_exec_idx_w[3]), .B(n50838), .Y(n42600) );
  AND2X1 U44640 ( .A(n50838), .B(n39766), .Y(n42601) );
  MX2X1 U44641 ( .A(n59045), .B(n59046), .S0(n43787), .Y(n14323) );
  AND2X1 U44642 ( .A(writeback_exec_idx_w[1]), .B(writeback_exec_idx_w[2]), 
        .Y(n42602) );
  AND2X1 U44643 ( .A(writeback_exec_idx_w[1]), .B(n50802), .Y(n42603) );
  AND2X1 U44644 ( .A(n50819), .B(n50824), .Y(n42604) );
  AND2X1 U44645 ( .A(n50826), .B(n50825), .Y(n42605) );
  MX2X1 U44646 ( .A(n58992), .B(n58993), .S0(n72786), .Y(n14410) );
  MX2X1 U44647 ( .A(n59025), .B(n59026), .S0(n43810), .Y(n14355) );
  MX2X1 U44648 ( .A(n59005), .B(n59006), .S0(n72806), .Y(n14387) );
  AND2X1 U44649 ( .A(n57437), .B(n58521), .Y(n42606) );
  AND2X1 U44650 ( .A(opcode_instr_w_40), .B(n73544), .Y(n42607) );
  AND2X1 U44651 ( .A(opcode_instr_w_35), .B(n57351), .Y(n42608) );
  OR2X1 U44652 ( .A(n42610), .B(n58189), .Y(n58190) );
  AND2X1 U44653 ( .A(u_mmu_itlb_entry_q_4), .B(n42611), .Y(n29681) );
  AND2X1 U44654 ( .A(u_csr_N3161), .B(n8835), .Y(n42611) );
  OR2X1 U44655 ( .A(n58457), .B(n25640), .Y(n58462) );
  OR2X1 U44656 ( .A(n1855), .B(n1849), .Y(n28943) );
  MX2X1 U44657 ( .A(u_mmu_itlb_entry_q[29]), .B(n14), .S0(n58179), .Y(
        mem_i_pc_o[29]) );
  INVX1 U44658 ( .A(n1953), .Y(n47972) );
  INVX1 U44659 ( .A(n42612), .Y(n48094) );
  INVX1 U44660 ( .A(n42613), .Y(n48089) );
  INVX1 U44661 ( .A(n42614), .Y(n61174) );
  INVX1 U44662 ( .A(opcode_instr_w_48), .Y(n57417) );
  NAND2X1 U44663 ( .A(n38492), .B(n46216), .Y(n42615) );
  NAND2X1 U44664 ( .A(n42883), .B(n46049), .Y(n42616) );
  INVX1 U44665 ( .A(n49587), .Y(n42617) );
  INVX1 U44666 ( .A(n42623), .Y(n42618) );
  INVX1 U44667 ( .A(n49587), .Y(n42619) );
  INVX1 U44668 ( .A(n42622), .Y(n42620) );
  INVX1 U44669 ( .A(n42622), .Y(n42621) );
  INVX1 U44670 ( .A(n42818), .Y(n42622) );
  INVX1 U44671 ( .A(n42818), .Y(n42623) );
  INVX1 U44672 ( .A(n49593), .Y(n42624) );
  INVX1 U44673 ( .A(n49593), .Y(n42625) );
  INVX1 U44674 ( .A(n49593), .Y(n42626) );
  INVX1 U44675 ( .A(n49593), .Y(n42627) );
  INVX1 U44676 ( .A(n42624), .Y(n42628) );
  INVX1 U44677 ( .A(n42624), .Y(n42629) );
  INVX1 U44678 ( .A(n42635), .Y(n42630) );
  INVX1 U44679 ( .A(n42634), .Y(n42631) );
  INVX1 U44680 ( .A(n42634), .Y(n42632) );
  INVX1 U44681 ( .A(n42635), .Y(n42633) );
  INVX1 U44682 ( .A(n42633), .Y(n42634) );
  INVX1 U44683 ( .A(n36499), .Y(n42635) );
  INVX1 U44684 ( .A(n38395), .Y(n42636) );
  INVX1 U44685 ( .A(n42630), .Y(n42637) );
  INVX1 U44686 ( .A(n42635), .Y(n42638) );
  INVX1 U44687 ( .A(n42637), .Y(n42639) );
  INVX1 U44688 ( .A(n42637), .Y(n42640) );
  INVX1 U44689 ( .A(n42637), .Y(n42641) );
  INVX1 U44690 ( .A(n42631), .Y(n42642) );
  INVX1 U44691 ( .A(n42642), .Y(n42643) );
  INVX1 U44692 ( .A(n42642), .Y(n42644) );
  NAND2X1 U44693 ( .A(n45535), .B(n42373), .Y(n42645) );
  NAND2X1 U44694 ( .A(n42696), .B(n39449), .Y(n42646) );
  NAND2X1 U44695 ( .A(n42696), .B(n39449), .Y(n42647) );
  INVX1 U44696 ( .A(n43762), .Y(n42648) );
  INVX1 U44697 ( .A(n42660), .Y(n42649) );
  INVX1 U44698 ( .A(n72783), .Y(n42650) );
  INVX1 U44699 ( .A(n42650), .Y(n42651) );
  INVX1 U44700 ( .A(n43762), .Y(n42652) );
  INVX1 U44701 ( .A(n42650), .Y(n42653) );
  INVX1 U44702 ( .A(n42650), .Y(n42654) );
  INVX1 U44703 ( .A(n42648), .Y(n42655) );
  INVX1 U44704 ( .A(n42648), .Y(n42656) );
  INVX1 U44705 ( .A(n42655), .Y(n42657) );
  INVX1 U44706 ( .A(n42655), .Y(n42658) );
  INVX1 U44707 ( .A(n42655), .Y(n42659) );
  INVX1 U44708 ( .A(n42656), .Y(n42660) );
  INVX1 U44709 ( .A(n42656), .Y(n42661) );
  INVX1 U44710 ( .A(opcode_opcode_w[18]), .Y(n42662) );
  INVX1 U44711 ( .A(opcode_opcode_w[18]), .Y(n42663) );
  INVX1 U44712 ( .A(opcode_opcode_w[18]), .Y(n42664) );
  INVX1 U44713 ( .A(opcode_opcode_w[18]), .Y(n42665) );
  INVX1 U44714 ( .A(n42666), .Y(n42667) );
  INVX1 U44715 ( .A(n42666), .Y(n42668) );
  INVX1 U44716 ( .A(n42666), .Y(n42669) );
  INVX1 U44717 ( .A(n40449), .Y(n42670) );
  INVX1 U44718 ( .A(n43019), .Y(n42672) );
  INVX1 U44719 ( .A(n48138), .Y(n42673) );
  INVX1 U44720 ( .A(n42673), .Y(n42674) );
  INVX1 U44721 ( .A(n49610), .Y(n42675) );
  INVX1 U44722 ( .A(n42868), .Y(n42676) );
  INVX1 U44723 ( .A(n49576), .Y(n42677) );
  INVX1 U44724 ( .A(n49576), .Y(n42678) );
  INVX1 U44725 ( .A(n38210), .Y(n42679) );
  INVX1 U44726 ( .A(n38210), .Y(n42680) );
  INVX1 U44727 ( .A(n49576), .Y(n42681) );
  INVX1 U44728 ( .A(n42677), .Y(n42682) );
  INVX1 U44729 ( .A(n42677), .Y(n42683) );
  INVX1 U44730 ( .A(n42677), .Y(n42684) );
  INVX1 U44731 ( .A(n42809), .Y(n42685) );
  INVX1 U44732 ( .A(n42809), .Y(n42686) );
  INVX1 U44733 ( .A(n42809), .Y(n42687) );
  INVX1 U44734 ( .A(opcode_opcode_w[17]), .Y(n42688) );
  INVX1 U44735 ( .A(opcode_opcode_w[17]), .Y(n42689) );
  INVX1 U44736 ( .A(n42780), .Y(n42690) );
  INVX1 U44737 ( .A(n42690), .Y(n42691) );
  INVX1 U44738 ( .A(n42690), .Y(n42692) );
  INVX1 U44739 ( .A(n42697), .Y(n42693) );
  INVX1 U44740 ( .A(n42697), .Y(n42694) );
  INVX1 U44741 ( .A(n42699), .Y(n42695) );
  INVX1 U44742 ( .A(n40498), .Y(n42696) );
  INVX1 U44743 ( .A(n40498), .Y(n42697) );
  INVX1 U44744 ( .A(n38768), .Y(n42698) );
  INVX1 U44745 ( .A(n38768), .Y(n42699) );
  INVX1 U44746 ( .A(n42698), .Y(n42700) );
  INVX1 U44747 ( .A(n43799), .Y(n42701) );
  NAND2X1 U44748 ( .A(n42759), .B(n42748), .Y(n42702) );
  INVX1 U44749 ( .A(n42780), .Y(n42703) );
  INVX1 U44750 ( .A(n42703), .Y(n42704) );
  INVX1 U44751 ( .A(n42703), .Y(n42705) );
  INVX1 U44752 ( .A(n49573), .Y(n42706) );
  INVX1 U44753 ( .A(n49573), .Y(n42707) );
  INVX1 U44754 ( .A(n40444), .Y(n42708) );
  INVX1 U44755 ( .A(n40444), .Y(n42709) );
  INVX1 U44756 ( .A(n42708), .Y(n42710) );
  INVX1 U44757 ( .A(n42710), .Y(n42711) );
  INVX1 U44758 ( .A(n42710), .Y(n42712) );
  INVX1 U44759 ( .A(n42709), .Y(n42713) );
  INVX1 U44760 ( .A(n42713), .Y(n42714) );
  INVX1 U44761 ( .A(n43462), .Y(n42715) );
  INVX1 U44762 ( .A(n43462), .Y(n42716) );
  INVX1 U44763 ( .A(n43462), .Y(n42717) );
  INVX1 U44764 ( .A(n43463), .Y(n42718) );
  INVX1 U44765 ( .A(n43461), .Y(n42719) );
  INVX1 U44766 ( .A(n43461), .Y(n42720) );
  INVX1 U44767 ( .A(n42721), .Y(n42722) );
  INVX1 U44768 ( .A(n42721), .Y(n42723) );
  INVX1 U44769 ( .A(n42721), .Y(n42724) );
  INVX1 U44770 ( .A(opcode_opcode_w[16]), .Y(n42725) );
  INVX1 U44771 ( .A(opcode_opcode_w[16]), .Y(n42726) );
  INVX1 U44772 ( .A(opcode_opcode_w[16]), .Y(n42727) );
  INVX1 U44773 ( .A(n42732), .Y(n42728) );
  INVX1 U44774 ( .A(n42732), .Y(n42729) );
  INVX1 U44775 ( .A(opcode_opcode_w[15]), .Y(n42730) );
  INVX1 U44776 ( .A(opcode_opcode_w[15]), .Y(n42731) );
  INVX1 U44777 ( .A(n42375), .Y(n42733) );
  INVX1 U44778 ( .A(n42733), .Y(n42734) );
  INVX1 U44779 ( .A(n42733), .Y(n42735) );
  INVX1 U44780 ( .A(n42375), .Y(n42736) );
  INVX1 U44781 ( .A(n38739), .Y(n42737) );
  INVX1 U44782 ( .A(n38739), .Y(n42738) );
  INVX1 U44783 ( .A(opcode_opcode_w[20]), .Y(n42739) );
  NAND2X1 U44784 ( .A(n38609), .B(n42771), .Y(n42741) );
  INVX1 U44785 ( .A(n48605), .Y(n42742) );
  INVX1 U44786 ( .A(n48605), .Y(n42743) );
  INVX1 U44787 ( .A(n48605), .Y(n42744) );
  INVX1 U44788 ( .A(n38806), .Y(n42745) );
  INVX1 U44789 ( .A(n38806), .Y(n42746) );
  INVX1 U44790 ( .A(n42750), .Y(n42747) );
  INVX1 U44791 ( .A(n42750), .Y(n42748) );
  INVX1 U44792 ( .A(opcode_opcode_w[24]), .Y(n42749) );
  INVX1 U44793 ( .A(n48612), .Y(n42751) );
  INVX1 U44794 ( .A(n42751), .Y(n42752) );
  INVX1 U44795 ( .A(n42751), .Y(n42753) );
  INVX1 U44796 ( .A(n42856), .Y(n42754) );
  INVX1 U44797 ( .A(n42856), .Y(n42755) );
  INVX1 U44798 ( .A(n42754), .Y(n42756) );
  INVX1 U44799 ( .A(n42755), .Y(n42757) );
  INVX1 U44800 ( .A(n42755), .Y(n42758) );
  INVX1 U44801 ( .A(n42761), .Y(n42759) );
  INVX1 U44802 ( .A(opcode_opcode_w[23]), .Y(n42760) );
  INVX1 U44803 ( .A(opcode_opcode_w[21]), .Y(n42762) );
  INVX1 U44804 ( .A(n42772), .Y(n42764) );
  INVX1 U44805 ( .A(n42773), .Y(n42765) );
  INVX1 U44806 ( .A(n42774), .Y(n42766) );
  INVX1 U44807 ( .A(n42774), .Y(n42767) );
  INVX1 U44808 ( .A(n40607), .Y(n42768) );
  INVX1 U44809 ( .A(n40607), .Y(n42769) );
  INVX1 U44810 ( .A(n42768), .Y(n42770) );
  INVX1 U44811 ( .A(n42768), .Y(n42771) );
  INVX1 U44812 ( .A(n42769), .Y(n42772) );
  INVX1 U44813 ( .A(n42769), .Y(n42773) );
  INVX1 U44814 ( .A(n42769), .Y(n42774) );
  INVX1 U44815 ( .A(n38740), .Y(n42775) );
  INVX1 U44816 ( .A(n38740), .Y(n42776) );
  INVX1 U44817 ( .A(n40107), .Y(n42777) );
  INVX1 U44818 ( .A(n40107), .Y(n42778) );
  INVX1 U44819 ( .A(n40107), .Y(n42779) );
  INVX1 U44820 ( .A(n49605), .Y(n42781) );
  INVX1 U44821 ( .A(n36759), .Y(n42782) );
  INVX1 U44822 ( .A(n36759), .Y(n42783) );
  INVX1 U44823 ( .A(n36759), .Y(n42784) );
  INVX1 U44824 ( .A(n42783), .Y(n42785) );
  INVX1 U44825 ( .A(opcode_opcode_w[19]), .Y(n42786) );
  INVX1 U44826 ( .A(opcode_opcode_w[19]), .Y(n42787) );
  INVX1 U44827 ( .A(opcode_opcode_w[19]), .Y(n42788) );
  INVX1 U44828 ( .A(opcode_opcode_w[19]), .Y(n42789) );
  INVX1 U44829 ( .A(opcode_opcode_w[19]), .Y(n42790) );
  INVX1 U44830 ( .A(n42791), .Y(n42792) );
  INVX1 U44831 ( .A(n42791), .Y(n42793) );
  INVX1 U44832 ( .A(n42791), .Y(n42794) );
  INVX1 U44833 ( .A(n42791), .Y(n42795) );
  NAND2X1 U44834 ( .A(n62905), .B(n45314), .Y(n42796) );
  NAND2X1 U44835 ( .A(n62905), .B(n45314), .Y(n42797) );
  INVX1 U44836 ( .A(n59145), .Y(n42798) );
  INVX1 U44837 ( .A(n59145), .Y(n42799) );
  INVX1 U44838 ( .A(n42805), .Y(n42800) );
  INVX1 U44839 ( .A(n42796), .Y(n42801) );
  INVX1 U44840 ( .A(n42796), .Y(n42802) );
  INVX1 U44841 ( .A(n42797), .Y(n42803) );
  INVX1 U44842 ( .A(n42797), .Y(n42804) );
  INVX1 U44843 ( .A(n64082), .Y(n42805) );
  INVX1 U44844 ( .A(n64082), .Y(n42806) );
  OR2X1 U44845 ( .A(n42807), .B(n42740), .Y(n46326) );
  OR2X1 U44846 ( .A(n42814), .B(n42763), .Y(n42807) );
  OR2X1 U44847 ( .A(n42808), .B(n42688), .Y(n48605) );
  OR2X1 U44848 ( .A(opcode_opcode_w[16]), .B(n42732), .Y(n42808) );
  OR2X1 U44849 ( .A(n46894), .B(n46915), .Y(n72783) );
  XNOR2X1 U44850 ( .A(n41973), .B(n64954), .Y(n64500) );
  XOR2X1 U44851 ( .A(n67546), .B(n42810), .Y(n66884) );
  INVX1 U44852 ( .A(n43583), .Y(n42810) );
  OR2X1 U44853 ( .A(n46626), .B(n45651), .Y(n46428) );
  NAND2X1 U44854 ( .A(n42811), .B(n45293), .Y(n42834) );
  OR2X1 U44855 ( .A(mem_d_resp_tag_i[1]), .B(n42763), .Y(n42811) );
  NOR2X1 U44856 ( .A(n42813), .B(n40378), .Y(n42812) );
  INVX1 U44857 ( .A(n40446), .Y(n42813) );
  XNOR2X1 U44858 ( .A(n59165), .B(n59192), .Y(n42815) );
  OR2X1 U44859 ( .A(n59883), .B(n59882), .Y(n42816) );
  INVX1 U44860 ( .A(n42817), .Y(n59221) );
  AND2X1 U44861 ( .A(n46183), .B(n36708), .Y(n42818) );
  INVX1 U44862 ( .A(n42818), .Y(n49587) );
  OR2X1 U44863 ( .A(n60960), .B(n60961), .Y(n60958) );
  NOR2X1 U44864 ( .A(n42881), .B(n45199), .Y(n42819) );
  OR2X1 U44865 ( .A(n42820), .B(n45870), .Y(n46766) );
  OR2X1 U44866 ( .A(n59496), .B(n36764), .Y(n59497) );
  OR2X1 U44867 ( .A(n59743), .B(n36770), .Y(n59745) );
  OR2X1 U44868 ( .A(n38768), .B(n42768), .Y(n49599) );
  AND2X1 U44869 ( .A(n60243), .B(n40391), .Y(n42822) );
  INVX1 U44870 ( .A(n42822), .Y(n59228) );
  OR2X1 U44871 ( .A(n46696), .B(n45651), .Y(n46759) );
  OR2X1 U44872 ( .A(n45176), .B(n38231), .Y(n49717) );
  AND2X1 U44873 ( .A(n61050), .B(n42823), .Y(n61054) );
  INVX1 U44874 ( .A(n61055), .Y(n42823) );
  AND2X1 U44875 ( .A(n49645), .B(n49644), .Y(n42824) );
  OR2X1 U44876 ( .A(n46364), .B(n46389), .Y(n59226) );
  AND2X1 U44877 ( .A(n59166), .B(n40229), .Y(n42825) );
  INVX1 U44878 ( .A(n38765), .Y(n59737) );
  AND2X1 U44879 ( .A(n42826), .B(n42827), .Y(n46784) );
  AND2X1 U44880 ( .A(n46757), .B(n46756), .Y(n42826) );
  AND2X1 U44881 ( .A(n46765), .B(n46764), .Y(n42827) );
  AND2X1 U44882 ( .A(n40379), .B(n59242), .Y(n42828) );
  INVX1 U44883 ( .A(n42829), .Y(n59322) );
  NOR2X1 U44884 ( .A(n42832), .B(n42831), .Y(n42830) );
  INVX1 U44885 ( .A(n46741), .Y(n42831) );
  OR2X1 U44886 ( .A(n40525), .B(n42690), .Y(n42832) );
  OR2X1 U44887 ( .A(n59474), .B(n59473), .Y(n59475) );
  OR2X1 U44888 ( .A(n59454), .B(n59455), .Y(n59456) );
  OR2X1 U44889 ( .A(n45199), .B(n46927), .Y(n49594) );
  OR2X1 U44890 ( .A(n59724), .B(n59725), .Y(n59729) );
  OR2X1 U44891 ( .A(n42867), .B(n46326), .Y(n49576) );
  OR2X1 U44892 ( .A(n45167), .B(n45166), .Y(n42833) );
  NOR2X1 U44893 ( .A(n42836), .B(n42837), .Y(n42835) );
  AND2X1 U44894 ( .A(n37390), .B(n38728), .Y(n42836) );
  AND2X1 U44895 ( .A(n42181), .B(n60206), .Y(n42837) );
  AND2X1 U44896 ( .A(n59405), .B(n59406), .Y(n42839) );
  INVX1 U44897 ( .A(n42839), .Y(n59467) );
  OR2X1 U44898 ( .A(n59265), .B(n59264), .Y(n59271) );
  INVX1 U44899 ( .A(n42840), .Y(n59211) );
  AND2X1 U44900 ( .A(n61251), .B(n61254), .Y(n42841) );
  NOR2X1 U44901 ( .A(n42844), .B(n42843), .Y(n42842) );
  INVX1 U44902 ( .A(n42842), .Y(n63602) );
  AND2X1 U44903 ( .A(n63334), .B(n63333), .Y(n42843) );
  AND2X1 U44904 ( .A(n63337), .B(n63335), .Y(n42844) );
  INVX1 U44905 ( .A(n38002), .Y(n42845) );
  INVX1 U44906 ( .A(n38002), .Y(n42846) );
  INVX1 U44907 ( .A(n37413), .Y(n42847) );
  INVX1 U44908 ( .A(n26912), .Y(n42848) );
  INVX1 U44909 ( .A(n26912), .Y(n42849) );
  INVX1 U44910 ( .A(n44837), .Y(n42850) );
  INVX1 U44911 ( .A(n42850), .Y(n42851) );
  INVX1 U44912 ( .A(n42850), .Y(n42852) );
  INVX1 U44913 ( .A(n42487), .Y(n42853) );
  INVX1 U44914 ( .A(n42487), .Y(n42854) );
  INVX1 U44915 ( .A(n42487), .Y(n42855) );
  INVX1 U44916 ( .A(n48612), .Y(n42856) );
  INVX1 U44917 ( .A(n42856), .Y(n42857) );
  INVX1 U44918 ( .A(n42224), .Y(n42858) );
  INVX1 U44919 ( .A(n42224), .Y(n42859) );
  INVX1 U44920 ( .A(n42504), .Y(n42860) );
  INVX1 U44921 ( .A(n42504), .Y(n42861) );
  INVX1 U44922 ( .A(n42504), .Y(n42862) );
  INVX1 U44923 ( .A(n39449), .Y(n42863) );
  INVX1 U44924 ( .A(n40248), .Y(n42864) );
  INVX1 U44925 ( .A(n40249), .Y(n42865) );
  INVX1 U44926 ( .A(n38659), .Y(n42866) );
  INVX1 U44927 ( .A(n38659), .Y(n42867) );
  INVX1 U44928 ( .A(n38659), .Y(n42868) );
  INVX1 U44929 ( .A(n42370), .Y(n42869) );
  INVX1 U44930 ( .A(n42370), .Y(n42870) );
  INVX1 U44931 ( .A(n42370), .Y(n42871) );
  INVX1 U44932 ( .A(n42292), .Y(n42872) );
  INVX1 U44933 ( .A(n42292), .Y(n42873) );
  INVX1 U44934 ( .A(n42292), .Y(n42874) );
  INVX1 U44935 ( .A(n42467), .Y(n42875) );
  INVX1 U44936 ( .A(n40843), .Y(n42876) );
  INVX1 U44937 ( .A(n40843), .Y(n42877) );
  INVX1 U44938 ( .A(n40843), .Y(n42878) );
  INVX1 U44939 ( .A(n42362), .Y(n42879) );
  INVX1 U44940 ( .A(n42362), .Y(n42880) );
  INVX1 U44941 ( .A(n42467), .Y(n42881) );
  INVX1 U44942 ( .A(n36600), .Y(n42882) );
  INVX1 U44943 ( .A(n36608), .Y(n42883) );
  INVX1 U44944 ( .A(n49699), .Y(n42884) );
  INVX1 U44945 ( .A(n40505), .Y(n42885) );
  INVX1 U44946 ( .A(n49621), .Y(n42886) );
  INVX1 U44947 ( .A(n49621), .Y(n42887) );
  INVX1 U44948 ( .A(n42884), .Y(n42888) );
  INVX1 U44949 ( .A(n38717), .Y(n42889) );
  INVX1 U44950 ( .A(n38717), .Y(n42890) );
  INVX1 U44951 ( .A(n42481), .Y(n42891) );
  INVX1 U44952 ( .A(n42481), .Y(n42892) );
  INVX1 U44953 ( .A(n42222), .Y(n42893) );
  INVX1 U44954 ( .A(n42222), .Y(n42894) );
  INVX1 U44955 ( .A(n42821), .Y(n42895) );
  INVX1 U44956 ( .A(n42821), .Y(n42896) );
  INVX1 U44957 ( .A(n49717), .Y(n42897) );
  INVX1 U44958 ( .A(n42897), .Y(n42898) );
  INVX1 U44959 ( .A(n42897), .Y(n42899) );
  NAND2X1 U44960 ( .A(n46412), .B(n46404), .Y(n42900) );
  NAND2X1 U44961 ( .A(n40590), .B(n46309), .Y(n42901) );
  INVX1 U44962 ( .A(n42147), .Y(n42902) );
  INVX1 U44963 ( .A(n42147), .Y(n42903) );
  INVX1 U44964 ( .A(n42223), .Y(n42904) );
  INVX1 U44965 ( .A(n42223), .Y(n42905) );
  INVX1 U44966 ( .A(n42223), .Y(n42906) );
  NAND2X1 U44967 ( .A(n42146), .B(n40404), .Y(n42907) );
  NAND2X1 U44968 ( .A(n42146), .B(n40404), .Y(n42908) );
  NAND2X1 U44969 ( .A(n36733), .B(n40447), .Y(n42909) );
  NAND2X1 U44970 ( .A(n40594), .B(n40447), .Y(n42910) );
  NAND2X1 U44971 ( .A(n40499), .B(n46736), .Y(n42911) );
  INVX1 U44972 ( .A(n38085), .Y(n42912) );
  INVX1 U44973 ( .A(n41740), .Y(n42913) );
  INVX1 U44974 ( .A(n41741), .Y(n42914) );
  INVX1 U44975 ( .A(n41741), .Y(n42915) );
  INVX1 U44976 ( .A(n41741), .Y(n42916) );
  INVX1 U44977 ( .A(n41742), .Y(n42917) );
  INVX1 U44978 ( .A(n41742), .Y(n42918) );
  INVX1 U44979 ( .A(n41742), .Y(n42919) );
  INVX1 U44980 ( .A(n50017), .Y(n42920) );
  INVX1 U44981 ( .A(n50017), .Y(n42921) );
  INVX1 U44982 ( .A(n42920), .Y(n42922) );
  INVX1 U44983 ( .A(n42920), .Y(n42923) );
  INVX1 U44984 ( .A(n42920), .Y(n42924) );
  INVX1 U44985 ( .A(n42921), .Y(n42925) );
  INVX1 U44986 ( .A(n42921), .Y(n42926) );
  INVX1 U44987 ( .A(n42921), .Y(n42927) );
  INVX1 U44988 ( .A(n42921), .Y(n42928) );
  INVX1 U44989 ( .A(n42579), .Y(n42929) );
  INVX1 U44990 ( .A(n42579), .Y(n42930) );
  INVX1 U44991 ( .A(n42579), .Y(n42931) );
  INVX1 U44992 ( .A(n42258), .Y(n42932) );
  INVX1 U44993 ( .A(n42258), .Y(n42933) );
  INVX1 U44994 ( .A(n42258), .Y(n42934) );
  NAND2X1 U44995 ( .A(opcode_instr_w[10]), .B(n50668), .Y(n42935) );
  NAND2X1 U44996 ( .A(opcode_instr_w[10]), .B(n50668), .Y(n42936) );
  NAND2X1 U44997 ( .A(n50697), .B(n50696), .Y(n42937) );
  NAND2X1 U44998 ( .A(n50697), .B(n50696), .Y(n42938) );
  INVX1 U44999 ( .A(n40680), .Y(n42939) );
  INVX1 U45000 ( .A(n40680), .Y(n42940) );
  INVX1 U45001 ( .A(n40680), .Y(n42941) );
  INVX1 U45002 ( .A(n362), .Y(n42942) );
  INVX1 U45003 ( .A(n42942), .Y(n42943) );
  NAND2X1 U45004 ( .A(n42315), .B(n73571), .Y(n42944) );
  NAND2X1 U45005 ( .A(n42315), .B(n73571), .Y(n42945) );
  NAND2X1 U45006 ( .A(n42310), .B(n73573), .Y(n42946) );
  INVX1 U45007 ( .A(n40690), .Y(n42947) );
  INVX1 U45008 ( .A(n40689), .Y(n42948) );
  INVX1 U45009 ( .A(n40691), .Y(n42949) );
  INVX1 U45010 ( .A(n58222), .Y(n42950) );
  INVX1 U45011 ( .A(n42950), .Y(n42951) );
  INVX1 U45012 ( .A(n42950), .Y(n42952) );
  INVX1 U45013 ( .A(n42950), .Y(n42953) );
  INVX1 U45014 ( .A(n58251), .Y(n42954) );
  INVX1 U45015 ( .A(n42954), .Y(n42955) );
  INVX1 U45016 ( .A(n42954), .Y(n42956) );
  INVX1 U45017 ( .A(n42954), .Y(n42957) );
  INVX1 U45018 ( .A(n15847), .Y(n42958) );
  INVX1 U45019 ( .A(n42958), .Y(n42959) );
  INVX1 U45020 ( .A(n42958), .Y(n42960) );
  INVX1 U45021 ( .A(n73503), .Y(n42961) );
  INVX1 U45022 ( .A(n42961), .Y(n42962) );
  INVX1 U45023 ( .A(n42131), .Y(n42963) );
  INVX1 U45024 ( .A(n42131), .Y(n42964) );
  INVX1 U45025 ( .A(n42135), .Y(n42965) );
  INVX1 U45026 ( .A(n42135), .Y(n42966) );
  INVX1 U45027 ( .A(n42135), .Y(n42967) );
  INVX1 U45028 ( .A(n37554), .Y(n42968) );
  INVX1 U45029 ( .A(n37554), .Y(n42969) );
  INVX1 U45030 ( .A(n37554), .Y(n42970) );
  OR2X1 U45031 ( .A(n15749), .B(n57298), .Y(n42971) );
  OR2X1 U45032 ( .A(n15749), .B(n57298), .Y(n42972) );
  INVX1 U45033 ( .A(n29961), .Y(n42973) );
  INVX1 U45034 ( .A(n42973), .Y(n42974) );
  INVX1 U45035 ( .A(n42973), .Y(n42975) );
  INVX1 U45036 ( .A(n42973), .Y(n42976) );
  INVX1 U45037 ( .A(n37587), .Y(n42977) );
  INVX1 U45038 ( .A(n37587), .Y(n42978) );
  INVX1 U45039 ( .A(n37587), .Y(n42979) );
  NAND2X1 U45040 ( .A(n42453), .B(n43607), .Y(n42980) );
  NAND2X1 U45041 ( .A(n42453), .B(n43607), .Y(n42981) );
  INVX1 U45042 ( .A(n41738), .Y(n42982) );
  INVX1 U45043 ( .A(n41738), .Y(n42983) );
  NAND2X1 U45044 ( .A(n43420), .B(n58542), .Y(n42984) );
  NAND2X1 U45045 ( .A(n43420), .B(n58542), .Y(n42985) );
  INVX1 U45046 ( .A(n37539), .Y(n42986) );
  INVX1 U45047 ( .A(n37539), .Y(n42987) );
  INVX1 U45048 ( .A(n37539), .Y(n42988) );
  INVX1 U45049 ( .A(n360), .Y(n42989) );
  INVX1 U45050 ( .A(n42989), .Y(n42990) );
  INVX1 U45051 ( .A(n42989), .Y(n42991) );
  INVX1 U45052 ( .A(n42185), .Y(n42992) );
  INVX1 U45053 ( .A(n42185), .Y(n42993) );
  INVX1 U45054 ( .A(n42185), .Y(n42994) );
  INVX1 U45055 ( .A(n42184), .Y(n42995) );
  INVX1 U45056 ( .A(n42184), .Y(n42996) );
  INVX1 U45057 ( .A(n42184), .Y(n42997) );
  INVX1 U45058 ( .A(n42187), .Y(n42998) );
  INVX1 U45059 ( .A(n42187), .Y(n42999) );
  INVX1 U45060 ( .A(n42188), .Y(n43000) );
  INVX1 U45061 ( .A(n42188), .Y(n43001) );
  INVX1 U45062 ( .A(n42216), .Y(n43002) );
  INVX1 U45063 ( .A(n42216), .Y(n43003) );
  INVX1 U45064 ( .A(n42216), .Y(n43004) );
  INVX1 U45065 ( .A(n15408), .Y(n43005) );
  INVX1 U45066 ( .A(n43005), .Y(n43006) );
  INVX1 U45067 ( .A(n43005), .Y(n43007) );
  NAND2X1 U45068 ( .A(n73573), .B(n73572), .Y(n43008) );
  INVX1 U45069 ( .A(n37341), .Y(n43009) );
  INVX1 U45070 ( .A(n37341), .Y(n43010) );
  INVX1 U45071 ( .A(n37341), .Y(n43011) );
  INVX1 U45072 ( .A(n43012), .Y(n43013) );
  INVX1 U45073 ( .A(n43012), .Y(n43014) );
  INVX1 U45074 ( .A(n40449), .Y(n43015) );
  INVX1 U45075 ( .A(n43018), .Y(n43016) );
  INVX1 U45076 ( .A(n48212), .Y(n43017) );
  INVX1 U45077 ( .A(n43015), .Y(n43018) );
  INVX1 U45078 ( .A(n48138), .Y(n43019) );
  INVX1 U45079 ( .A(n49715), .Y(n43020) );
  INVX1 U45080 ( .A(n43024), .Y(n43021) );
  INVX1 U45081 ( .A(n43024), .Y(n43022) );
  INVX1 U45082 ( .A(n43024), .Y(n43023) );
  INVX1 U45083 ( .A(n49806), .Y(n43024) );
  INVX1 U45084 ( .A(n49806), .Y(n43025) );
  INVX1 U45085 ( .A(n49806), .Y(n43026) );
  INVX1 U45086 ( .A(n45317), .Y(n43027) );
  INVX1 U45087 ( .A(n45317), .Y(n43028) );
  INVX1 U45088 ( .A(n47624), .Y(n43029) );
  INVX1 U45089 ( .A(n47624), .Y(n43030) );
  INVX1 U45090 ( .A(n47624), .Y(n43031) );
  INVX1 U45091 ( .A(n43035), .Y(n43032) );
  INVX1 U45092 ( .A(n43035), .Y(n43033) );
  INVX1 U45093 ( .A(n43035), .Y(n43034) );
  INVX1 U45094 ( .A(n42158), .Y(n43035) );
  INVX1 U45095 ( .A(n45324), .Y(n43036) );
  INVX1 U45096 ( .A(n45324), .Y(n43037) );
  INVX1 U45097 ( .A(n43041), .Y(n43038) );
  INVX1 U45098 ( .A(n43041), .Y(n43039) );
  INVX1 U45099 ( .A(n43041), .Y(n43040) );
  INVX1 U45100 ( .A(n40023), .Y(n43041) );
  INVX1 U45101 ( .A(n57609), .Y(n43042) );
  INVX1 U45102 ( .A(n57609), .Y(n43043) );
  INVX1 U45103 ( .A(n43046), .Y(n43044) );
  INVX1 U45104 ( .A(n43046), .Y(n43045) );
  INVX1 U45105 ( .A(n39630), .Y(n43046) );
  INVX1 U45106 ( .A(n45347), .Y(n43047) );
  INVX1 U45107 ( .A(n45347), .Y(n43048) );
  INVX1 U45108 ( .A(n45350), .Y(n43049) );
  INVX1 U45109 ( .A(n45350), .Y(n43050) );
  INVX1 U45110 ( .A(n48386), .Y(n43051) );
  INVX1 U45111 ( .A(n48386), .Y(n43052) );
  INVX1 U45112 ( .A(n47668), .Y(n43053) );
  INVX1 U45113 ( .A(n57625), .Y(n43054) );
  INVX1 U45114 ( .A(n57625), .Y(n43055) );
  INVX1 U45115 ( .A(n43059), .Y(n43056) );
  INVX1 U45116 ( .A(n43059), .Y(n43057) );
  INVX1 U45117 ( .A(n43059), .Y(n43058) );
  INVX1 U45118 ( .A(n39620), .Y(n43059) );
  INVX1 U45119 ( .A(n48373), .Y(n43060) );
  INVX1 U45120 ( .A(n48373), .Y(n43061) );
  INVX1 U45121 ( .A(n48373), .Y(n43062) );
  INVX1 U45122 ( .A(n57604), .Y(n43063) );
  INVX1 U45123 ( .A(n57604), .Y(n43064) );
  INVX1 U45124 ( .A(n57604), .Y(n43065) );
  INVX1 U45125 ( .A(n45363), .Y(n43066) );
  INVX1 U45126 ( .A(n45363), .Y(n43067) );
  INVX1 U45127 ( .A(n45363), .Y(n43068) );
  INVX1 U45128 ( .A(n48357), .Y(n43069) );
  INVX1 U45129 ( .A(n48357), .Y(n43070) );
  INVX1 U45130 ( .A(n37396), .Y(n43071) );
  INVX1 U45131 ( .A(n37396), .Y(n43072) );
  INVX1 U45132 ( .A(n37396), .Y(n43073) );
  INVX1 U45133 ( .A(n47618), .Y(n43074) );
  INVX1 U45134 ( .A(n47618), .Y(n43075) );
  INVX1 U45135 ( .A(n47618), .Y(n43076) );
  INVX1 U45136 ( .A(n43079), .Y(n43077) );
  INVX1 U45137 ( .A(n43079), .Y(n43078) );
  INVX1 U45138 ( .A(n37664), .Y(n43079) );
  INVX1 U45139 ( .A(n62903), .Y(n43080) );
  INVX1 U45140 ( .A(n62903), .Y(n43081) );
  INVX1 U45141 ( .A(n62903), .Y(n43082) );
  INVX1 U45142 ( .A(n43085), .Y(n43083) );
  INVX1 U45143 ( .A(n43085), .Y(n43084) );
  INVX1 U45144 ( .A(n37666), .Y(n43085) );
  INVX1 U45145 ( .A(n37788), .Y(n43086) );
  INVX1 U45146 ( .A(n37788), .Y(n43087) );
  INVX1 U45147 ( .A(n37788), .Y(n43088) );
  INVX1 U45148 ( .A(n43091), .Y(n43089) );
  INVX1 U45149 ( .A(n43091), .Y(n43090) );
  INVX1 U45150 ( .A(n37670), .Y(n43091) );
  INVX1 U45151 ( .A(n37782), .Y(n43092) );
  INVX1 U45152 ( .A(n37782), .Y(n43093) );
  INVX1 U45153 ( .A(n37782), .Y(n43094) );
  INVX1 U45154 ( .A(n43097), .Y(n43095) );
  INVX1 U45155 ( .A(n43097), .Y(n43096) );
  INVX1 U45156 ( .A(n37671), .Y(n43097) );
  INVX1 U45157 ( .A(n37786), .Y(n43098) );
  INVX1 U45158 ( .A(n37786), .Y(n43099) );
  INVX1 U45159 ( .A(n37786), .Y(n43100) );
  INVX1 U45160 ( .A(writeback_exec_value_w[8]), .Y(n43101) );
  INVX1 U45161 ( .A(writeback_exec_value_w[8]), .Y(n43102) );
  INVX1 U45162 ( .A(n37790), .Y(n43103) );
  INVX1 U45163 ( .A(n37790), .Y(n43104) );
  INVX1 U45164 ( .A(n37790), .Y(n43105) );
  INVX1 U45165 ( .A(writeback_exec_value_w[7]), .Y(n43106) );
  INVX1 U45166 ( .A(writeback_exec_value_w[7]), .Y(n43107) );
  INVX1 U45167 ( .A(n48676), .Y(n43108) );
  INVX1 U45168 ( .A(n48676), .Y(n43109) );
  INVX1 U45169 ( .A(n48676), .Y(n43110) );
  INVX1 U45170 ( .A(n43113), .Y(n43111) );
  INVX1 U45171 ( .A(n43113), .Y(n43112) );
  INVX1 U45172 ( .A(n37667), .Y(n43113) );
  INVX1 U45173 ( .A(n48516), .Y(n43114) );
  INVX1 U45174 ( .A(n48516), .Y(n43115) );
  INVX1 U45175 ( .A(n48516), .Y(n43116) );
  INVX1 U45176 ( .A(n43119), .Y(n43117) );
  INVX1 U45177 ( .A(n43119), .Y(n43118) );
  INVX1 U45178 ( .A(n37668), .Y(n43119) );
  INVX1 U45179 ( .A(n37787), .Y(n43120) );
  INVX1 U45180 ( .A(n37787), .Y(n43121) );
  INVX1 U45181 ( .A(n37787), .Y(n43122) );
  INVX1 U45182 ( .A(writeback_exec_value_w[9]), .Y(n43123) );
  INVX1 U45183 ( .A(writeback_exec_value_w[9]), .Y(n43124) );
  INVX1 U45184 ( .A(n37783), .Y(n43125) );
  INVX1 U45185 ( .A(n37783), .Y(n43126) );
  INVX1 U45186 ( .A(n37783), .Y(n43127) );
  INVX1 U45187 ( .A(writeback_exec_value_w[10]), .Y(n43128) );
  INVX1 U45188 ( .A(writeback_exec_value_w[10]), .Y(n43129) );
  INVX1 U45189 ( .A(n37784), .Y(n43130) );
  INVX1 U45190 ( .A(n37784), .Y(n43131) );
  INVX1 U45191 ( .A(n37784), .Y(n43132) );
  INVX1 U45192 ( .A(n43135), .Y(n43133) );
  INVX1 U45193 ( .A(n43135), .Y(n43134) );
  INVX1 U45194 ( .A(n37676), .Y(n43135) );
  INVX1 U45195 ( .A(n37785), .Y(n43136) );
  INVX1 U45196 ( .A(n37785), .Y(n43137) );
  INVX1 U45197 ( .A(n37785), .Y(n43138) );
  INVX1 U45198 ( .A(n43141), .Y(n43139) );
  INVX1 U45199 ( .A(n43141), .Y(n43140) );
  INVX1 U45200 ( .A(n37677), .Y(n43141) );
  INVX1 U45201 ( .A(n37789), .Y(n43142) );
  INVX1 U45202 ( .A(n37789), .Y(n43143) );
  INVX1 U45203 ( .A(n37789), .Y(n43144) );
  INVX1 U45204 ( .A(n43147), .Y(n43145) );
  INVX1 U45205 ( .A(n43147), .Y(n43146) );
  INVX1 U45206 ( .A(n37678), .Y(n43147) );
  INVX1 U45207 ( .A(n37795), .Y(n43148) );
  INVX1 U45208 ( .A(n37795), .Y(n43149) );
  INVX1 U45209 ( .A(n37795), .Y(n43150) );
  INVX1 U45210 ( .A(n43153), .Y(n43151) );
  INVX1 U45211 ( .A(n43153), .Y(n43152) );
  INVX1 U45212 ( .A(n37679), .Y(n43153) );
  INVX1 U45213 ( .A(n37792), .Y(n43154) );
  INVX1 U45214 ( .A(n37792), .Y(n43155) );
  INVX1 U45215 ( .A(n37792), .Y(n43156) );
  INVX1 U45216 ( .A(n43159), .Y(n43157) );
  INVX1 U45217 ( .A(n43159), .Y(n43158) );
  INVX1 U45218 ( .A(n37680), .Y(n43159) );
  INVX1 U45219 ( .A(n37793), .Y(n43160) );
  INVX1 U45220 ( .A(n37793), .Y(n43161) );
  INVX1 U45221 ( .A(n37793), .Y(n43162) );
  INVX1 U45222 ( .A(n43165), .Y(n43163) );
  INVX1 U45223 ( .A(n43165), .Y(n43164) );
  INVX1 U45224 ( .A(n37681), .Y(n43165) );
  INVX1 U45225 ( .A(n37354), .Y(n43166) );
  INVX1 U45226 ( .A(n37354), .Y(n43167) );
  INVX1 U45227 ( .A(n37354), .Y(n43168) );
  INVX1 U45228 ( .A(writeback_exec_value_w[19]), .Y(n43169) );
  INVX1 U45229 ( .A(writeback_exec_value_w[19]), .Y(n43170) );
  INVX1 U45230 ( .A(n40844), .Y(n43171) );
  INVX1 U45231 ( .A(n40844), .Y(n43172) );
  INVX1 U45232 ( .A(n40844), .Y(n43173) );
  INVX1 U45233 ( .A(writeback_exec_value_w[20]), .Y(n43174) );
  INVX1 U45234 ( .A(writeback_exec_value_w[20]), .Y(n43175) );
  INVX1 U45235 ( .A(n40845), .Y(n43176) );
  INVX1 U45236 ( .A(n40845), .Y(n43177) );
  INVX1 U45237 ( .A(n40845), .Y(n43178) );
  INVX1 U45238 ( .A(n43181), .Y(n43179) );
  INVX1 U45239 ( .A(n43181), .Y(n43180) );
  INVX1 U45240 ( .A(n37682), .Y(n43181) );
  INVX1 U45241 ( .A(n43184), .Y(n43182) );
  INVX1 U45242 ( .A(n43184), .Y(n43183) );
  INVX1 U45243 ( .A(n53762), .Y(n43184) );
  INVX1 U45244 ( .A(n43187), .Y(n43185) );
  INVX1 U45245 ( .A(n43187), .Y(n43186) );
  INVX1 U45246 ( .A(n37683), .Y(n43187) );
  INVX1 U45247 ( .A(n43190), .Y(n43188) );
  INVX1 U45248 ( .A(n43190), .Y(n43189) );
  INVX1 U45249 ( .A(n53889), .Y(n43190) );
  INVX1 U45250 ( .A(n43193), .Y(n43191) );
  INVX1 U45251 ( .A(n43193), .Y(n43192) );
  INVX1 U45252 ( .A(n37684), .Y(n43193) );
  INVX1 U45253 ( .A(n40941), .Y(n43194) );
  INVX1 U45254 ( .A(n40941), .Y(n43195) );
  INVX1 U45255 ( .A(n40941), .Y(n43196) );
  INVX1 U45256 ( .A(writeback_exec_value_w[24]), .Y(n43197) );
  INVX1 U45257 ( .A(writeback_exec_value_w[24]), .Y(n43198) );
  INVX1 U45258 ( .A(n40939), .Y(n43199) );
  INVX1 U45259 ( .A(n40939), .Y(n43200) );
  INVX1 U45260 ( .A(n40939), .Y(n43201) );
  INVX1 U45261 ( .A(writeback_exec_value_w[25]), .Y(n43202) );
  INVX1 U45262 ( .A(writeback_exec_value_w[25]), .Y(n43203) );
  INVX1 U45263 ( .A(n37794), .Y(n43204) );
  INVX1 U45264 ( .A(n37794), .Y(n43205) );
  INVX1 U45265 ( .A(n37794), .Y(n43206) );
  INVX1 U45266 ( .A(n37406), .Y(n43207) );
  INVX1 U45267 ( .A(n37406), .Y(n43208) );
  INVX1 U45268 ( .A(n37406), .Y(n43209) );
  INVX1 U45269 ( .A(n43212), .Y(n43210) );
  INVX1 U45270 ( .A(n43212), .Y(n43211) );
  INVX1 U45271 ( .A(n55947), .Y(n43212) );
  INVX1 U45272 ( .A(n43216), .Y(n43213) );
  INVX1 U45273 ( .A(n43216), .Y(n43214) );
  INVX1 U45274 ( .A(n43216), .Y(n43215) );
  INVX1 U45275 ( .A(n43219), .Y(n43217) );
  INVX1 U45276 ( .A(n43219), .Y(n43218) );
  INVX1 U45277 ( .A(n56124), .Y(n43219) );
  INVX1 U45278 ( .A(n43222), .Y(n43220) );
  INVX1 U45279 ( .A(n43222), .Y(n43221) );
  INVX1 U45280 ( .A(n37685), .Y(n43222) );
  INVX1 U45281 ( .A(n40940), .Y(n43223) );
  INVX1 U45282 ( .A(n40940), .Y(n43224) );
  INVX1 U45283 ( .A(n40940), .Y(n43225) );
  INVX1 U45284 ( .A(n43228), .Y(n43226) );
  INVX1 U45285 ( .A(n43228), .Y(n43227) );
  INVX1 U45286 ( .A(n37686), .Y(n43228) );
  INVX1 U45287 ( .A(n37355), .Y(n43229) );
  INVX1 U45288 ( .A(n37355), .Y(n43230) );
  INVX1 U45289 ( .A(n37355), .Y(n43231) );
  INVX1 U45290 ( .A(n43235), .Y(n43232) );
  INVX1 U45291 ( .A(n43235), .Y(n43233) );
  INVX1 U45292 ( .A(n43235), .Y(n43234) );
  INVX1 U45293 ( .A(n43238), .Y(n43236) );
  INVX1 U45294 ( .A(n43238), .Y(n43237) );
  INVX1 U45295 ( .A(n42136), .Y(n43238) );
  INVX1 U45296 ( .A(n43241), .Y(n43239) );
  INVX1 U45297 ( .A(n43241), .Y(n43240) );
  INVX1 U45298 ( .A(n56578), .Y(n43241) );
  INVX1 U45299 ( .A(n56578), .Y(n43242) );
  INVX1 U45300 ( .A(n54405), .Y(n43243) );
  INVX1 U45301 ( .A(n54405), .Y(n43244) );
  INVX1 U45302 ( .A(n54405), .Y(n43245) );
  INVX1 U45303 ( .A(n57240), .Y(n43246) );
  INVX1 U45304 ( .A(n57240), .Y(n43247) );
  INVX1 U45305 ( .A(n57240), .Y(n43248) );
  INVX1 U45306 ( .A(n43251), .Y(n43249) );
  INVX1 U45307 ( .A(n43251), .Y(n43250) );
  INVX1 U45308 ( .A(n56590), .Y(n43251) );
  INVX1 U45309 ( .A(n56590), .Y(n43252) );
  INVX1 U45310 ( .A(n43255), .Y(n43253) );
  INVX1 U45311 ( .A(n43255), .Y(n43254) );
  INVX1 U45312 ( .A(n42137), .Y(n43255) );
  INVX1 U45313 ( .A(n54418), .Y(n43256) );
  INVX1 U45314 ( .A(n54418), .Y(n43257) );
  INVX1 U45315 ( .A(n54418), .Y(n43258) );
  INVX1 U45316 ( .A(n57254), .Y(n43259) );
  INVX1 U45317 ( .A(n57254), .Y(n43260) );
  INVX1 U45318 ( .A(n48452), .Y(n43261) );
  INVX1 U45319 ( .A(n48452), .Y(n43262) );
  INVX1 U45320 ( .A(n48452), .Y(n43263) );
  INVX1 U45321 ( .A(n43266), .Y(n43264) );
  INVX1 U45322 ( .A(n43266), .Y(n43265) );
  INVX1 U45323 ( .A(n37669), .Y(n43266) );
  INVX1 U45324 ( .A(n42433), .Y(n43267) );
  INVX1 U45325 ( .A(n42433), .Y(n43268) );
  INVX1 U45326 ( .A(n42433), .Y(n43269) );
  INVX1 U45327 ( .A(n43272), .Y(n43270) );
  INVX1 U45328 ( .A(n43272), .Y(n43271) );
  INVX1 U45329 ( .A(n57131), .Y(n43272) );
  INVX1 U45330 ( .A(n43275), .Y(n43273) );
  INVX1 U45331 ( .A(n43275), .Y(n43274) );
  INVX1 U45332 ( .A(n57144), .Y(n43275) );
  INVX1 U45333 ( .A(n43278), .Y(n43276) );
  INVX1 U45334 ( .A(n43278), .Y(n43277) );
  INVX1 U45335 ( .A(n57209), .Y(n43278) );
  INVX1 U45336 ( .A(n40942), .Y(n43279) );
  INVX1 U45337 ( .A(n40942), .Y(n43280) );
  INVX1 U45338 ( .A(n40942), .Y(n43281) );
  INVX1 U45339 ( .A(n43285), .Y(n43282) );
  INVX1 U45340 ( .A(n43285), .Y(n43283) );
  INVX1 U45341 ( .A(n43285), .Y(n43284) );
  INVX1 U45342 ( .A(n57234), .Y(n43285) );
  INVX1 U45343 ( .A(n42595), .Y(n43286) );
  INVX1 U45344 ( .A(n42595), .Y(n43287) );
  INVX1 U45345 ( .A(n42595), .Y(n43288) );
  INVX1 U45346 ( .A(n42268), .Y(n43289) );
  INVX1 U45347 ( .A(n42268), .Y(n43290) );
  INVX1 U45348 ( .A(n42268), .Y(n43291) );
  INVX1 U45349 ( .A(n42447), .Y(n43292) );
  INVX1 U45350 ( .A(n42447), .Y(n43293) );
  INVX1 U45351 ( .A(n42447), .Y(n43294) );
  INVX1 U45352 ( .A(n42583), .Y(n43295) );
  INVX1 U45353 ( .A(n42583), .Y(n43296) );
  INVX1 U45354 ( .A(n42583), .Y(n43297) );
  INVX1 U45355 ( .A(n37410), .Y(n43298) );
  INVX1 U45356 ( .A(n37410), .Y(n43299) );
  INVX1 U45357 ( .A(n37410), .Y(n43300) );
  INVX1 U45358 ( .A(n37411), .Y(n43301) );
  INVX1 U45359 ( .A(n37411), .Y(n43302) );
  INVX1 U45360 ( .A(n37411), .Y(n43303) );
  INVX1 U45361 ( .A(n42521), .Y(n43304) );
  INVX1 U45362 ( .A(n42521), .Y(n43305) );
  INVX1 U45363 ( .A(n42521), .Y(n43306) );
  INVX1 U45364 ( .A(n43310), .Y(n43307) );
  INVX1 U45365 ( .A(n43310), .Y(n43308) );
  INVX1 U45366 ( .A(n43310), .Y(n43309) );
  INVX1 U45367 ( .A(n42596), .Y(n43310) );
  INVX1 U45368 ( .A(n37409), .Y(n43311) );
  INVX1 U45369 ( .A(n37409), .Y(n43312) );
  INVX1 U45370 ( .A(n37409), .Y(n43313) );
  INVX1 U45371 ( .A(n38002), .Y(n43314) );
  INVX1 U45372 ( .A(n43318), .Y(n43315) );
  INVX1 U45373 ( .A(n43318), .Y(n43316) );
  INVX1 U45374 ( .A(n43318), .Y(n43317) );
  INVX1 U45375 ( .A(n57280), .Y(n43318) );
  INVX1 U45376 ( .A(n57280), .Y(n43319) );
  INVX1 U45377 ( .A(n42263), .Y(n43320) );
  INVX1 U45378 ( .A(n42263), .Y(n43321) );
  INVX1 U45379 ( .A(n42263), .Y(n43322) );
  INVX1 U45380 ( .A(n42426), .Y(n43323) );
  INVX1 U45381 ( .A(n42426), .Y(n43324) );
  INVX1 U45382 ( .A(n42426), .Y(n43325) );
  INVX1 U45383 ( .A(n42427), .Y(n43326) );
  INVX1 U45384 ( .A(n42427), .Y(n43327) );
  INVX1 U45385 ( .A(n42427), .Y(n43328) );
  INVX1 U45386 ( .A(n37791), .Y(n43329) );
  INVX1 U45387 ( .A(n37791), .Y(n43330) );
  INVX1 U45388 ( .A(n37791), .Y(n43331) );
  INVX1 U45389 ( .A(n43334), .Y(n43332) );
  INVX1 U45390 ( .A(n43334), .Y(n43333) );
  INVX1 U45391 ( .A(n37687), .Y(n43334) );
  INVX1 U45392 ( .A(n43337), .Y(n43335) );
  INVX1 U45393 ( .A(n43337), .Y(n43336) );
  INVX1 U45394 ( .A(n37665), .Y(n43337) );
  INVX1 U45395 ( .A(n43341), .Y(n43338) );
  INVX1 U45396 ( .A(n43341), .Y(n43339) );
  INVX1 U45397 ( .A(n43341), .Y(n43340) );
  INVX1 U45398 ( .A(n41791), .Y(n43341) );
  INVX1 U45399 ( .A(n37398), .Y(n43342) );
  INVX1 U45400 ( .A(n37398), .Y(n43343) );
  INVX1 U45401 ( .A(n37398), .Y(n43344) );
  INVX1 U45402 ( .A(n43348), .Y(n43345) );
  INVX1 U45403 ( .A(n43348), .Y(n43346) );
  INVX1 U45404 ( .A(n43348), .Y(n43347) );
  INVX1 U45405 ( .A(n41782), .Y(n43348) );
  INVX1 U45406 ( .A(n47621), .Y(n43349) );
  INVX1 U45407 ( .A(n47621), .Y(n43350) );
  INVX1 U45408 ( .A(n43353), .Y(n43351) );
  INVX1 U45409 ( .A(n43353), .Y(n43352) );
  INVX1 U45410 ( .A(n42165), .Y(n43353) );
  INVX1 U45411 ( .A(n43357), .Y(n43354) );
  INVX1 U45412 ( .A(n43357), .Y(n43355) );
  INVX1 U45413 ( .A(n43357), .Y(n43356) );
  INVX1 U45414 ( .A(n41786), .Y(n43357) );
  INVX1 U45415 ( .A(n37399), .Y(n43358) );
  INVX1 U45416 ( .A(n37399), .Y(n43359) );
  INVX1 U45417 ( .A(n37399), .Y(n43360) );
  INVX1 U45418 ( .A(n43364), .Y(n43361) );
  INVX1 U45419 ( .A(n43364), .Y(n43362) );
  INVX1 U45420 ( .A(n43364), .Y(n43363) );
  INVX1 U45421 ( .A(n42164), .Y(n43364) );
  INVX1 U45422 ( .A(n43368), .Y(n43365) );
  INVX1 U45423 ( .A(n43368), .Y(n43366) );
  INVX1 U45424 ( .A(n43368), .Y(n43367) );
  INVX1 U45425 ( .A(n42159), .Y(n43368) );
  INVX1 U45426 ( .A(n38764), .Y(n43369) );
  INVX1 U45427 ( .A(n38764), .Y(n43370) );
  INVX1 U45428 ( .A(n38764), .Y(n43371) );
  INVX1 U45429 ( .A(n47637), .Y(n43372) );
  INVX1 U45430 ( .A(n47637), .Y(n43373) );
  INVX1 U45431 ( .A(n43376), .Y(n43374) );
  INVX1 U45432 ( .A(n43376), .Y(n43375) );
  INVX1 U45433 ( .A(n57902), .Y(n43376) );
  INVX1 U45434 ( .A(n57902), .Y(n43377) );
  INVX1 U45435 ( .A(n57397), .Y(n43378) );
  INVX1 U45436 ( .A(n57397), .Y(n43379) );
  INVX1 U45437 ( .A(n57397), .Y(n43380) );
  INVX1 U45438 ( .A(n57899), .Y(n43381) );
  INVX1 U45439 ( .A(n57899), .Y(n43382) );
  INVX1 U45440 ( .A(n37469), .Y(n43383) );
  INVX1 U45441 ( .A(n37469), .Y(n43384) );
  INVX1 U45442 ( .A(n37469), .Y(n43385) );
  INVX1 U45443 ( .A(n42586), .Y(n43386) );
  INVX1 U45444 ( .A(n42586), .Y(n43387) );
  INVX1 U45445 ( .A(n42586), .Y(n43388) );
  INVX1 U45446 ( .A(n37473), .Y(n43389) );
  INVX1 U45447 ( .A(n37473), .Y(n43390) );
  INVX1 U45448 ( .A(n37473), .Y(n43391) );
  INVX1 U45449 ( .A(n42217), .Y(n43392) );
  INVX1 U45450 ( .A(n42217), .Y(n43393) );
  INVX1 U45451 ( .A(n42217), .Y(n43394) );
  INVX1 U45452 ( .A(n42307), .Y(n43395) );
  INVX1 U45453 ( .A(n42307), .Y(n43396) );
  INVX1 U45454 ( .A(n42307), .Y(n43397) );
  INVX1 U45455 ( .A(n36766), .Y(n43398) );
  INVX1 U45456 ( .A(n36766), .Y(n43399) );
  INVX1 U45457 ( .A(n36766), .Y(n43400) );
  INVX1 U45458 ( .A(n43403), .Y(n43401) );
  INVX1 U45459 ( .A(n43403), .Y(n43402) );
  INVX1 U45460 ( .A(n42138), .Y(n43403) );
  INVX1 U45461 ( .A(n42262), .Y(n43404) );
  INVX1 U45462 ( .A(n42262), .Y(n43405) );
  INVX1 U45463 ( .A(n8801), .Y(n43406) );
  INVX1 U45464 ( .A(n8801), .Y(n43407) );
  INVX1 U45465 ( .A(n43411), .Y(n43408) );
  INVX1 U45466 ( .A(n43411), .Y(n43409) );
  INVX1 U45467 ( .A(n43411), .Y(n43410) );
  INVX1 U45468 ( .A(n58556), .Y(n43411) );
  INVX1 U45469 ( .A(n58556), .Y(n43412) );
  INVX1 U45470 ( .A(n42451), .Y(n43413) );
  INVX1 U45471 ( .A(n43415), .Y(n43414) );
  INVX1 U45472 ( .A(n43413), .Y(n43415) );
  INVX1 U45473 ( .A(n42435), .Y(n43416) );
  INVX1 U45474 ( .A(n43419), .Y(n43417) );
  INVX1 U45475 ( .A(n43419), .Y(n43418) );
  INVX1 U45476 ( .A(n43416), .Y(n43419) );
  INVX1 U45477 ( .A(n43416), .Y(n43420) );
  INVX1 U45478 ( .A(n42316), .Y(n43421) );
  INVX1 U45479 ( .A(n42316), .Y(n43422) );
  INVX1 U45480 ( .A(n42316), .Y(n43423) );
  INVX1 U45481 ( .A(n43421), .Y(n43424) );
  INVX1 U45482 ( .A(n43422), .Y(n43425) );
  INVX1 U45483 ( .A(n43431), .Y(n43426) );
  INVX1 U45484 ( .A(n43430), .Y(n43427) );
  INVX1 U45485 ( .A(n43430), .Y(n43428) );
  INVX1 U45486 ( .A(n43430), .Y(n43429) );
  INVX1 U45487 ( .A(n58801), .Y(n43430) );
  INVX1 U45488 ( .A(n58801), .Y(n43431) );
  INVX1 U45489 ( .A(n58802), .Y(n43432) );
  INVX1 U45490 ( .A(n58802), .Y(n43433) );
  INVX1 U45491 ( .A(n58802), .Y(n43434) );
  INVX1 U45492 ( .A(n43440), .Y(n43435) );
  INVX1 U45493 ( .A(n43440), .Y(n43436) );
  INVX1 U45494 ( .A(n43434), .Y(n43437) );
  INVX1 U45495 ( .A(n43440), .Y(n43438) );
  INVX1 U45496 ( .A(n43440), .Y(n43439) );
  INVX1 U45497 ( .A(n58802), .Y(n43440) );
  INVX1 U45498 ( .A(n58759), .Y(n43441) );
  INVX1 U45499 ( .A(n58759), .Y(n43442) );
  INVX1 U45500 ( .A(n73383), .Y(n43443) );
  INVX1 U45501 ( .A(n73383), .Y(n43444) );
  INVX1 U45502 ( .A(n58977), .Y(n43445) );
  INVX1 U45503 ( .A(n58977), .Y(n43446) );
  INVX1 U45504 ( .A(n59112), .Y(n43447) );
  INVX1 U45505 ( .A(n42980), .Y(n43448) );
  INVX1 U45506 ( .A(n42981), .Y(n43449) );
  INVX1 U45507 ( .A(n59145), .Y(n43450) );
  INVX1 U45508 ( .A(n62904), .Y(n43451) );
  INVX1 U45509 ( .A(n62904), .Y(n43452) );
  INVX1 U45510 ( .A(n62904), .Y(n43453) );
  INVX1 U45511 ( .A(n38271), .Y(n43454) );
  INVX1 U45512 ( .A(n38271), .Y(n43455) );
  INVX1 U45513 ( .A(n39626), .Y(n43456) );
  INVX1 U45514 ( .A(n43459), .Y(n43457) );
  INVX1 U45515 ( .A(n39626), .Y(n43458) );
  INVX1 U45516 ( .A(n62659), .Y(n43459) );
  INVX1 U45517 ( .A(n62659), .Y(n43460) );
  INVX1 U45518 ( .A(n40228), .Y(n43461) );
  INVX1 U45519 ( .A(n63824), .Y(n43462) );
  INVX1 U45520 ( .A(n40524), .Y(n43463) );
  INVX1 U45521 ( .A(n43469), .Y(n43464) );
  INVX1 U45522 ( .A(n43468), .Y(n43465) );
  INVX1 U45523 ( .A(n43468), .Y(n43466) );
  INVX1 U45524 ( .A(n43468), .Y(n43467) );
  INVX1 U45525 ( .A(n62923), .Y(n43468) );
  INVX1 U45526 ( .A(n62923), .Y(n43469) );
  INVX1 U45527 ( .A(n62923), .Y(n43470) );
  INVX1 U45528 ( .A(n43473), .Y(n43471) );
  INVX1 U45529 ( .A(n43473), .Y(n43472) );
  INVX1 U45530 ( .A(n63222), .Y(n43473) );
  INVX1 U45531 ( .A(n38592), .Y(n43474) );
  INVX1 U45532 ( .A(n38644), .Y(n43475) );
  INVX1 U45533 ( .A(n63209), .Y(n43476) );
  INVX1 U45534 ( .A(n43480), .Y(n43477) );
  INVX1 U45535 ( .A(n43480), .Y(n43478) );
  INVX1 U45536 ( .A(n43480), .Y(n43479) );
  INVX1 U45537 ( .A(n70051), .Y(n43480) );
  INVX1 U45538 ( .A(n70051), .Y(n43481) );
  INVX1 U45539 ( .A(n43485), .Y(n43482) );
  INVX1 U45540 ( .A(n43485), .Y(n43483) );
  INVX1 U45541 ( .A(n43485), .Y(n43484) );
  INVX1 U45542 ( .A(n70371), .Y(n43485) );
  INVX1 U45543 ( .A(n43489), .Y(n43486) );
  INVX1 U45544 ( .A(n43489), .Y(n43487) );
  INVX1 U45545 ( .A(n43490), .Y(n43488) );
  INVX1 U45546 ( .A(n70671), .Y(n43489) );
  INVX1 U45547 ( .A(n70671), .Y(n43490) );
  INVX1 U45548 ( .A(n43495), .Y(n43491) );
  INVX1 U45549 ( .A(n43494), .Y(n43492) );
  INVX1 U45550 ( .A(n43494), .Y(n43493) );
  INVX1 U45551 ( .A(n39959), .Y(n43494) );
  INVX1 U45552 ( .A(n39959), .Y(n43495) );
  INVX1 U45553 ( .A(n40500), .Y(n43496) );
  INVX1 U45554 ( .A(n43499), .Y(n43497) );
  INVX1 U45555 ( .A(n71297), .Y(n43498) );
  INVX1 U45556 ( .A(n71297), .Y(n43499) );
  INVX1 U45557 ( .A(n43504), .Y(n43500) );
  INVX1 U45558 ( .A(n43504), .Y(n43501) );
  INVX1 U45559 ( .A(n43503), .Y(n43502) );
  INVX1 U45560 ( .A(n71546), .Y(n43503) );
  INVX1 U45561 ( .A(n71546), .Y(n43504) );
  INVX1 U45562 ( .A(n43511), .Y(n43505) );
  INVX1 U45563 ( .A(n43511), .Y(n43506) );
  INVX1 U45564 ( .A(n43510), .Y(n43507) );
  INVX1 U45565 ( .A(n43510), .Y(n43508) );
  INVX1 U45566 ( .A(n43510), .Y(n43509) );
  INVX1 U45567 ( .A(n43516), .Y(n43510) );
  INVX1 U45568 ( .A(n43516), .Y(n43511) );
  INVX1 U45569 ( .A(n41417), .Y(n43512) );
  INVX1 U45570 ( .A(n43515), .Y(n43513) );
  INVX1 U45571 ( .A(n43515), .Y(n43514) );
  INVX1 U45572 ( .A(n71734), .Y(n43515) );
  INVX1 U45573 ( .A(n71734), .Y(n43516) );
  INVX1 U45574 ( .A(n43519), .Y(n43517) );
  INVX1 U45575 ( .A(n43519), .Y(n43518) );
  INVX1 U45576 ( .A(n39868), .Y(n43519) );
  INVX1 U45577 ( .A(n39961), .Y(n43520) );
  INVX1 U45578 ( .A(n43526), .Y(n43521) );
  INVX1 U45579 ( .A(n43525), .Y(n43522) );
  INVX1 U45580 ( .A(n43525), .Y(n43523) );
  INVX1 U45581 ( .A(n43525), .Y(n43524) );
  INVX1 U45582 ( .A(n43533), .Y(n43525) );
  INVX1 U45583 ( .A(n43534), .Y(n43526) );
  INVX1 U45584 ( .A(n40345), .Y(n43527) );
  INVX1 U45585 ( .A(n39838), .Y(n43528) );
  INVX1 U45586 ( .A(n39838), .Y(n43529) );
  INVX1 U45587 ( .A(n39838), .Y(n43530) );
  INVX1 U45588 ( .A(n43534), .Y(n43531) );
  INVX1 U45589 ( .A(n43533), .Y(n43532) );
  INVX1 U45590 ( .A(n72139), .Y(n43533) );
  INVX1 U45591 ( .A(n72139), .Y(n43534) );
  INVX1 U45592 ( .A(n43539), .Y(n43535) );
  INVX1 U45593 ( .A(n72145), .Y(n43536) );
  INVX1 U45594 ( .A(n72145), .Y(n43537) );
  INVX1 U45595 ( .A(n43543), .Y(n43538) );
  INVX1 U45596 ( .A(n43543), .Y(n43539) );
  INVX1 U45597 ( .A(n43543), .Y(n43540) );
  INVX1 U45598 ( .A(n41317), .Y(n43541) );
  INVX1 U45599 ( .A(n43543), .Y(n43542) );
  INVX1 U45600 ( .A(n72145), .Y(n43543) );
  INVX1 U45601 ( .A(n43550), .Y(n43544) );
  INVX1 U45602 ( .A(n43548), .Y(n43545) );
  INVX1 U45603 ( .A(n72153), .Y(n43546) );
  INVX1 U45604 ( .A(n43554), .Y(n43547) );
  INVX1 U45605 ( .A(n43555), .Y(n43548) );
  INVX1 U45606 ( .A(n43555), .Y(n43549) );
  INVX1 U45607 ( .A(n43555), .Y(n43550) );
  INVX1 U45608 ( .A(n43554), .Y(n43551) );
  INVX1 U45609 ( .A(n43554), .Y(n43552) );
  INVX1 U45610 ( .A(n43554), .Y(n43553) );
  INVX1 U45611 ( .A(n72153), .Y(n43554) );
  INVX1 U45612 ( .A(n72153), .Y(n43555) );
  INVX1 U45613 ( .A(n36760), .Y(n43556) );
  INVX1 U45614 ( .A(n36760), .Y(n43557) );
  INVX1 U45615 ( .A(n36760), .Y(n43558) );
  INVX1 U45616 ( .A(n43561), .Y(n43559) );
  INVX1 U45617 ( .A(n36760), .Y(n43560) );
  INVX1 U45618 ( .A(n43556), .Y(n43561) );
  INVX1 U45619 ( .A(n43556), .Y(n43562) );
  INVX1 U45620 ( .A(n43557), .Y(n43563) );
  INVX1 U45621 ( .A(n43557), .Y(n43564) );
  INVX1 U45622 ( .A(n43557), .Y(n43565) );
  INVX1 U45623 ( .A(n43558), .Y(n43566) );
  INVX1 U45624 ( .A(n72168), .Y(n43567) );
  INVX1 U45625 ( .A(n72168), .Y(n43568) );
  INVX1 U45626 ( .A(n72168), .Y(n43569) );
  INVX1 U45627 ( .A(n42191), .Y(n43570) );
  INVX1 U45628 ( .A(n42191), .Y(n43571) );
  INVX1 U45629 ( .A(n42191), .Y(n43572) );
  INVX1 U45630 ( .A(n43575), .Y(n43573) );
  INVX1 U45631 ( .A(n43575), .Y(n43574) );
  INVX1 U45632 ( .A(n43570), .Y(n43575) );
  INVX1 U45633 ( .A(n43571), .Y(n43576) );
  INVX1 U45634 ( .A(n43571), .Y(n43577) );
  INVX1 U45635 ( .A(n43572), .Y(n43578) );
  INVX1 U45636 ( .A(n43572), .Y(n43579) );
  INVX1 U45637 ( .A(n43572), .Y(n43580) );
  INVX1 U45638 ( .A(n43584), .Y(n43581) );
  INVX1 U45639 ( .A(n43584), .Y(n43582) );
  INVX1 U45640 ( .A(n43584), .Y(n43583) );
  INVX1 U45641 ( .A(n43591), .Y(n43584) );
  INVX1 U45642 ( .A(n43590), .Y(n43585) );
  INVX1 U45643 ( .A(n43590), .Y(n43586) );
  INVX1 U45644 ( .A(n43590), .Y(n43587) );
  INVX1 U45645 ( .A(n43590), .Y(n43588) );
  INVX1 U45646 ( .A(n43590), .Y(n43589) );
  INVX1 U45647 ( .A(n72182), .Y(n43590) );
  INVX1 U45648 ( .A(n72182), .Y(n43591) );
  INVX1 U45649 ( .A(n42993), .Y(n43592) );
  INVX1 U45650 ( .A(n42992), .Y(n43593) );
  INVX1 U45651 ( .A(n42994), .Y(n43594) );
  INVX1 U45652 ( .A(n42190), .Y(n43595) );
  INVX1 U45653 ( .A(n42190), .Y(n43596) );
  INVX1 U45654 ( .A(n43599), .Y(n43597) );
  INVX1 U45655 ( .A(n42190), .Y(n43598) );
  INVX1 U45656 ( .A(n43595), .Y(n43599) );
  INVX1 U45657 ( .A(n43596), .Y(n43600) );
  INVX1 U45658 ( .A(n43596), .Y(n43601) );
  INVX1 U45659 ( .A(n43596), .Y(n43602) );
  INVX1 U45660 ( .A(n43606), .Y(n43603) );
  INVX1 U45661 ( .A(n43606), .Y(n43604) );
  INVX1 U45662 ( .A(n43606), .Y(n43605) );
  INVX1 U45663 ( .A(n72336), .Y(n43606) );
  INVX1 U45664 ( .A(n43611), .Y(n43607) );
  INVX1 U45665 ( .A(n43610), .Y(n43608) );
  INVX1 U45666 ( .A(n43610), .Y(n43609) );
  INVX1 U45667 ( .A(n72348), .Y(n43610) );
  INVX1 U45668 ( .A(n72348), .Y(n43611) );
  INVX1 U45669 ( .A(n37415), .Y(n43612) );
  INVX1 U45670 ( .A(n37415), .Y(n43613) );
  INVX1 U45671 ( .A(n37415), .Y(n43614) );
  INVX1 U45672 ( .A(n72536), .Y(n43615) );
  INVX1 U45673 ( .A(n72536), .Y(n43616) );
  INVX1 U45674 ( .A(n42996), .Y(n43617) );
  INVX1 U45675 ( .A(n42997), .Y(n43618) );
  INVX1 U45676 ( .A(n43622), .Y(n43619) );
  INVX1 U45677 ( .A(n43622), .Y(n43620) );
  INVX1 U45678 ( .A(n43622), .Y(n43621) );
  INVX1 U45679 ( .A(n43629), .Y(n43622) );
  INVX1 U45680 ( .A(n43630), .Y(n43623) );
  INVX1 U45681 ( .A(n43630), .Y(n43624) );
  INVX1 U45682 ( .A(n43630), .Y(n43625) );
  INVX1 U45683 ( .A(n43630), .Y(n43626) );
  INVX1 U45684 ( .A(n43629), .Y(n43627) );
  INVX1 U45685 ( .A(n43629), .Y(n43628) );
  INVX1 U45686 ( .A(n72558), .Y(n43629) );
  INVX1 U45687 ( .A(n72558), .Y(n43630) );
  INVX1 U45688 ( .A(n43634), .Y(n43631) );
  INVX1 U45689 ( .A(n43634), .Y(n43632) );
  INVX1 U45690 ( .A(n43634), .Y(n43633) );
  INVX1 U45691 ( .A(n43641), .Y(n43634) );
  INVX1 U45692 ( .A(n43640), .Y(n43635) );
  INVX1 U45693 ( .A(n43640), .Y(n43636) );
  INVX1 U45694 ( .A(n40276), .Y(n43637) );
  INVX1 U45695 ( .A(n43641), .Y(n43638) );
  INVX1 U45696 ( .A(n43640), .Y(n43639) );
  INVX1 U45697 ( .A(n72591), .Y(n43640) );
  INVX1 U45698 ( .A(n72591), .Y(n43641) );
  INVX1 U45699 ( .A(n43645), .Y(n43642) );
  INVX1 U45700 ( .A(n43645), .Y(n43643) );
  INVX1 U45701 ( .A(n43645), .Y(n43644) );
  INVX1 U45702 ( .A(n43652), .Y(n43645) );
  INVX1 U45703 ( .A(n43651), .Y(n43646) );
  INVX1 U45704 ( .A(n43651), .Y(n43647) );
  INVX1 U45705 ( .A(n43651), .Y(n43648) );
  INVX1 U45706 ( .A(n43651), .Y(n43649) );
  INVX1 U45707 ( .A(n43644), .Y(n43650) );
  INVX1 U45708 ( .A(n72613), .Y(n43651) );
  INVX1 U45709 ( .A(n72613), .Y(n43652) );
  INVX1 U45710 ( .A(n43660), .Y(n43653) );
  INVX1 U45711 ( .A(n72620), .Y(n43654) );
  INVX1 U45712 ( .A(n43660), .Y(n43655) );
  INVX1 U45713 ( .A(n43663), .Y(n43656) );
  INVX1 U45714 ( .A(n43663), .Y(n43657) );
  INVX1 U45715 ( .A(n43663), .Y(n43658) );
  INVX1 U45716 ( .A(n43662), .Y(n43659) );
  INVX1 U45717 ( .A(n43662), .Y(n43660) );
  INVX1 U45718 ( .A(n43663), .Y(n43661) );
  INVX1 U45719 ( .A(n72620), .Y(n43662) );
  INVX1 U45720 ( .A(n72620), .Y(n43663) );
  INVX1 U45721 ( .A(n43671), .Y(n43664) );
  INVX1 U45722 ( .A(n43670), .Y(n43665) );
  INVX1 U45723 ( .A(n72626), .Y(n43666) );
  INVX1 U45724 ( .A(n43669), .Y(n43667) );
  INVX1 U45725 ( .A(n43675), .Y(n43668) );
  INVX1 U45726 ( .A(n43675), .Y(n43669) );
  INVX1 U45727 ( .A(n43674), .Y(n43670) );
  INVX1 U45728 ( .A(n43674), .Y(n43671) );
  INVX1 U45729 ( .A(n43674), .Y(n43672) );
  INVX1 U45730 ( .A(n43667), .Y(n43673) );
  INVX1 U45731 ( .A(n72626), .Y(n43674) );
  INVX1 U45732 ( .A(n72626), .Y(n43675) );
  INVX1 U45733 ( .A(n43681), .Y(n43676) );
  INVX1 U45734 ( .A(n43681), .Y(n43677) );
  INVX1 U45735 ( .A(n43680), .Y(n43678) );
  INVX1 U45736 ( .A(n43680), .Y(n43679) );
  INVX1 U45737 ( .A(n43690), .Y(n43680) );
  INVX1 U45738 ( .A(n43690), .Y(n43681) );
  INVX1 U45739 ( .A(n43689), .Y(n43682) );
  INVX1 U45740 ( .A(n43689), .Y(n43683) );
  INVX1 U45741 ( .A(n43689), .Y(n43684) );
  INVX1 U45742 ( .A(n41374), .Y(n43685) );
  INVX1 U45743 ( .A(n43689), .Y(n43686) );
  INVX1 U45744 ( .A(n37975), .Y(n43687) );
  INVX1 U45745 ( .A(n43689), .Y(n43688) );
  INVX1 U45746 ( .A(n72675), .Y(n43689) );
  INVX1 U45747 ( .A(n72675), .Y(n43690) );
  INVX1 U45748 ( .A(n43702), .Y(n43691) );
  INVX1 U45749 ( .A(n43695), .Y(n43692) );
  INVX1 U45750 ( .A(n43695), .Y(n43693) );
  INVX1 U45751 ( .A(n43695), .Y(n43694) );
  INVX1 U45752 ( .A(n43704), .Y(n43695) );
  INVX1 U45753 ( .A(n41454), .Y(n43696) );
  INVX1 U45754 ( .A(n41454), .Y(n43697) );
  INVX1 U45755 ( .A(n43691), .Y(n43698) );
  INVX1 U45756 ( .A(n43703), .Y(n43699) );
  INVX1 U45757 ( .A(n43704), .Y(n43700) );
  INVX1 U45758 ( .A(n43704), .Y(n43701) );
  INVX1 U45759 ( .A(n43703), .Y(n43702) );
  INVX1 U45760 ( .A(n72698), .Y(n43703) );
  INVX1 U45761 ( .A(n72698), .Y(n43704) );
  INVX1 U45762 ( .A(n43710), .Y(n43705) );
  INVX1 U45763 ( .A(n72708), .Y(n43706) );
  INVX1 U45764 ( .A(n43713), .Y(n43707) );
  INVX1 U45765 ( .A(n40456), .Y(n43708) );
  INVX1 U45766 ( .A(n40456), .Y(n43709) );
  INVX1 U45767 ( .A(n43717), .Y(n43710) );
  INVX1 U45768 ( .A(n43717), .Y(n43711) );
  INVX1 U45769 ( .A(n43716), .Y(n43712) );
  INVX1 U45770 ( .A(n43716), .Y(n43713) );
  INVX1 U45771 ( .A(n43716), .Y(n43714) );
  INVX1 U45772 ( .A(n43717), .Y(n43715) );
  INVX1 U45773 ( .A(n72708), .Y(n43716) );
  INVX1 U45774 ( .A(n72708), .Y(n43717) );
  INVX1 U45775 ( .A(n43721), .Y(n43718) );
  INVX1 U45776 ( .A(n43721), .Y(n43719) );
  INVX1 U45777 ( .A(n43721), .Y(n43720) );
  INVX1 U45778 ( .A(n72728), .Y(n43721) );
  INVX1 U45779 ( .A(n72741), .Y(n43722) );
  INVX1 U45780 ( .A(n72741), .Y(n43723) );
  INVX1 U45781 ( .A(n43728), .Y(n43724) );
  INVX1 U45782 ( .A(n43728), .Y(n43725) );
  INVX1 U45783 ( .A(n43725), .Y(n43726) );
  INVX1 U45784 ( .A(n38110), .Y(n43727) );
  INVX1 U45785 ( .A(n38111), .Y(n43728) );
  INVX1 U45786 ( .A(n43734), .Y(n43729) );
  INVX1 U45787 ( .A(n43733), .Y(n43730) );
  INVX1 U45788 ( .A(n43733), .Y(n43731) );
  INVX1 U45789 ( .A(n43733), .Y(n43732) );
  INVX1 U45790 ( .A(n72759), .Y(n43733) );
  INVX1 U45791 ( .A(n72759), .Y(n43734) );
  INVX1 U45792 ( .A(n43740), .Y(n43735) );
  INVX1 U45793 ( .A(n43739), .Y(n43736) );
  INVX1 U45794 ( .A(n43739), .Y(n43737) );
  INVX1 U45795 ( .A(n43739), .Y(n43738) );
  INVX1 U45796 ( .A(n72760), .Y(n43739) );
  INVX1 U45797 ( .A(n72760), .Y(n43740) );
  INVX1 U45798 ( .A(n43746), .Y(n43741) );
  INVX1 U45799 ( .A(n43745), .Y(n43742) );
  INVX1 U45800 ( .A(n43745), .Y(n43743) );
  INVX1 U45801 ( .A(n43745), .Y(n43744) );
  INVX1 U45802 ( .A(n72765), .Y(n43745) );
  INVX1 U45803 ( .A(n72765), .Y(n43746) );
  INVX1 U45804 ( .A(n72765), .Y(n43747) );
  INVX1 U45805 ( .A(n72766), .Y(n43748) );
  INVX1 U45806 ( .A(n72766), .Y(n43749) );
  INVX1 U45807 ( .A(n43755), .Y(n43750) );
  INVX1 U45808 ( .A(n43754), .Y(n43751) );
  INVX1 U45809 ( .A(n43754), .Y(n43752) );
  INVX1 U45810 ( .A(n43754), .Y(n43753) );
  INVX1 U45811 ( .A(n72779), .Y(n43754) );
  INVX1 U45812 ( .A(n72779), .Y(n43755) );
  INVX1 U45813 ( .A(n72779), .Y(n43756) );
  INVX1 U45814 ( .A(n43761), .Y(n43757) );
  INVX1 U45815 ( .A(n43760), .Y(n43758) );
  INVX1 U45816 ( .A(n43760), .Y(n43759) );
  INVX1 U45817 ( .A(n72780), .Y(n43760) );
  INVX1 U45818 ( .A(n72780), .Y(n43761) );
  INVX1 U45819 ( .A(n72783), .Y(n43762) );
  INVX1 U45820 ( .A(n43768), .Y(n43763) );
  INVX1 U45821 ( .A(n43767), .Y(n43764) );
  INVX1 U45822 ( .A(n43767), .Y(n43765) );
  INVX1 U45823 ( .A(n43767), .Y(n43766) );
  INVX1 U45824 ( .A(n72786), .Y(n43767) );
  INVX1 U45825 ( .A(n72786), .Y(n43768) );
  INVX1 U45826 ( .A(n72786), .Y(n43769) );
  INVX1 U45827 ( .A(n72787), .Y(n43770) );
  INVX1 U45828 ( .A(n72787), .Y(n43771) );
  INVX1 U45829 ( .A(n42824), .Y(n43772) );
  INVX1 U45830 ( .A(n42824), .Y(n43773) );
  INVX1 U45831 ( .A(n43777), .Y(n43774) );
  INVX1 U45832 ( .A(n43777), .Y(n43775) );
  INVX1 U45833 ( .A(n43777), .Y(n43776) );
  INVX1 U45834 ( .A(n72803), .Y(n43777) );
  INVX1 U45835 ( .A(n72803), .Y(n43778) );
  INVX1 U45836 ( .A(n43785), .Y(n43779) );
  INVX1 U45837 ( .A(n43784), .Y(n43780) );
  INVX1 U45838 ( .A(n43784), .Y(n43781) );
  INVX1 U45839 ( .A(n43783), .Y(n43782) );
  INVX1 U45840 ( .A(n72806), .Y(n43783) );
  INVX1 U45841 ( .A(n72806), .Y(n43784) );
  INVX1 U45842 ( .A(n72806), .Y(n43785) );
  INVX1 U45843 ( .A(n43790), .Y(n43786) );
  INVX1 U45844 ( .A(n43789), .Y(n43787) );
  INVX1 U45845 ( .A(n43789), .Y(n43788) );
  INVX1 U45846 ( .A(n72807), .Y(n43789) );
  INVX1 U45847 ( .A(n72807), .Y(n43790) );
  INVX1 U45848 ( .A(n43794), .Y(n43791) );
  INVX1 U45849 ( .A(n43793), .Y(n43792) );
  INVX1 U45850 ( .A(n72810), .Y(n43793) );
  INVX1 U45851 ( .A(n72810), .Y(n43794) );
  INVX1 U45852 ( .A(n43797), .Y(n43795) );
  INVX1 U45853 ( .A(n43797), .Y(n43796) );
  INVX1 U45854 ( .A(n72811), .Y(n43797) );
  INVX1 U45855 ( .A(n43801), .Y(n43798) );
  INVX1 U45856 ( .A(n43801), .Y(n43799) );
  INVX1 U45857 ( .A(n43801), .Y(n43800) );
  INVX1 U45858 ( .A(n72815), .Y(n43801) );
  INVX1 U45859 ( .A(n43808), .Y(n43802) );
  INVX1 U45860 ( .A(n43806), .Y(n43803) );
  INVX1 U45861 ( .A(n43806), .Y(n43804) );
  INVX1 U45862 ( .A(n43806), .Y(n43805) );
  INVX1 U45863 ( .A(n72819), .Y(n43806) );
  INVX1 U45864 ( .A(n72819), .Y(n43807) );
  INVX1 U45865 ( .A(n72819), .Y(n43808) );
  INVX1 U45866 ( .A(n43813), .Y(n43809) );
  INVX1 U45867 ( .A(n40543), .Y(n43810) );
  INVX1 U45868 ( .A(n40543), .Y(n43811) );
  INVX1 U45869 ( .A(n43813), .Y(n43812) );
  INVX1 U45870 ( .A(n43810), .Y(n43813) );
  INVX1 U45871 ( .A(n43818), .Y(n43814) );
  INVX1 U45872 ( .A(n43817), .Y(n43815) );
  INVX1 U45873 ( .A(n43817), .Y(n43816) );
  INVX1 U45874 ( .A(n38106), .Y(n43817) );
  INVX1 U45875 ( .A(n38105), .Y(n43818) );
  INVX1 U45876 ( .A(n43822), .Y(n43819) );
  INVX1 U45877 ( .A(n43822), .Y(n43820) );
  INVX1 U45878 ( .A(n43822), .Y(n43821) );
  INVX1 U45879 ( .A(n72825), .Y(n43822) );
  INVX1 U45880 ( .A(n37444), .Y(n43823) );
  INVX1 U45881 ( .A(n37444), .Y(n43824) );
  INVX1 U45882 ( .A(n37444), .Y(n43825) );
  INVX1 U45883 ( .A(n43828), .Y(n43826) );
  INVX1 U45884 ( .A(n43828), .Y(n43827) );
  INVX1 U45885 ( .A(n42140), .Y(n43828) );
  INVX1 U45886 ( .A(n42132), .Y(n43829) );
  INVX1 U45887 ( .A(n42132), .Y(n43830) );
  INVX1 U45888 ( .A(n42132), .Y(n43831) );
  INVX1 U45889 ( .A(n43834), .Y(n43832) );
  INVX1 U45890 ( .A(n43834), .Y(n43833) );
  INVX1 U45891 ( .A(n42212), .Y(n43834) );
  INVX1 U45892 ( .A(n43837), .Y(n43835) );
  INVX1 U45893 ( .A(n43837), .Y(n43836) );
  INVX1 U45894 ( .A(n42304), .Y(n43837) );
  INVX1 U45895 ( .A(n42228), .Y(n43838) );
  INVX1 U45896 ( .A(n42228), .Y(n43839) );
  INVX1 U45897 ( .A(n43845), .Y(n43840) );
  INVX1 U45898 ( .A(n43844), .Y(n43841) );
  INVX1 U45899 ( .A(n43844), .Y(n43842) );
  INVX1 U45900 ( .A(n43844), .Y(n43843) );
  INVX1 U45901 ( .A(n43838), .Y(n43844) );
  INVX1 U45902 ( .A(n43838), .Y(n43845) );
  INVX1 U45903 ( .A(n43839), .Y(n43846) );
  INVX1 U45904 ( .A(n43839), .Y(n43847) );
  INVX1 U45905 ( .A(n42239), .Y(n43848) );
  INVX1 U45906 ( .A(n42239), .Y(n43849) );
  INVX1 U45907 ( .A(n42239), .Y(n43850) );
  INVX1 U45908 ( .A(n43854), .Y(n43851) );
  INVX1 U45909 ( .A(n43854), .Y(n43852) );
  INVX1 U45910 ( .A(n43854), .Y(n43853) );
  INVX1 U45911 ( .A(n43848), .Y(n43854) );
  INVX1 U45912 ( .A(n43849), .Y(n43855) );
  INVX1 U45913 ( .A(n43849), .Y(n43856) );
  INVX1 U45914 ( .A(n42241), .Y(n43857) );
  INVX1 U45915 ( .A(n42241), .Y(n43858) );
  INVX1 U45916 ( .A(n43864), .Y(n43859) );
  INVX1 U45917 ( .A(n43863), .Y(n43860) );
  INVX1 U45918 ( .A(n43863), .Y(n43861) );
  INVX1 U45919 ( .A(n43863), .Y(n43862) );
  INVX1 U45920 ( .A(n43857), .Y(n43863) );
  INVX1 U45921 ( .A(n43857), .Y(n43864) );
  INVX1 U45922 ( .A(n43858), .Y(n43865) );
  INVX1 U45923 ( .A(n43858), .Y(n43866) );
  INVX1 U45924 ( .A(n42243), .Y(n43867) );
  INVX1 U45925 ( .A(n42243), .Y(n43868) );
  INVX1 U45926 ( .A(n42243), .Y(n43869) );
  INVX1 U45927 ( .A(n43873), .Y(n43870) );
  INVX1 U45928 ( .A(n43873), .Y(n43871) );
  INVX1 U45929 ( .A(n43873), .Y(n43872) );
  INVX1 U45930 ( .A(n43867), .Y(n43873) );
  INVX1 U45931 ( .A(n43868), .Y(n43874) );
  INVX1 U45932 ( .A(n43868), .Y(n43875) );
  INVX1 U45933 ( .A(n43868), .Y(n43876) );
  INVX1 U45934 ( .A(n42246), .Y(n43877) );
  INVX1 U45935 ( .A(n42246), .Y(n43878) );
  INVX1 U45936 ( .A(n42246), .Y(n43879) );
  INVX1 U45937 ( .A(n43883), .Y(n43880) );
  INVX1 U45938 ( .A(n43883), .Y(n43881) );
  INVX1 U45939 ( .A(n43883), .Y(n43882) );
  INVX1 U45940 ( .A(n43877), .Y(n43883) );
  INVX1 U45941 ( .A(n43877), .Y(n43884) );
  INVX1 U45942 ( .A(n43878), .Y(n43885) );
  INVX1 U45943 ( .A(n43878), .Y(n43886) );
  INVX1 U45944 ( .A(n42249), .Y(n43887) );
  INVX1 U45945 ( .A(n42249), .Y(n43888) );
  INVX1 U45946 ( .A(n42249), .Y(n43889) );
  INVX1 U45947 ( .A(n43893), .Y(n43890) );
  INVX1 U45948 ( .A(n43893), .Y(n43891) );
  INVX1 U45949 ( .A(n43893), .Y(n43892) );
  INVX1 U45950 ( .A(n43887), .Y(n43893) );
  INVX1 U45951 ( .A(n43887), .Y(n43894) );
  INVX1 U45952 ( .A(n43888), .Y(n43895) );
  INVX1 U45953 ( .A(n43902), .Y(n43896) );
  INVX1 U45954 ( .A(n43900), .Y(n43897) );
  INVX1 U45955 ( .A(n43900), .Y(n43898) );
  INVX1 U45956 ( .A(n43900), .Y(n43899) );
  INVX1 U45957 ( .A(n73216), .Y(n43900) );
  INVX1 U45958 ( .A(n73216), .Y(n43901) );
  INVX1 U45959 ( .A(n73216), .Y(n43902) );
  INVX1 U45960 ( .A(n43907), .Y(n43903) );
  INVX1 U45961 ( .A(n43907), .Y(n43904) );
  INVX1 U45962 ( .A(n43907), .Y(n43905) );
  INVX1 U45963 ( .A(n43907), .Y(n43906) );
  INVX1 U45964 ( .A(n73224), .Y(n43907) );
  INVX1 U45965 ( .A(n73224), .Y(n43908) );
  INVX1 U45966 ( .A(n43914), .Y(n43909) );
  INVX1 U45967 ( .A(n43913), .Y(n43910) );
  INVX1 U45968 ( .A(n43913), .Y(n43911) );
  INVX1 U45969 ( .A(n43913), .Y(n43912) );
  INVX1 U45970 ( .A(n73232), .Y(n43913) );
  INVX1 U45971 ( .A(n73232), .Y(n43914) );
  INVX1 U45972 ( .A(n73232), .Y(n43915) );
  INVX1 U45973 ( .A(n42255), .Y(n43916) );
  INVX1 U45974 ( .A(n42255), .Y(n43917) );
  INVX1 U45975 ( .A(n42255), .Y(n43918) );
  INVX1 U45976 ( .A(n43924), .Y(n43919) );
  INVX1 U45977 ( .A(n43922), .Y(n43920) );
  INVX1 U45978 ( .A(n43923), .Y(n43921) );
  INVX1 U45979 ( .A(n43916), .Y(n43922) );
  INVX1 U45980 ( .A(n43917), .Y(n43923) );
  INVX1 U45981 ( .A(n43917), .Y(n43924) );
  INVX1 U45982 ( .A(n42259), .Y(n43925) );
  INVX1 U45983 ( .A(n43932), .Y(n43926) );
  INVX1 U45984 ( .A(n42259), .Y(n43927) );
  INVX1 U45985 ( .A(n43932), .Y(n43928) );
  INVX1 U45986 ( .A(n43930), .Y(n43929) );
  INVX1 U45987 ( .A(n43925), .Y(n43930) );
  INVX1 U45988 ( .A(n43925), .Y(n43931) );
  INVX1 U45989 ( .A(n43925), .Y(n43932) );
  INVX1 U45990 ( .A(n43938), .Y(n43933) );
  INVX1 U45991 ( .A(n43937), .Y(n43934) );
  INVX1 U45992 ( .A(n43937), .Y(n43935) );
  INVX1 U45993 ( .A(n43937), .Y(n43936) );
  INVX1 U45994 ( .A(n73254), .Y(n43937) );
  INVX1 U45995 ( .A(n73254), .Y(n43938) );
  INVX1 U45996 ( .A(n73254), .Y(n43939) );
  INVX1 U45997 ( .A(n42265), .Y(n43940) );
  INVX1 U45998 ( .A(n42265), .Y(n43941) );
  INVX1 U45999 ( .A(n42265), .Y(n43942) );
  INVX1 U46000 ( .A(n43946), .Y(n43943) );
  INVX1 U46001 ( .A(n43946), .Y(n43944) );
  INVX1 U46002 ( .A(n43946), .Y(n43945) );
  INVX1 U46003 ( .A(n43940), .Y(n43946) );
  INVX1 U46004 ( .A(n43940), .Y(n43947) );
  INVX1 U46005 ( .A(n43941), .Y(n43948) );
  INVX1 U46006 ( .A(n43941), .Y(n43949) );
  INVX1 U46007 ( .A(n42240), .Y(n43950) );
  INVX1 U46008 ( .A(n42240), .Y(n43951) );
  INVX1 U46009 ( .A(n42240), .Y(n43952) );
  INVX1 U46010 ( .A(n43956), .Y(n43953) );
  INVX1 U46011 ( .A(n43956), .Y(n43954) );
  INVX1 U46012 ( .A(n43956), .Y(n43955) );
  INVX1 U46013 ( .A(n43950), .Y(n43956) );
  INVX1 U46014 ( .A(n43951), .Y(n43957) );
  INVX1 U46015 ( .A(n43951), .Y(n43958) );
  INVX1 U46016 ( .A(n43951), .Y(n43959) );
  INVX1 U46017 ( .A(n42242), .Y(n43960) );
  INVX1 U46018 ( .A(n42242), .Y(n43961) );
  INVX1 U46019 ( .A(n42242), .Y(n43962) );
  INVX1 U46020 ( .A(n43966), .Y(n43963) );
  INVX1 U46021 ( .A(n43966), .Y(n43964) );
  INVX1 U46022 ( .A(n43966), .Y(n43965) );
  INVX1 U46023 ( .A(n43960), .Y(n43966) );
  INVX1 U46024 ( .A(n43961), .Y(n43967) );
  INVX1 U46025 ( .A(n43961), .Y(n43968) );
  INVX1 U46026 ( .A(n43961), .Y(n43969) );
  INVX1 U46027 ( .A(n42269), .Y(n43970) );
  INVX1 U46028 ( .A(n42269), .Y(n43971) );
  INVX1 U46029 ( .A(n42269), .Y(n43972) );
  INVX1 U46030 ( .A(n43976), .Y(n43973) );
  INVX1 U46031 ( .A(n43976), .Y(n43974) );
  INVX1 U46032 ( .A(n43976), .Y(n43975) );
  INVX1 U46033 ( .A(n43970), .Y(n43976) );
  INVX1 U46034 ( .A(n43971), .Y(n43977) );
  INVX1 U46035 ( .A(n43971), .Y(n43978) );
  INVX1 U46036 ( .A(n43971), .Y(n43979) );
  INVX1 U46037 ( .A(n42272), .Y(n43980) );
  INVX1 U46038 ( .A(n42272), .Y(n43981) );
  INVX1 U46039 ( .A(n42272), .Y(n43982) );
  INVX1 U46040 ( .A(n43986), .Y(n43983) );
  INVX1 U46041 ( .A(n43986), .Y(n43984) );
  INVX1 U46042 ( .A(n43986), .Y(n43985) );
  INVX1 U46043 ( .A(n43980), .Y(n43986) );
  INVX1 U46044 ( .A(n43981), .Y(n43987) );
  INVX1 U46045 ( .A(n43981), .Y(n43988) );
  INVX1 U46046 ( .A(n43981), .Y(n43989) );
  INVX1 U46047 ( .A(n42275), .Y(n43990) );
  INVX1 U46048 ( .A(n42275), .Y(n43991) );
  INVX1 U46049 ( .A(n42275), .Y(n43992) );
  INVX1 U46050 ( .A(n43996), .Y(n43993) );
  INVX1 U46051 ( .A(n43995), .Y(n43994) );
  INVX1 U46052 ( .A(n43990), .Y(n43995) );
  INVX1 U46053 ( .A(n43990), .Y(n43996) );
  INVX1 U46054 ( .A(n42278), .Y(n43997) );
  INVX1 U46055 ( .A(n42278), .Y(n43998) );
  INVX1 U46056 ( .A(n42278), .Y(n43999) );
  INVX1 U46057 ( .A(n44003), .Y(n44000) );
  INVX1 U46058 ( .A(n44003), .Y(n44001) );
  INVX1 U46059 ( .A(n44003), .Y(n44002) );
  INVX1 U46060 ( .A(n43997), .Y(n44003) );
  INVX1 U46061 ( .A(n43997), .Y(n44004) );
  INVX1 U46062 ( .A(n43998), .Y(n44005) );
  INVX1 U46063 ( .A(n43998), .Y(n44006) );
  INVX1 U46064 ( .A(n44012), .Y(n44007) );
  INVX1 U46065 ( .A(n44011), .Y(n44008) );
  INVX1 U46066 ( .A(n44011), .Y(n44009) );
  INVX1 U46067 ( .A(n44011), .Y(n44010) );
  INVX1 U46068 ( .A(n73311), .Y(n44011) );
  INVX1 U46069 ( .A(n73311), .Y(n44012) );
  INVX1 U46070 ( .A(n73311), .Y(n44013) );
  INVX1 U46071 ( .A(n42281), .Y(n44014) );
  INVX1 U46072 ( .A(n42281), .Y(n44015) );
  INVX1 U46073 ( .A(n44022), .Y(n44016) );
  INVX1 U46074 ( .A(n42281), .Y(n44017) );
  INVX1 U46075 ( .A(n44021), .Y(n44018) );
  INVX1 U46076 ( .A(n44020), .Y(n44019) );
  INVX1 U46077 ( .A(n44014), .Y(n44020) );
  INVX1 U46078 ( .A(n44015), .Y(n44021) );
  INVX1 U46079 ( .A(n44015), .Y(n44022) );
  INVX1 U46080 ( .A(n42284), .Y(n44023) );
  INVX1 U46081 ( .A(n44029), .Y(n44024) );
  INVX1 U46082 ( .A(n42284), .Y(n44025) );
  INVX1 U46083 ( .A(n44029), .Y(n44026) );
  INVX1 U46084 ( .A(n42284), .Y(n44027) );
  INVX1 U46085 ( .A(n44023), .Y(n44028) );
  INVX1 U46086 ( .A(n44023), .Y(n44029) );
  INVX1 U46087 ( .A(n44032), .Y(n44030) );
  INVX1 U46088 ( .A(n44032), .Y(n44031) );
  INVX1 U46089 ( .A(n42141), .Y(n44032) );
  INVX1 U46090 ( .A(n42238), .Y(n44033) );
  INVX1 U46091 ( .A(n42238), .Y(n44034) );
  INVX1 U46092 ( .A(n42238), .Y(n44035) );
  INVX1 U46093 ( .A(n44039), .Y(n44036) );
  INVX1 U46094 ( .A(n44039), .Y(n44037) );
  INVX1 U46095 ( .A(n44039), .Y(n44038) );
  INVX1 U46096 ( .A(n44033), .Y(n44039) );
  INVX1 U46097 ( .A(n44033), .Y(n44040) );
  INVX1 U46098 ( .A(n44034), .Y(n44041) );
  INVX1 U46099 ( .A(n44044), .Y(n44042) );
  INVX1 U46100 ( .A(n44044), .Y(n44043) );
  INVX1 U46101 ( .A(n42139), .Y(n44044) );
  INVX1 U46102 ( .A(n42289), .Y(n44045) );
  INVX1 U46103 ( .A(n42289), .Y(n44046) );
  INVX1 U46104 ( .A(n44051), .Y(n44047) );
  INVX1 U46105 ( .A(n42289), .Y(n44048) );
  INVX1 U46106 ( .A(n44052), .Y(n44049) );
  INVX1 U46107 ( .A(n44053), .Y(n44050) );
  INVX1 U46108 ( .A(n44045), .Y(n44051) );
  INVX1 U46109 ( .A(n44046), .Y(n44052) );
  INVX1 U46110 ( .A(n44046), .Y(n44053) );
  INVX1 U46111 ( .A(n44059), .Y(n44054) );
  INVX1 U46112 ( .A(n44058), .Y(n44055) );
  INVX1 U46113 ( .A(n44058), .Y(n44056) );
  INVX1 U46114 ( .A(n44058), .Y(n44057) );
  INVX1 U46115 ( .A(n73379), .Y(n44058) );
  INVX1 U46116 ( .A(n73379), .Y(n44059) );
  INVX1 U46117 ( .A(n73379), .Y(n44060) );
  INVX1 U46118 ( .A(n73382), .Y(n44061) );
  INVX1 U46119 ( .A(n73382), .Y(n44062) );
  INVX1 U46120 ( .A(n73382), .Y(n44063) );
  INVX1 U46121 ( .A(n44068), .Y(n44064) );
  INVX1 U46122 ( .A(n44068), .Y(n44065) );
  INVX1 U46123 ( .A(n44068), .Y(n44066) );
  INVX1 U46124 ( .A(n44068), .Y(n44067) );
  INVX1 U46125 ( .A(n73382), .Y(n44068) );
  INVX1 U46126 ( .A(n39358), .Y(n44069) );
  INVX1 U46127 ( .A(n39358), .Y(n44070) );
  INVX1 U46128 ( .A(n44072), .Y(n44071) );
  INVX1 U46129 ( .A(n44069), .Y(n44072) );
  INVX1 U46130 ( .A(n58179), .Y(n44073) );
  INVX1 U46131 ( .A(n58179), .Y(n44074) );
  INVX1 U46132 ( .A(n44077), .Y(n44075) );
  INVX1 U46133 ( .A(n44077), .Y(n44076) );
  INVX1 U46134 ( .A(n42210), .Y(n44077) );
  INVX1 U46135 ( .A(n58275), .Y(n44078) );
  INVX1 U46136 ( .A(n58275), .Y(n44079) );
  INVX1 U46137 ( .A(n26912), .Y(n44080) );
  INVX1 U46138 ( .A(n26912), .Y(n44081) );
  INVX1 U46139 ( .A(n27964), .Y(n44082) );
  INVX1 U46140 ( .A(n27964), .Y(n44083) );
  INVX1 U46141 ( .A(n27964), .Y(n44084) );
  INVX1 U46142 ( .A(n57600), .Y(n44085) );
  INVX1 U46143 ( .A(n57600), .Y(n44086) );
  INVX1 U46144 ( .A(rst_i), .Y(n44087) );
  INVX1 U46145 ( .A(n44233), .Y(n44088) );
  INVX1 U46146 ( .A(n44246), .Y(n44089) );
  INVX1 U46147 ( .A(n44246), .Y(n44090) );
  INVX1 U46148 ( .A(n44246), .Y(n44091) );
  INVX1 U46149 ( .A(n44245), .Y(n44092) );
  INVX1 U46150 ( .A(n44245), .Y(n44093) );
  INVX1 U46151 ( .A(n44245), .Y(n44094) );
  INVX1 U46152 ( .A(n44244), .Y(n44095) );
  INVX1 U46153 ( .A(n44244), .Y(n44096) );
  INVX1 U46154 ( .A(n44244), .Y(n44097) );
  INVX1 U46155 ( .A(n44243), .Y(n44098) );
  INVX1 U46156 ( .A(n44243), .Y(n44099) );
  INVX1 U46157 ( .A(n44243), .Y(n44100) );
  INVX1 U46158 ( .A(n44242), .Y(n44101) );
  INVX1 U46159 ( .A(n44242), .Y(n44102) );
  INVX1 U46160 ( .A(n44242), .Y(n44103) );
  INVX1 U46161 ( .A(n44241), .Y(n44104) );
  INVX1 U46162 ( .A(n44241), .Y(n44105) );
  INVX1 U46163 ( .A(n44241), .Y(n44106) );
  INVX1 U46164 ( .A(n44240), .Y(n44107) );
  INVX1 U46165 ( .A(n44240), .Y(n44108) );
  INVX1 U46166 ( .A(n44240), .Y(n44109) );
  INVX1 U46167 ( .A(n44239), .Y(n44110) );
  INVX1 U46168 ( .A(n44239), .Y(n44111) );
  INVX1 U46169 ( .A(n44239), .Y(n44112) );
  INVX1 U46170 ( .A(n44238), .Y(n44113) );
  INVX1 U46171 ( .A(n44238), .Y(n44114) );
  INVX1 U46172 ( .A(n44238), .Y(n44115) );
  INVX1 U46173 ( .A(n44237), .Y(n44116) );
  INVX1 U46174 ( .A(n44237), .Y(n44117) );
  INVX1 U46175 ( .A(n44237), .Y(n44118) );
  INVX1 U46176 ( .A(n44236), .Y(n44119) );
  INVX1 U46177 ( .A(n44236), .Y(n44120) );
  INVX1 U46178 ( .A(n44236), .Y(n44121) );
  INVX1 U46179 ( .A(n44235), .Y(n44122) );
  INVX1 U46180 ( .A(n44235), .Y(n44123) );
  INVX1 U46181 ( .A(n44235), .Y(n44124) );
  INVX1 U46182 ( .A(n44234), .Y(n44125) );
  INVX1 U46183 ( .A(n44234), .Y(n44126) );
  INVX1 U46184 ( .A(n44234), .Y(n44127) );
  INVX1 U46185 ( .A(n44232), .Y(n44128) );
  INVX1 U46186 ( .A(n44232), .Y(n44129) );
  INVX1 U46187 ( .A(n44239), .Y(n44130) );
  INVX1 U46188 ( .A(n44241), .Y(n44131) );
  INVX1 U46189 ( .A(n44223), .Y(n44132) );
  INVX1 U46190 ( .A(n44215), .Y(n44133) );
  INVX1 U46191 ( .A(n44214), .Y(n44134) );
  INVX1 U46192 ( .A(n44240), .Y(n44135) );
  INVX1 U46193 ( .A(n44215), .Y(n44136) );
  INVX1 U46194 ( .A(n44233), .Y(n44137) );
  INVX1 U46195 ( .A(rst_i), .Y(n44138) );
  INVX1 U46196 ( .A(n44230), .Y(n44139) );
  INVX1 U46197 ( .A(n44232), .Y(n44140) );
  INVX1 U46198 ( .A(n44246), .Y(n44141) );
  INVX1 U46199 ( .A(n44253), .Y(n44142) );
  INVX1 U46200 ( .A(n44254), .Y(n44143) );
  INVX1 U46201 ( .A(n44245), .Y(n44144) );
  INVX1 U46202 ( .A(n44231), .Y(n44145) );
  INVX1 U46203 ( .A(n44231), .Y(n44146) );
  INVX1 U46204 ( .A(n44231), .Y(n44147) );
  INVX1 U46205 ( .A(n44230), .Y(n44148) );
  INVX1 U46206 ( .A(n44230), .Y(n44149) );
  INVX1 U46207 ( .A(n44229), .Y(n44150) );
  INVX1 U46208 ( .A(n44229), .Y(n44151) );
  INVX1 U46209 ( .A(n44229), .Y(n44152) );
  INVX1 U46210 ( .A(n44228), .Y(n44153) );
  INVX1 U46211 ( .A(n44228), .Y(n44154) );
  INVX1 U46212 ( .A(n44228), .Y(n44155) );
  INVX1 U46213 ( .A(n44227), .Y(n44156) );
  INVX1 U46214 ( .A(n44227), .Y(n44157) );
  INVX1 U46215 ( .A(n44227), .Y(n44158) );
  INVX1 U46216 ( .A(n44226), .Y(n44159) );
  INVX1 U46217 ( .A(n44226), .Y(n44160) );
  INVX1 U46218 ( .A(n44226), .Y(n44161) );
  INVX1 U46219 ( .A(n44225), .Y(n44162) );
  INVX1 U46220 ( .A(n44225), .Y(n44163) );
  INVX1 U46221 ( .A(n44225), .Y(n44164) );
  INVX1 U46222 ( .A(n44224), .Y(n44165) );
  INVX1 U46223 ( .A(n44224), .Y(n44166) );
  INVX1 U46224 ( .A(n44224), .Y(n44167) );
  INVX1 U46225 ( .A(n44223), .Y(n44168) );
  INVX1 U46226 ( .A(n44223), .Y(n44169) );
  INVX1 U46227 ( .A(n44223), .Y(n44170) );
  INVX1 U46228 ( .A(n44222), .Y(n44171) );
  INVX1 U46229 ( .A(n44222), .Y(n44172) );
  INVX1 U46230 ( .A(n44222), .Y(n44173) );
  INVX1 U46231 ( .A(n44221), .Y(n44174) );
  INVX1 U46232 ( .A(n44221), .Y(n44175) );
  INVX1 U46233 ( .A(n44221), .Y(n44176) );
  INVX1 U46234 ( .A(n44220), .Y(n44177) );
  INVX1 U46235 ( .A(n44220), .Y(n44178) );
  INVX1 U46236 ( .A(n44220), .Y(n44179) );
  INVX1 U46237 ( .A(n44219), .Y(n44180) );
  INVX1 U46238 ( .A(n44219), .Y(n44181) );
  INVX1 U46239 ( .A(n44219), .Y(n44182) );
  INVX1 U46240 ( .A(n44218), .Y(n44183) );
  INVX1 U46241 ( .A(n44218), .Y(n44184) );
  INVX1 U46242 ( .A(n44218), .Y(n44185) );
  INVX1 U46243 ( .A(n44217), .Y(n44186) );
  INVX1 U46244 ( .A(n44217), .Y(n44187) );
  INVX1 U46245 ( .A(n44217), .Y(n44188) );
  INVX1 U46246 ( .A(n44243), .Y(n44189) );
  INVX1 U46247 ( .A(n44244), .Y(n44190) );
  INVX1 U46248 ( .A(n44233), .Y(n44191) );
  INVX1 U46249 ( .A(n44235), .Y(n44192) );
  INVX1 U46250 ( .A(n44234), .Y(n44193) );
  INVX1 U46251 ( .A(n44216), .Y(n44194) );
  INVX1 U46252 ( .A(n44233), .Y(n44195) );
  INVX1 U46253 ( .A(n44212), .Y(n44196) );
  INVX1 U46254 ( .A(n44213), .Y(n44197) );
  INVX1 U46255 ( .A(n44216), .Y(n44198) );
  INVX1 U46256 ( .A(n44216), .Y(n44199) );
  INVX1 U46257 ( .A(n44216), .Y(n44200) );
  INVX1 U46258 ( .A(n44215), .Y(n44201) );
  INVX1 U46259 ( .A(n44215), .Y(n44202) );
  INVX1 U46260 ( .A(n44214), .Y(n44203) );
  INVX1 U46261 ( .A(n44214), .Y(n44204) );
  INVX1 U46262 ( .A(n44214), .Y(n44205) );
  INVX1 U46263 ( .A(n44213), .Y(n44206) );
  INVX1 U46264 ( .A(n44213), .Y(n44207) );
  INVX1 U46265 ( .A(n44213), .Y(n44208) );
  INVX1 U46266 ( .A(n44212), .Y(n44209) );
  INVX1 U46267 ( .A(n44212), .Y(n44210) );
  INVX1 U46268 ( .A(n44212), .Y(n44211) );
  INVX1 U46269 ( .A(n44252), .Y(n44212) );
  INVX1 U46270 ( .A(n44252), .Y(n44213) );
  INVX1 U46271 ( .A(n38345), .Y(n44214) );
  INVX1 U46272 ( .A(n38346), .Y(n44215) );
  INVX1 U46273 ( .A(n38347), .Y(n44216) );
  INVX1 U46274 ( .A(n38341), .Y(n44217) );
  INVX1 U46275 ( .A(n38342), .Y(n44218) );
  INVX1 U46276 ( .A(n38343), .Y(n44219) );
  INVX1 U46277 ( .A(n38327), .Y(n44220) );
  INVX1 U46278 ( .A(n38328), .Y(n44221) );
  INVX1 U46279 ( .A(n38325), .Y(n44222) );
  INVX1 U46280 ( .A(n44249), .Y(n44223) );
  INVX1 U46281 ( .A(n44249), .Y(n44224) );
  INVX1 U46282 ( .A(n44249), .Y(n44225) );
  INVX1 U46283 ( .A(n38333), .Y(n44226) );
  INVX1 U46284 ( .A(n38330), .Y(n44227) );
  INVX1 U46285 ( .A(n38331), .Y(n44228) );
  INVX1 U46286 ( .A(n38357), .Y(n44229) );
  INVX1 U46287 ( .A(n38354), .Y(n44230) );
  INVX1 U46288 ( .A(n38355), .Y(n44231) );
  INVX1 U46289 ( .A(n38320), .Y(n44232) );
  INVX1 U46290 ( .A(n38352), .Y(n44233) );
  INVX1 U46291 ( .A(n38349), .Y(n44234) );
  INVX1 U46292 ( .A(n38350), .Y(n44235) );
  INVX1 U46293 ( .A(n38337), .Y(n44236) );
  INVX1 U46294 ( .A(n38338), .Y(n44237) );
  INVX1 U46295 ( .A(n38335), .Y(n44238) );
  INVX1 U46296 ( .A(n38361), .Y(n44239) );
  INVX1 U46297 ( .A(n38362), .Y(n44240) );
  INVX1 U46298 ( .A(n38359), .Y(n44241) );
  INVX1 U46299 ( .A(n44248), .Y(n44242) );
  INVX1 U46300 ( .A(n44248), .Y(n44243) );
  INVX1 U46301 ( .A(n44248), .Y(n44244) );
  INVX1 U46302 ( .A(n44247), .Y(n44245) );
  INVX1 U46303 ( .A(n44247), .Y(n44246) );
  INVX1 U46304 ( .A(n44254), .Y(n44247) );
  INVX1 U46305 ( .A(n44254), .Y(n44248) );
  INVX1 U46306 ( .A(n44253), .Y(n44249) );
  INVX1 U46307 ( .A(n44253), .Y(n44250) );
  INVX1 U46308 ( .A(n44253), .Y(n44251) );
  INVX1 U46309 ( .A(n44242), .Y(n44252) );
  INVX1 U46310 ( .A(n73547), .Y(n44253) );
  INVX1 U46311 ( .A(n73547), .Y(n44254) );
  INVX1 U46312 ( .A(n36758), .Y(n44255) );
  INVX1 U46313 ( .A(n44263), .Y(n44256) );
  INVX1 U46314 ( .A(n36758), .Y(n44257) );
  INVX1 U46315 ( .A(n36758), .Y(n44258) );
  INVX1 U46316 ( .A(n44263), .Y(n44259) );
  INVX1 U46317 ( .A(n44264), .Y(n44260) );
  INVX1 U46318 ( .A(n44255), .Y(n44261) );
  INVX1 U46319 ( .A(n44255), .Y(n44262) );
  INVX1 U46320 ( .A(n44255), .Y(n44263) );
  INVX1 U46321 ( .A(n44256), .Y(n44264) );
  INVX1 U46322 ( .A(n44256), .Y(n44265) );
  INVX1 U46323 ( .A(n37459), .Y(n44266) );
  INVX1 U46324 ( .A(n37459), .Y(n44267) );
  INVX1 U46325 ( .A(n37459), .Y(n44268) );
  INVX1 U46326 ( .A(n44271), .Y(n44269) );
  INVX1 U46327 ( .A(n44271), .Y(n44270) );
  INVX1 U46328 ( .A(n28264), .Y(n44271) );
  INVX1 U46329 ( .A(n42207), .Y(n44272) );
  INVX1 U46330 ( .A(n42207), .Y(n44273) );
  INVX1 U46331 ( .A(n42207), .Y(n44274) );
  INVX1 U46332 ( .A(n42213), .Y(n44275) );
  INVX1 U46333 ( .A(n42213), .Y(n44276) );
  INVX1 U46334 ( .A(n42213), .Y(n44277) );
  INVX1 U46335 ( .A(n42206), .Y(n44278) );
  INVX1 U46336 ( .A(n42206), .Y(n44279) );
  INVX1 U46337 ( .A(n42206), .Y(n44280) );
  INVX1 U46338 ( .A(n42444), .Y(n44281) );
  INVX1 U46339 ( .A(n42444), .Y(n44282) );
  INVX1 U46340 ( .A(n42133), .Y(n44283) );
  INVX1 U46341 ( .A(n42133), .Y(n44284) );
  INVX1 U46342 ( .A(n42133), .Y(n44285) );
  INVX1 U46343 ( .A(n44287), .Y(n44286) );
  INVX1 U46344 ( .A(n42144), .Y(n44287) );
  INVX1 U46345 ( .A(n37449), .Y(n44288) );
  INVX1 U46346 ( .A(n37449), .Y(n44289) );
  INVX1 U46347 ( .A(n37450), .Y(n44290) );
  INVX1 U46348 ( .A(n37450), .Y(n44291) );
  INVX1 U46349 ( .A(n37450), .Y(n44292) );
  INVX1 U46350 ( .A(n42209), .Y(n44293) );
  INVX1 U46351 ( .A(n42209), .Y(n44294) );
  INVX1 U46352 ( .A(n36765), .Y(n44295) );
  INVX1 U46353 ( .A(n36765), .Y(n44296) );
  INVX1 U46354 ( .A(n36765), .Y(n44297) );
  INVX1 U46355 ( .A(n37479), .Y(n44298) );
  INVX1 U46356 ( .A(n37479), .Y(n44299) );
  INVX1 U46357 ( .A(n37479), .Y(n44300) );
  INVX1 U46358 ( .A(n37524), .Y(n44301) );
  INVX1 U46359 ( .A(n37524), .Y(n44302) );
  INVX1 U46360 ( .A(n37524), .Y(n44303) );
  INVX1 U46361 ( .A(n44306), .Y(n44304) );
  INVX1 U46362 ( .A(n44306), .Y(n44305) );
  INVX1 U46363 ( .A(n23761), .Y(n44306) );
  INVX1 U46364 ( .A(n37523), .Y(n44307) );
  INVX1 U46365 ( .A(n37523), .Y(n44308) );
  INVX1 U46366 ( .A(n37523), .Y(n44309) );
  INVX1 U46367 ( .A(n37478), .Y(n44310) );
  INVX1 U46368 ( .A(n37478), .Y(n44311) );
  INVX1 U46369 ( .A(n37478), .Y(n44312) );
  INVX1 U46370 ( .A(n37500), .Y(n44313) );
  INVX1 U46371 ( .A(n37500), .Y(n44314) );
  INVX1 U46372 ( .A(n37500), .Y(n44315) );
  INVX1 U46373 ( .A(n44318), .Y(n44316) );
  INVX1 U46374 ( .A(n44318), .Y(n44317) );
  INVX1 U46375 ( .A(n23541), .Y(n44318) );
  INVX1 U46376 ( .A(n37499), .Y(n44319) );
  INVX1 U46377 ( .A(n37499), .Y(n44320) );
  INVX1 U46378 ( .A(n37499), .Y(n44321) );
  INVX1 U46379 ( .A(n37477), .Y(n44322) );
  INVX1 U46380 ( .A(n37477), .Y(n44323) );
  INVX1 U46381 ( .A(n37477), .Y(n44324) );
  INVX1 U46382 ( .A(n37503), .Y(n44325) );
  INVX1 U46383 ( .A(n37503), .Y(n44326) );
  INVX1 U46384 ( .A(n37503), .Y(n44327) );
  INVX1 U46385 ( .A(n44330), .Y(n44328) );
  INVX1 U46386 ( .A(n44330), .Y(n44329) );
  INVX1 U46387 ( .A(n23321), .Y(n44330) );
  INVX1 U46388 ( .A(n37504), .Y(n44331) );
  INVX1 U46389 ( .A(n37504), .Y(n44332) );
  INVX1 U46390 ( .A(n37504), .Y(n44333) );
  INVX1 U46391 ( .A(n37475), .Y(n44334) );
  INVX1 U46392 ( .A(n37475), .Y(n44335) );
  INVX1 U46393 ( .A(n37475), .Y(n44336) );
  INVX1 U46394 ( .A(n37497), .Y(n44337) );
  INVX1 U46395 ( .A(n37497), .Y(n44338) );
  INVX1 U46396 ( .A(n37497), .Y(n44339) );
  INVX1 U46397 ( .A(n44342), .Y(n44340) );
  INVX1 U46398 ( .A(n44342), .Y(n44341) );
  INVX1 U46399 ( .A(n23107), .Y(n44342) );
  INVX1 U46400 ( .A(n37498), .Y(n44343) );
  INVX1 U46401 ( .A(n37498), .Y(n44344) );
  INVX1 U46402 ( .A(n37498), .Y(n44345) );
  INVX1 U46403 ( .A(n37476), .Y(n44346) );
  INVX1 U46404 ( .A(n37476), .Y(n44347) );
  INVX1 U46405 ( .A(n37476), .Y(n44348) );
  INVX1 U46406 ( .A(n37520), .Y(n44349) );
  INVX1 U46407 ( .A(n37520), .Y(n44350) );
  INVX1 U46408 ( .A(n37520), .Y(n44351) );
  INVX1 U46409 ( .A(n44354), .Y(n44352) );
  INVX1 U46410 ( .A(n44354), .Y(n44353) );
  INVX1 U46411 ( .A(n22887), .Y(n44354) );
  INVX1 U46412 ( .A(n37519), .Y(n44355) );
  INVX1 U46413 ( .A(n37519), .Y(n44356) );
  INVX1 U46414 ( .A(n37519), .Y(n44357) );
  INVX1 U46415 ( .A(n37467), .Y(n44358) );
  INVX1 U46416 ( .A(n37467), .Y(n44359) );
  INVX1 U46417 ( .A(n37467), .Y(n44360) );
  INVX1 U46418 ( .A(n37502), .Y(n44361) );
  INVX1 U46419 ( .A(n37502), .Y(n44362) );
  INVX1 U46420 ( .A(n37502), .Y(n44363) );
  INVX1 U46421 ( .A(n44366), .Y(n44364) );
  INVX1 U46422 ( .A(n44366), .Y(n44365) );
  INVX1 U46423 ( .A(n22667), .Y(n44366) );
  INVX1 U46424 ( .A(n37501), .Y(n44367) );
  INVX1 U46425 ( .A(n37501), .Y(n44368) );
  INVX1 U46426 ( .A(n37501), .Y(n44369) );
  INVX1 U46427 ( .A(n37480), .Y(n44370) );
  INVX1 U46428 ( .A(n37480), .Y(n44371) );
  INVX1 U46429 ( .A(n37480), .Y(n44372) );
  INVX1 U46430 ( .A(n37474), .Y(n44373) );
  INVX1 U46431 ( .A(n37474), .Y(n44374) );
  INVX1 U46432 ( .A(n37474), .Y(n44375) );
  INVX1 U46433 ( .A(n37492), .Y(n44376) );
  INVX1 U46434 ( .A(n37492), .Y(n44377) );
  INVX1 U46435 ( .A(n37492), .Y(n44378) );
  INVX1 U46436 ( .A(n37529), .Y(n44379) );
  INVX1 U46437 ( .A(n37529), .Y(n44380) );
  INVX1 U46438 ( .A(n37529), .Y(n44381) );
  INVX1 U46439 ( .A(n44384), .Y(n44382) );
  INVX1 U46440 ( .A(n44384), .Y(n44383) );
  INVX1 U46441 ( .A(n22425), .Y(n44384) );
  INVX1 U46442 ( .A(n37530), .Y(n44385) );
  INVX1 U46443 ( .A(n37530), .Y(n44386) );
  INVX1 U46444 ( .A(n37530), .Y(n44387) );
  INVX1 U46445 ( .A(n37493), .Y(n44388) );
  INVX1 U46446 ( .A(n37493), .Y(n44389) );
  INVX1 U46447 ( .A(n37493), .Y(n44390) );
  INVX1 U46448 ( .A(n37513), .Y(n44391) );
  INVX1 U46449 ( .A(n37513), .Y(n44392) );
  INVX1 U46450 ( .A(n37513), .Y(n44393) );
  INVX1 U46451 ( .A(n44396), .Y(n44394) );
  INVX1 U46452 ( .A(n44396), .Y(n44395) );
  INVX1 U46453 ( .A(n22229), .Y(n44396) );
  INVX1 U46454 ( .A(n37514), .Y(n44397) );
  INVX1 U46455 ( .A(n37514), .Y(n44398) );
  INVX1 U46456 ( .A(n37514), .Y(n44399) );
  INVX1 U46457 ( .A(n37494), .Y(n44400) );
  INVX1 U46458 ( .A(n37494), .Y(n44401) );
  INVX1 U46459 ( .A(n37494), .Y(n44402) );
  INVX1 U46460 ( .A(n37505), .Y(n44403) );
  INVX1 U46461 ( .A(n37505), .Y(n44404) );
  INVX1 U46462 ( .A(n37505), .Y(n44405) );
  INVX1 U46463 ( .A(n44408), .Y(n44406) );
  INVX1 U46464 ( .A(n44408), .Y(n44407) );
  INVX1 U46465 ( .A(n22033), .Y(n44408) );
  INVX1 U46466 ( .A(n37506), .Y(n44409) );
  INVX1 U46467 ( .A(n37506), .Y(n44410) );
  INVX1 U46468 ( .A(n37506), .Y(n44411) );
  INVX1 U46469 ( .A(n37490), .Y(n44412) );
  INVX1 U46470 ( .A(n37490), .Y(n44413) );
  INVX1 U46471 ( .A(n37490), .Y(n44414) );
  INVX1 U46472 ( .A(n37511), .Y(n44415) );
  INVX1 U46473 ( .A(n37511), .Y(n44416) );
  INVX1 U46474 ( .A(n37511), .Y(n44417) );
  INVX1 U46475 ( .A(n44420), .Y(n44418) );
  INVX1 U46476 ( .A(n44420), .Y(n44419) );
  INVX1 U46477 ( .A(n21837), .Y(n44420) );
  INVX1 U46478 ( .A(n37512), .Y(n44421) );
  INVX1 U46479 ( .A(n37512), .Y(n44422) );
  INVX1 U46480 ( .A(n37512), .Y(n44423) );
  INVX1 U46481 ( .A(n37491), .Y(n44424) );
  INVX1 U46482 ( .A(n37491), .Y(n44425) );
  INVX1 U46483 ( .A(n37491), .Y(n44426) );
  INVX1 U46484 ( .A(n37527), .Y(n44427) );
  INVX1 U46485 ( .A(n37527), .Y(n44428) );
  INVX1 U46486 ( .A(n37527), .Y(n44429) );
  INVX1 U46487 ( .A(n44432), .Y(n44430) );
  INVX1 U46488 ( .A(n44432), .Y(n44431) );
  INVX1 U46489 ( .A(n21641), .Y(n44432) );
  INVX1 U46490 ( .A(n37528), .Y(n44433) );
  INVX1 U46491 ( .A(n37528), .Y(n44434) );
  INVX1 U46492 ( .A(n37528), .Y(n44435) );
  INVX1 U46493 ( .A(n37470), .Y(n44436) );
  INVX1 U46494 ( .A(n37470), .Y(n44437) );
  INVX1 U46495 ( .A(n37470), .Y(n44438) );
  INVX1 U46496 ( .A(n37508), .Y(n44439) );
  INVX1 U46497 ( .A(n37508), .Y(n44440) );
  INVX1 U46498 ( .A(n37508), .Y(n44441) );
  INVX1 U46499 ( .A(n44444), .Y(n44442) );
  INVX1 U46500 ( .A(n44444), .Y(n44443) );
  INVX1 U46501 ( .A(n21445), .Y(n44444) );
  INVX1 U46502 ( .A(n37507), .Y(n44445) );
  INVX1 U46503 ( .A(n37507), .Y(n44446) );
  INVX1 U46504 ( .A(n37507), .Y(n44447) );
  INVX1 U46505 ( .A(n37465), .Y(n44448) );
  INVX1 U46506 ( .A(n37465), .Y(n44449) );
  INVX1 U46507 ( .A(n37465), .Y(n44450) );
  INVX1 U46508 ( .A(n37458), .Y(n44451) );
  INVX1 U46509 ( .A(n37458), .Y(n44452) );
  INVX1 U46510 ( .A(n37458), .Y(n44453) );
  INVX1 U46511 ( .A(n37466), .Y(n44454) );
  INVX1 U46512 ( .A(n37466), .Y(n44455) );
  INVX1 U46513 ( .A(n37466), .Y(n44456) );
  INVX1 U46514 ( .A(n37463), .Y(n44457) );
  INVX1 U46515 ( .A(n37463), .Y(n44458) );
  INVX1 U46516 ( .A(n37463), .Y(n44459) );
  INVX1 U46517 ( .A(n44462), .Y(n44460) );
  INVX1 U46518 ( .A(n44462), .Y(n44461) );
  INVX1 U46519 ( .A(n21051), .Y(n44462) );
  INVX1 U46520 ( .A(n37462), .Y(n44463) );
  INVX1 U46521 ( .A(n37462), .Y(n44464) );
  INVX1 U46522 ( .A(n37462), .Y(n44465) );
  INVX1 U46523 ( .A(n37486), .Y(n44466) );
  INVX1 U46524 ( .A(n37486), .Y(n44467) );
  INVX1 U46525 ( .A(n37486), .Y(n44468) );
  INVX1 U46526 ( .A(n37526), .Y(n44469) );
  INVX1 U46527 ( .A(n37526), .Y(n44470) );
  INVX1 U46528 ( .A(n37526), .Y(n44471) );
  INVX1 U46529 ( .A(n37584), .Y(n44472) );
  INVX1 U46530 ( .A(n37584), .Y(n44473) );
  INVX1 U46531 ( .A(n37584), .Y(n44474) );
  INVX1 U46532 ( .A(n37525), .Y(n44475) );
  INVX1 U46533 ( .A(n37525), .Y(n44476) );
  INVX1 U46534 ( .A(n37525), .Y(n44477) );
  INVX1 U46535 ( .A(n37487), .Y(n44478) );
  INVX1 U46536 ( .A(n37487), .Y(n44479) );
  INVX1 U46537 ( .A(n37487), .Y(n44480) );
  INVX1 U46538 ( .A(n37518), .Y(n44481) );
  INVX1 U46539 ( .A(n37518), .Y(n44482) );
  INVX1 U46540 ( .A(n37518), .Y(n44483) );
  INVX1 U46541 ( .A(n44486), .Y(n44484) );
  INVX1 U46542 ( .A(n44486), .Y(n44485) );
  INVX1 U46543 ( .A(n20659), .Y(n44486) );
  INVX1 U46544 ( .A(n37517), .Y(n44487) );
  INVX1 U46545 ( .A(n37517), .Y(n44488) );
  INVX1 U46546 ( .A(n37517), .Y(n44489) );
  INVX1 U46547 ( .A(n37481), .Y(n44490) );
  INVX1 U46548 ( .A(n37481), .Y(n44491) );
  INVX1 U46549 ( .A(n37481), .Y(n44492) );
  INVX1 U46550 ( .A(n37468), .Y(n44493) );
  INVX1 U46551 ( .A(n37468), .Y(n44494) );
  INVX1 U46552 ( .A(n37468), .Y(n44495) );
  INVX1 U46553 ( .A(n37488), .Y(n44496) );
  INVX1 U46554 ( .A(n37488), .Y(n44497) );
  INVX1 U46555 ( .A(n37488), .Y(n44498) );
  INVX1 U46556 ( .A(n37515), .Y(n44499) );
  INVX1 U46557 ( .A(n37515), .Y(n44500) );
  INVX1 U46558 ( .A(n37515), .Y(n44501) );
  INVX1 U46559 ( .A(n44504), .Y(n44502) );
  INVX1 U46560 ( .A(n44504), .Y(n44503) );
  INVX1 U46561 ( .A(n20267), .Y(n44504) );
  INVX1 U46562 ( .A(n37516), .Y(n44505) );
  INVX1 U46563 ( .A(n37516), .Y(n44506) );
  INVX1 U46564 ( .A(n37516), .Y(n44507) );
  INVX1 U46565 ( .A(n37489), .Y(n44508) );
  INVX1 U46566 ( .A(n37489), .Y(n44509) );
  INVX1 U46567 ( .A(n37489), .Y(n44510) );
  INVX1 U46568 ( .A(n37522), .Y(n44511) );
  INVX1 U46569 ( .A(n37522), .Y(n44512) );
  INVX1 U46570 ( .A(n37522), .Y(n44513) );
  INVX1 U46571 ( .A(n44516), .Y(n44514) );
  INVX1 U46572 ( .A(n44516), .Y(n44515) );
  INVX1 U46573 ( .A(n20071), .Y(n44516) );
  INVX1 U46574 ( .A(n37521), .Y(n44517) );
  INVX1 U46575 ( .A(n37521), .Y(n44518) );
  INVX1 U46576 ( .A(n37521), .Y(n44519) );
  INVX1 U46577 ( .A(n37471), .Y(n44520) );
  INVX1 U46578 ( .A(n37471), .Y(n44521) );
  INVX1 U46579 ( .A(n37471), .Y(n44522) );
  INVX1 U46580 ( .A(n37510), .Y(n44523) );
  INVX1 U46581 ( .A(n37510), .Y(n44524) );
  INVX1 U46582 ( .A(n37510), .Y(n44525) );
  INVX1 U46583 ( .A(n44528), .Y(n44526) );
  INVX1 U46584 ( .A(n44528), .Y(n44527) );
  INVX1 U46585 ( .A(n19875), .Y(n44528) );
  INVX1 U46586 ( .A(n37509), .Y(n44529) );
  INVX1 U46587 ( .A(n37509), .Y(n44530) );
  INVX1 U46588 ( .A(n37509), .Y(n44531) );
  INVX1 U46589 ( .A(n37484), .Y(n44532) );
  INVX1 U46590 ( .A(n37484), .Y(n44533) );
  INVX1 U46591 ( .A(n37484), .Y(n44534) );
  INVX1 U46592 ( .A(n42599), .Y(n44535) );
  INVX1 U46593 ( .A(n42599), .Y(n44536) );
  INVX1 U46594 ( .A(n42599), .Y(n44537) );
  INVX1 U46595 ( .A(n44540), .Y(n44538) );
  INVX1 U46596 ( .A(n44540), .Y(n44539) );
  INVX1 U46597 ( .A(n19678), .Y(n44540) );
  INVX1 U46598 ( .A(n37532), .Y(n44541) );
  INVX1 U46599 ( .A(n37532), .Y(n44542) );
  INVX1 U46600 ( .A(n37532), .Y(n44543) );
  INVX1 U46601 ( .A(n37464), .Y(n44544) );
  INVX1 U46602 ( .A(n37464), .Y(n44545) );
  INVX1 U46603 ( .A(n37464), .Y(n44546) );
  INVX1 U46604 ( .A(n37457), .Y(n44547) );
  INVX1 U46605 ( .A(n37457), .Y(n44548) );
  INVX1 U46606 ( .A(n37457), .Y(n44549) );
  INVX1 U46607 ( .A(n44552), .Y(n44550) );
  INVX1 U46608 ( .A(n44552), .Y(n44551) );
  INVX1 U46609 ( .A(n19481), .Y(n44552) );
  INVX1 U46610 ( .A(n37456), .Y(n44553) );
  INVX1 U46611 ( .A(n37456), .Y(n44554) );
  INVX1 U46612 ( .A(n37456), .Y(n44555) );
  INVX1 U46613 ( .A(n37535), .Y(n44556) );
  INVX1 U46614 ( .A(n37535), .Y(n44557) );
  INVX1 U46615 ( .A(n37535), .Y(n44558) );
  INVX1 U46616 ( .A(n37579), .Y(n44559) );
  INVX1 U46617 ( .A(n37579), .Y(n44560) );
  INVX1 U46618 ( .A(n37579), .Y(n44561) );
  INVX1 U46619 ( .A(n37496), .Y(n44562) );
  INVX1 U46620 ( .A(n37496), .Y(n44563) );
  INVX1 U46621 ( .A(n37496), .Y(n44564) );
  INVX1 U46622 ( .A(n44567), .Y(n44565) );
  INVX1 U46623 ( .A(n44567), .Y(n44566) );
  INVX1 U46624 ( .A(n19088), .Y(n44567) );
  INVX1 U46625 ( .A(n37534), .Y(n44568) );
  INVX1 U46626 ( .A(n37534), .Y(n44569) );
  INVX1 U46627 ( .A(n37534), .Y(n44570) );
  INVX1 U46628 ( .A(n37580), .Y(n44571) );
  INVX1 U46629 ( .A(n37580), .Y(n44572) );
  INVX1 U46630 ( .A(n37580), .Y(n44573) );
  INVX1 U46631 ( .A(n37495), .Y(n44574) );
  INVX1 U46632 ( .A(n37495), .Y(n44575) );
  INVX1 U46633 ( .A(n37495), .Y(n44576) );
  INVX1 U46634 ( .A(n44579), .Y(n44577) );
  INVX1 U46635 ( .A(n44579), .Y(n44578) );
  INVX1 U46636 ( .A(n18696), .Y(n44579) );
  INVX1 U46637 ( .A(n37536), .Y(n44580) );
  INVX1 U46638 ( .A(n37536), .Y(n44581) );
  INVX1 U46639 ( .A(n37536), .Y(n44582) );
  INVX1 U46640 ( .A(n37581), .Y(n44583) );
  INVX1 U46641 ( .A(n37581), .Y(n44584) );
  INVX1 U46642 ( .A(n37581), .Y(n44585) );
  INVX1 U46643 ( .A(n37460), .Y(n44586) );
  INVX1 U46644 ( .A(n37460), .Y(n44587) );
  INVX1 U46645 ( .A(n37460), .Y(n44588) );
  INVX1 U46646 ( .A(n37455), .Y(n44589) );
  INVX1 U46647 ( .A(n37455), .Y(n44590) );
  INVX1 U46648 ( .A(n37455), .Y(n44591) );
  INVX1 U46649 ( .A(n44594), .Y(n44592) );
  INVX1 U46650 ( .A(n44594), .Y(n44593) );
  INVX1 U46651 ( .A(n18305), .Y(n44594) );
  INVX1 U46652 ( .A(n37454), .Y(n44595) );
  INVX1 U46653 ( .A(n37454), .Y(n44596) );
  INVX1 U46654 ( .A(n37454), .Y(n44597) );
  INVX1 U46655 ( .A(n42604), .Y(n44598) );
  INVX1 U46656 ( .A(n42604), .Y(n44599) );
  INVX1 U46657 ( .A(n42604), .Y(n44600) );
  INVX1 U46658 ( .A(n37577), .Y(n44601) );
  INVX1 U46659 ( .A(n37577), .Y(n44602) );
  INVX1 U46660 ( .A(n37577), .Y(n44603) );
  INVX1 U46661 ( .A(n42605), .Y(n44604) );
  INVX1 U46662 ( .A(n42605), .Y(n44605) );
  INVX1 U46663 ( .A(n42605), .Y(n44606) );
  INVX1 U46664 ( .A(n44609), .Y(n44607) );
  INVX1 U46665 ( .A(n44609), .Y(n44608) );
  INVX1 U46666 ( .A(n18002), .Y(n44609) );
  INVX1 U46667 ( .A(n44619), .Y(n44610) );
  INVX1 U46668 ( .A(n44626), .Y(n44611) );
  INVX1 U46669 ( .A(n44620), .Y(n44612) );
  INVX1 U46670 ( .A(n44623), .Y(n44613) );
  INVX1 U46671 ( .A(n44619), .Y(n44614) );
  INVX1 U46672 ( .A(n44619), .Y(n44615) );
  INVX1 U46673 ( .A(n44619), .Y(n44616) );
  INVX1 U46674 ( .A(n44619), .Y(n44617) );
  INVX1 U46675 ( .A(n44619), .Y(n44618) );
  INVX1 U46676 ( .A(n44627), .Y(n44619) );
  INVX1 U46677 ( .A(n44627), .Y(n44620) );
  INVX1 U46678 ( .A(n44627), .Y(n44621) );
  INVX1 U46679 ( .A(n44627), .Y(n44622) );
  INVX1 U46680 ( .A(n44627), .Y(n44623) );
  INVX1 U46681 ( .A(n42598), .Y(n44624) );
  INVX1 U46682 ( .A(n44627), .Y(n44625) );
  INVX1 U46683 ( .A(n44627), .Y(n44626) );
  INVX1 U46684 ( .A(n44624), .Y(n44627) );
  INVX1 U46685 ( .A(n37575), .Y(n44628) );
  INVX1 U46686 ( .A(n37575), .Y(n44629) );
  INVX1 U46687 ( .A(n37575), .Y(n44630) );
  INVX1 U46688 ( .A(n37333), .Y(n44631) );
  INVX1 U46689 ( .A(n37333), .Y(n44632) );
  INVX1 U46690 ( .A(n37333), .Y(n44633) );
  INVX1 U46691 ( .A(n40930), .Y(n44634) );
  INVX1 U46692 ( .A(n40930), .Y(n44635) );
  INVX1 U46693 ( .A(n40930), .Y(n44636) );
  INVX1 U46694 ( .A(n40930), .Y(n44637) );
  INVX1 U46695 ( .A(n40930), .Y(n44638) );
  INVX1 U46696 ( .A(n8805), .Y(n44639) );
  INVX1 U46697 ( .A(n8805), .Y(n44640) );
  INVX1 U46698 ( .A(writeback_csr_value_w[30]), .Y(n44641) );
  INVX1 U46699 ( .A(writeback_csr_value_w[30]), .Y(n44642) );
  INVX1 U46700 ( .A(writeback_csr_value_w[15]), .Y(n44643) );
  INVX1 U46701 ( .A(writeback_csr_value_w[15]), .Y(n44644) );
  INVX1 U46702 ( .A(writeback_csr_value_w[14]), .Y(n44645) );
  INVX1 U46703 ( .A(writeback_csr_value_w[14]), .Y(n44646) );
  INVX1 U46704 ( .A(writeback_csr_value_w[29]), .Y(n44647) );
  INVX1 U46705 ( .A(writeback_csr_value_w[29]), .Y(n44648) );
  INVX1 U46706 ( .A(writeback_csr_value_w[28]), .Y(n44649) );
  INVX1 U46707 ( .A(writeback_csr_value_w[28]), .Y(n44650) );
  INVX1 U46708 ( .A(writeback_csr_value_w[19]), .Y(n44651) );
  INVX1 U46709 ( .A(writeback_csr_value_w[19]), .Y(n44652) );
  INVX1 U46710 ( .A(writeback_csr_value_w[20]), .Y(n44653) );
  INVX1 U46711 ( .A(writeback_csr_value_w[20]), .Y(n44654) );
  INVX1 U46712 ( .A(writeback_csr_value_w[23]), .Y(n44655) );
  INVX1 U46713 ( .A(writeback_csr_value_w[23]), .Y(n44656) );
  INVX1 U46714 ( .A(writeback_csr_value_w[22]), .Y(n44657) );
  INVX1 U46715 ( .A(writeback_csr_value_w[22]), .Y(n44658) );
  INVX1 U46716 ( .A(writeback_csr_value_w[16]), .Y(n44659) );
  INVX1 U46717 ( .A(writeback_csr_value_w[16]), .Y(n44660) );
  INVX1 U46718 ( .A(writeback_csr_value_w[21]), .Y(n44661) );
  INVX1 U46719 ( .A(writeback_csr_value_w[21]), .Y(n44662) );
  INVX1 U46720 ( .A(writeback_csr_value_w[26]), .Y(n44663) );
  INVX1 U46721 ( .A(writeback_csr_value_w[26]), .Y(n44664) );
  INVX1 U46722 ( .A(writeback_csr_value_w[18]), .Y(n44665) );
  INVX1 U46723 ( .A(writeback_csr_value_w[18]), .Y(n44666) );
  INVX1 U46724 ( .A(writeback_csr_value_w[12]), .Y(n44667) );
  INVX1 U46725 ( .A(writeback_csr_value_w[12]), .Y(n44668) );
  INVX1 U46726 ( .A(writeback_csr_value_w[13]), .Y(n44669) );
  INVX1 U46727 ( .A(writeback_csr_value_w[13]), .Y(n44670) );
  INVX1 U46728 ( .A(writeback_csr_value_w[27]), .Y(n44671) );
  INVX1 U46729 ( .A(writeback_csr_value_w[27]), .Y(n44672) );
  INVX1 U46730 ( .A(writeback_csr_value_w[25]), .Y(n44673) );
  INVX1 U46731 ( .A(writeback_csr_value_w[25]), .Y(n44674) );
  INVX1 U46732 ( .A(writeback_csr_value_w[24]), .Y(n44675) );
  INVX1 U46733 ( .A(writeback_csr_value_w[24]), .Y(n44676) );
  INVX1 U46734 ( .A(writeback_csr_value_w[17]), .Y(n44677) );
  INVX1 U46735 ( .A(writeback_csr_value_w[17]), .Y(n44678) );
  INVX1 U46736 ( .A(writeback_csr_value_w[31]), .Y(n44679) );
  INVX1 U46737 ( .A(writeback_csr_value_w[31]), .Y(n44680) );
  INVX1 U46738 ( .A(writeback_csr_value_w[0]), .Y(n44681) );
  INVX1 U46739 ( .A(writeback_csr_value_w[0]), .Y(n44682) );
  INVX1 U46740 ( .A(writeback_csr_value_w[1]), .Y(n44683) );
  INVX1 U46741 ( .A(writeback_csr_value_w[1]), .Y(n44684) );
  INVX1 U46742 ( .A(writeback_csr_value_w[2]), .Y(n44685) );
  INVX1 U46743 ( .A(writeback_csr_value_w[2]), .Y(n44686) );
  INVX1 U46744 ( .A(writeback_csr_value_w[3]), .Y(n44687) );
  INVX1 U46745 ( .A(writeback_csr_value_w[3]), .Y(n44688) );
  INVX1 U46746 ( .A(writeback_csr_value_w[4]), .Y(n44689) );
  INVX1 U46747 ( .A(writeback_csr_value_w[4]), .Y(n44690) );
  INVX1 U46748 ( .A(writeback_csr_value_w[5]), .Y(n44691) );
  INVX1 U46749 ( .A(writeback_csr_value_w[5]), .Y(n44692) );
  INVX1 U46750 ( .A(writeback_csr_value_w[11]), .Y(n44693) );
  INVX1 U46751 ( .A(writeback_csr_value_w[11]), .Y(n44694) );
  INVX1 U46752 ( .A(writeback_csr_value_w[6]), .Y(n44695) );
  INVX1 U46753 ( .A(writeback_csr_value_w[6]), .Y(n44696) );
  INVX1 U46754 ( .A(writeback_csr_value_w[10]), .Y(n44697) );
  INVX1 U46755 ( .A(writeback_csr_value_w[10]), .Y(n44698) );
  INVX1 U46756 ( .A(writeback_csr_value_w[9]), .Y(n44699) );
  INVX1 U46757 ( .A(writeback_csr_value_w[9]), .Y(n44700) );
  INVX1 U46758 ( .A(writeback_csr_value_w[7]), .Y(n44701) );
  INVX1 U46759 ( .A(writeback_csr_value_w[7]), .Y(n44702) );
  INVX1 U46760 ( .A(writeback_csr_value_w[8]), .Y(n44703) );
  INVX1 U46761 ( .A(writeback_csr_value_w[8]), .Y(n44704) );
  INVX1 U46762 ( .A(writeback_muldiv_value_w[30]), .Y(n44705) );
  INVX1 U46763 ( .A(writeback_muldiv_value_w[30]), .Y(n44706) );
  INVX1 U46764 ( .A(writeback_muldiv_value_w[31]), .Y(n44707) );
  INVX1 U46765 ( .A(writeback_muldiv_value_w[31]), .Y(n44708) );
  INVX1 U46766 ( .A(writeback_muldiv_value_w[15]), .Y(n44709) );
  INVX1 U46767 ( .A(writeback_muldiv_value_w[15]), .Y(n44710) );
  INVX1 U46768 ( .A(writeback_muldiv_value_w[14]), .Y(n44711) );
  INVX1 U46769 ( .A(writeback_muldiv_value_w[14]), .Y(n44712) );
  INVX1 U46770 ( .A(writeback_muldiv_value_w[29]), .Y(n44713) );
  INVX1 U46771 ( .A(writeback_muldiv_value_w[29]), .Y(n44714) );
  INVX1 U46772 ( .A(writeback_muldiv_value_w[28]), .Y(n44715) );
  INVX1 U46773 ( .A(writeback_muldiv_value_w[28]), .Y(n44716) );
  INVX1 U46774 ( .A(writeback_muldiv_value_w[19]), .Y(n44717) );
  INVX1 U46775 ( .A(writeback_muldiv_value_w[19]), .Y(n44718) );
  INVX1 U46776 ( .A(writeback_muldiv_value_w[20]), .Y(n44719) );
  INVX1 U46777 ( .A(writeback_muldiv_value_w[20]), .Y(n44720) );
  INVX1 U46778 ( .A(writeback_muldiv_value_w[23]), .Y(n44721) );
  INVX1 U46779 ( .A(writeback_muldiv_value_w[23]), .Y(n44722) );
  INVX1 U46780 ( .A(writeback_muldiv_value_w[22]), .Y(n44723) );
  INVX1 U46781 ( .A(writeback_muldiv_value_w[22]), .Y(n44724) );
  INVX1 U46782 ( .A(writeback_muldiv_value_w[16]), .Y(n44725) );
  INVX1 U46783 ( .A(writeback_muldiv_value_w[16]), .Y(n44726) );
  INVX1 U46784 ( .A(writeback_muldiv_value_w[21]), .Y(n44727) );
  INVX1 U46785 ( .A(writeback_muldiv_value_w[21]), .Y(n44728) );
  INVX1 U46786 ( .A(writeback_muldiv_value_w[26]), .Y(n44729) );
  INVX1 U46787 ( .A(writeback_muldiv_value_w[26]), .Y(n44730) );
  INVX1 U46788 ( .A(writeback_muldiv_value_w[18]), .Y(n44731) );
  INVX1 U46789 ( .A(writeback_muldiv_value_w[18]), .Y(n44732) );
  INVX1 U46790 ( .A(writeback_muldiv_value_w[12]), .Y(n44733) );
  INVX1 U46791 ( .A(writeback_muldiv_value_w[12]), .Y(n44734) );
  INVX1 U46792 ( .A(writeback_muldiv_value_w[13]), .Y(n44735) );
  INVX1 U46793 ( .A(writeback_muldiv_value_w[13]), .Y(n44736) );
  INVX1 U46794 ( .A(writeback_muldiv_value_w[27]), .Y(n44737) );
  INVX1 U46795 ( .A(writeback_muldiv_value_w[27]), .Y(n44738) );
  INVX1 U46796 ( .A(writeback_muldiv_value_w[25]), .Y(n44739) );
  INVX1 U46797 ( .A(writeback_muldiv_value_w[25]), .Y(n44740) );
  INVX1 U46798 ( .A(writeback_muldiv_value_w[24]), .Y(n44741) );
  INVX1 U46799 ( .A(writeback_muldiv_value_w[24]), .Y(n44742) );
  INVX1 U46800 ( .A(writeback_muldiv_value_w[17]), .Y(n44743) );
  INVX1 U46801 ( .A(writeback_muldiv_value_w[17]), .Y(n44744) );
  INVX1 U46802 ( .A(writeback_muldiv_value_w[0]), .Y(n44745) );
  INVX1 U46803 ( .A(writeback_muldiv_value_w[0]), .Y(n44746) );
  INVX1 U46804 ( .A(writeback_muldiv_value_w[5]), .Y(n44747) );
  INVX1 U46805 ( .A(writeback_muldiv_value_w[5]), .Y(n44748) );
  INVX1 U46806 ( .A(writeback_muldiv_value_w[1]), .Y(n44749) );
  INVX1 U46807 ( .A(writeback_muldiv_value_w[1]), .Y(n44750) );
  INVX1 U46808 ( .A(writeback_muldiv_value_w[4]), .Y(n44751) );
  INVX1 U46809 ( .A(writeback_muldiv_value_w[4]), .Y(n44752) );
  INVX1 U46810 ( .A(writeback_muldiv_value_w[3]), .Y(n44753) );
  INVX1 U46811 ( .A(writeback_muldiv_value_w[3]), .Y(n44754) );
  INVX1 U46812 ( .A(writeback_muldiv_value_w[2]), .Y(n44755) );
  INVX1 U46813 ( .A(writeback_muldiv_value_w[2]), .Y(n44756) );
  INVX1 U46814 ( .A(writeback_muldiv_value_w[11]), .Y(n44757) );
  INVX1 U46815 ( .A(writeback_muldiv_value_w[11]), .Y(n44758) );
  INVX1 U46816 ( .A(writeback_muldiv_value_w[6]), .Y(n44759) );
  INVX1 U46817 ( .A(writeback_muldiv_value_w[6]), .Y(n44760) );
  INVX1 U46818 ( .A(writeback_muldiv_value_w[10]), .Y(n44761) );
  INVX1 U46819 ( .A(writeback_muldiv_value_w[10]), .Y(n44762) );
  INVX1 U46820 ( .A(writeback_muldiv_value_w[9]), .Y(n44763) );
  INVX1 U46821 ( .A(writeback_muldiv_value_w[9]), .Y(n44764) );
  INVX1 U46822 ( .A(writeback_muldiv_value_w[7]), .Y(n44765) );
  INVX1 U46823 ( .A(writeback_muldiv_value_w[7]), .Y(n44766) );
  INVX1 U46824 ( .A(writeback_muldiv_value_w[8]), .Y(n44767) );
  INVX1 U46825 ( .A(writeback_muldiv_value_w[8]), .Y(n44768) );
  INVX1 U46826 ( .A(n19276), .Y(n44769) );
  INVX1 U46827 ( .A(n19276), .Y(n44770) );
  INVX1 U46828 ( .A(n19276), .Y(n44771) );
  INVX1 U46829 ( .A(n19279), .Y(n44772) );
  INVX1 U46830 ( .A(n19279), .Y(n44773) );
  INVX1 U46831 ( .A(n19279), .Y(n44774) );
  INVX1 U46832 ( .A(n18884), .Y(n44775) );
  INVX1 U46833 ( .A(n18884), .Y(n44776) );
  INVX1 U46834 ( .A(n18884), .Y(n44777) );
  INVX1 U46835 ( .A(n18887), .Y(n44778) );
  INVX1 U46836 ( .A(n18887), .Y(n44779) );
  INVX1 U46837 ( .A(n18887), .Y(n44780) );
  INVX1 U46838 ( .A(n19472), .Y(n44781) );
  INVX1 U46839 ( .A(n19472), .Y(n44782) );
  INVX1 U46840 ( .A(n19475), .Y(n44783) );
  INVX1 U46841 ( .A(n19475), .Y(n44784) );
  INVX1 U46842 ( .A(n18688), .Y(n44785) );
  INVX1 U46843 ( .A(n18688), .Y(n44786) );
  INVX1 U46844 ( .A(n18688), .Y(n44787) );
  INVX1 U46845 ( .A(n18691), .Y(n44788) );
  INVX1 U46846 ( .A(n18691), .Y(n44789) );
  INVX1 U46847 ( .A(n18691), .Y(n44790) );
  INVX1 U46848 ( .A(n19080), .Y(n44791) );
  INVX1 U46849 ( .A(n19080), .Y(n44792) );
  INVX1 U46850 ( .A(n19080), .Y(n44793) );
  INVX1 U46851 ( .A(n19083), .Y(n44794) );
  INVX1 U46852 ( .A(n19083), .Y(n44795) );
  INVX1 U46853 ( .A(n19083), .Y(n44796) );
  INVX1 U46854 ( .A(n18295), .Y(n44797) );
  INVX1 U46855 ( .A(n18295), .Y(n44798) );
  INVX1 U46856 ( .A(n18295), .Y(n44799) );
  INVX1 U46857 ( .A(n18299), .Y(n44800) );
  INVX1 U46858 ( .A(n18299), .Y(n44801) );
  INVX1 U46859 ( .A(n18299), .Y(n44802) );
  INVX1 U46860 ( .A(n24100), .Y(n44803) );
  INVX1 U46861 ( .A(n24100), .Y(n44804) );
  INVX1 U46862 ( .A(n24100), .Y(n44805) );
  INVX1 U46863 ( .A(n24104), .Y(n44806) );
  INVX1 U46864 ( .A(n24104), .Y(n44807) );
  INVX1 U46865 ( .A(n24104), .Y(n44808) );
  INVX1 U46866 ( .A(n44810), .Y(n44809) );
  INVX1 U46867 ( .A(n44818), .Y(n44811) );
  INVX1 U46868 ( .A(n44810), .Y(n44812) );
  INVX1 U46869 ( .A(n44818), .Y(n44813) );
  INVX1 U46870 ( .A(n44809), .Y(n44814) );
  INVX1 U46871 ( .A(n44809), .Y(n44815) );
  INVX1 U46872 ( .A(n44809), .Y(n44816) );
  INVX1 U46873 ( .A(n44809), .Y(n44817) );
  INVX1 U46874 ( .A(n36761), .Y(n44818) );
  INVX1 U46875 ( .A(n44821), .Y(n44819) );
  INVX1 U46876 ( .A(n44821), .Y(n44820) );
  INVX1 U46877 ( .A(u_muldiv_div_inst_q), .Y(n44821) );
  INVX1 U46878 ( .A(n44828), .Y(n44822) );
  INVX1 U46879 ( .A(n44824), .Y(n44823) );
  INVX1 U46880 ( .A(n44819), .Y(n44824) );
  INVX1 U46881 ( .A(n44819), .Y(n44825) );
  INVX1 U46882 ( .A(n44819), .Y(n44826) );
  INVX1 U46883 ( .A(n44820), .Y(n44827) );
  INVX1 U46884 ( .A(n44820), .Y(n44828) );
  INVX1 U46885 ( .A(n44820), .Y(n44829) );
  INVX1 U46886 ( .A(n44819), .Y(n44830) );
  INVX1 U46887 ( .A(n44832), .Y(n44831) );
  INVX1 U46888 ( .A(n44832), .Y(n44833) );
  INVX1 U46889 ( .A(n42850), .Y(n44834) );
  INVX1 U46890 ( .A(n44839), .Y(n44835) );
  INVX1 U46891 ( .A(n44839), .Y(n44836) );
  INVX1 U46892 ( .A(n44843), .Y(n44837) );
  INVX1 U46893 ( .A(n44841), .Y(n44838) );
  INVX1 U46894 ( .A(opcode_opcode_w[31]), .Y(n44839) );
  INVX1 U46895 ( .A(n44838), .Y(n44840) );
  INVX1 U46896 ( .A(n44831), .Y(n44841) );
  INVX1 U46897 ( .A(n44831), .Y(n44842) );
  INVX1 U46898 ( .A(n44831), .Y(n44843) );
  INVX1 U46899 ( .A(opcode_opcode_w[31]), .Y(n44844) );
  INVX1 U46900 ( .A(n42851), .Y(n44845) );
  INVX1 U46901 ( .A(n44847), .Y(n44846) );
  INVX1 U46902 ( .A(wm_select), .Y(n44847) );
  INVX1 U46903 ( .A(n44847), .Y(n44848) );
  INVX1 U46904 ( .A(n44856), .Y(n44849) );
  INVX1 U46905 ( .A(n44856), .Y(n44850) );
  INVX1 U46906 ( .A(n44856), .Y(n44851) );
  INVX1 U46907 ( .A(n44856), .Y(n44852) );
  INVX1 U46908 ( .A(n44858), .Y(n44853) );
  INVX1 U46909 ( .A(n44856), .Y(n44854) );
  INVX1 U46910 ( .A(n44862), .Y(n44855) );
  INVX1 U46911 ( .A(n44846), .Y(n44856) );
  INVX1 U46912 ( .A(n44846), .Y(n44857) );
  INVX1 U46913 ( .A(wm_select), .Y(n44858) );
  INVX1 U46914 ( .A(wm_select), .Y(n44859) );
  INVX1 U46915 ( .A(wm_select), .Y(n44860) );
  INVX1 U46916 ( .A(n44846), .Y(n44861) );
  INVX1 U46917 ( .A(n44846), .Y(n44862) );
  INVX1 U46918 ( .A(n44846), .Y(n44863) );
  INVX1 U46919 ( .A(clk_i), .Y(n73546) );
  INVX1 U46920 ( .A(mem_d_resp_tag_i[0]), .Y(n73557) );
  INVX1 U46921 ( .A(mem_d_resp_tag_i[1]), .Y(n73556) );
  INVX1 U46922 ( .A(mem_d_resp_tag_i[2]), .Y(n73555) );
  NAND2X1 U46923 ( .A(n36249), .B(mem_d_ack_i), .Y(n28544) );
  INVX1 U46924 ( .A(n28544), .Y(n44990) );
  NAND2X1 U46925 ( .A(mem_d_resp_tag_i[3]), .B(n44990), .Y(n45297) );
  INVX1 U46926 ( .A(n45297), .Y(n45163) );
  NAND2X1 U46927 ( .A(n36247), .B(n44990), .Y(n35922) );
  NOR2X1 U46928 ( .A(mem_d_resp_tag_i[2]), .B(n73556), .Y(n44864) );
  NAND2X1 U46929 ( .A(n44864), .B(n44990), .Y(n45076) );
  INVX1 U46930 ( .A(n45076), .Y(n57519) );
  NAND2X1 U46931 ( .A(n36244), .B(n44990), .Y(n57534) );
  NAND2X1 U46932 ( .A(n57519), .B(n57534), .Y(n24196) );
  INVX1 U46933 ( .A(n35952), .Y(n44865) );
  NOR2X1 U46934 ( .A(n37433), .B(n44865), .Y(n44946) );
  XNOR2X1 U46935 ( .A(n56553), .B(u_mmu_dtlb_va_addr_q[30]), .Y(n44867) );
  XNOR2X1 U46936 ( .A(n56708), .B(u_mmu_dtlb_va_addr_q[28]), .Y(n44866) );
  NAND2X1 U46937 ( .A(n44867), .B(n44866), .Y(n44873) );
  XNOR2X1 U46938 ( .A(u_mmu_dtlb_va_addr_q[23]), .B(n8320), .Y(n44869) );
  XNOR2X1 U46939 ( .A(u_mmu_dtlb_va_addr_q[25]), .B(n8324), .Y(n44868) );
  NOR2X1 U46940 ( .A(n44869), .B(n44868), .Y(n44871) );
  XNOR2X1 U46941 ( .A(n56367), .B(u_mmu_dtlb_va_addr_q[29]), .Y(n44870) );
  NAND2X1 U46942 ( .A(n44871), .B(n44870), .Y(n44872) );
  NOR2X1 U46943 ( .A(n44873), .B(n44872), .Y(n44883) );
  XOR2X1 U46944 ( .A(n8314), .B(u_mmu_dtlb_va_addr_q[20]), .Y(n44875) );
  XOR2X1 U46945 ( .A(n8308), .B(u_mmu_dtlb_va_addr_q[18]), .Y(n44874) );
  NAND2X1 U46946 ( .A(n44875), .B(n44874), .Y(n44881) );
  XNOR2X1 U46947 ( .A(u_mmu_dtlb_va_addr_q[14]), .B(n8300), .Y(n44877) );
  XNOR2X1 U46948 ( .A(u_mmu_dtlb_va_addr_q[16]), .B(n8304), .Y(n44876) );
  NOR2X1 U46949 ( .A(n44877), .B(n44876), .Y(n44879) );
  XOR2X1 U46950 ( .A(n8310), .B(u_mmu_dtlb_va_addr_q[19]), .Y(n44878) );
  NAND2X1 U46951 ( .A(n44879), .B(n44878), .Y(n44880) );
  NOR2X1 U46952 ( .A(n44881), .B(n44880), .Y(n44882) );
  NAND2X1 U46953 ( .A(n44883), .B(n44882), .Y(n44901) );
  XNOR2X1 U46954 ( .A(u_mmu_dtlb_va_addr_q[26]), .B(n8326), .Y(n44885) );
  XNOR2X1 U46955 ( .A(u_mmu_dtlb_va_addr_q[22]), .B(n8318), .Y(n44884) );
  NOR2X1 U46956 ( .A(n44885), .B(n44884), .Y(n44887) );
  XNOR2X1 U46957 ( .A(n56627), .B(u_mmu_dtlb_va_addr_q[31]), .Y(n44886) );
  NAND2X1 U46958 ( .A(n44887), .B(n44886), .Y(n44888) );
  NOR2X1 U46959 ( .A(n44889), .B(n44888), .Y(n44899) );
  XOR2X1 U46960 ( .A(n8322), .B(u_mmu_dtlb_va_addr_q[24]), .Y(n44891) );
  XOR2X1 U46961 ( .A(n8306), .B(u_mmu_dtlb_va_addr_q[17]), .Y(n44890) );
  NAND2X1 U46962 ( .A(n44891), .B(n44890), .Y(n44897) );
  XNOR2X1 U46963 ( .A(u_mmu_dtlb_va_addr_q[13]), .B(n8298), .Y(n44893) );
  XNOR2X1 U46964 ( .A(u_mmu_dtlb_va_addr_q[15]), .B(n8302), .Y(n44892) );
  NOR2X1 U46965 ( .A(n44893), .B(n44892), .Y(n44895) );
  XOR2X1 U46966 ( .A(n8316), .B(u_mmu_dtlb_va_addr_q[21]), .Y(n44894) );
  NAND2X1 U46967 ( .A(n44895), .B(n44894), .Y(n44896) );
  NOR2X1 U46968 ( .A(n44897), .B(n44896), .Y(n44898) );
  NAND2X1 U46969 ( .A(n44899), .B(n44898), .Y(n44900) );
  NOR2X1 U46970 ( .A(n44901), .B(n44900), .Y(n44944) );
  XNOR2X1 U46971 ( .A(u_mmu_dtlb_va_addr_q[21]), .B(n2549), .Y(n44903) );
  XNOR2X1 U46972 ( .A(u_mmu_dtlb_va_addr_q[13]), .B(n2753), .Y(n44902) );
  NOR2X1 U46973 ( .A(n44903), .B(n44902), .Y(n44905) );
  XOR2X1 U46974 ( .A(n2617), .B(u_mmu_dtlb_va_addr_q[26]), .Y(n44904) );
  NAND2X1 U46975 ( .A(n44905), .B(n44904), .Y(n44906) );
  NOR2X1 U46976 ( .A(n44907), .B(n44906), .Y(n44917) );
  XOR2X1 U46977 ( .A(n2383), .B(u_mmu_dtlb_va_addr_q[20]), .Y(n44909) );
  XOR2X1 U46978 ( .A(n2516), .B(u_mmu_dtlb_va_addr_q[16]), .Y(n44908) );
  NAND2X1 U46979 ( .A(n44909), .B(n44908), .Y(n44915) );
  XNOR2X1 U46980 ( .A(n1872), .B(u_mmu_dtlb_va_addr_q[31]), .Y(n44911) );
  XNOR2X1 U46981 ( .A(u_mmu_dtlb_va_addr_q[29]), .B(n1801), .Y(n44910) );
  NOR2X1 U46982 ( .A(n44911), .B(n44910), .Y(n44913) );
  XOR2X1 U46983 ( .A(n2283), .B(u_mmu_dtlb_va_addr_q[19]), .Y(n44912) );
  NAND2X1 U46984 ( .A(n44913), .B(n44912), .Y(n44914) );
  NOR2X1 U46985 ( .A(n44915), .B(n44914), .Y(n44916) );
  NAND2X1 U46986 ( .A(n44917), .B(n44916), .Y(n44935) );
  XNOR2X1 U46987 ( .A(u_mmu_dtlb_va_addr_q[18]), .B(n2650), .Y(n44919) );
  XNOR2X1 U46988 ( .A(u_mmu_dtlb_va_addr_q[12]), .B(n2683), .Y(n44918) );
  NOR2X1 U46989 ( .A(n44919), .B(n44918), .Y(n44921) );
  XOR2X1 U46990 ( .A(n2850), .B(u_mmu_dtlb_va_addr_q[24]), .Y(n44920) );
  NAND2X1 U46991 ( .A(n44921), .B(n44920), .Y(n44922) );
  NOR2X1 U46992 ( .A(n44923), .B(n44922), .Y(n44933) );
  XOR2X1 U46993 ( .A(n2483), .B(u_mmu_dtlb_va_addr_q[22]), .Y(n44925) );
  XOR2X1 U46994 ( .A(n2451), .B(u_mmu_dtlb_va_addr_q[23]), .Y(n44924) );
  NAND2X1 U46995 ( .A(n44925), .B(n44924), .Y(n44931) );
  XNOR2X1 U46996 ( .A(u_mmu_dtlb_va_addr_q[14]), .B(n1797), .Y(n44927) );
  XNOR2X1 U46997 ( .A(n1871), .B(u_mmu_dtlb_va_addr_q[30]), .Y(n44926) );
  NOR2X1 U46998 ( .A(n44927), .B(n44926), .Y(n44929) );
  XOR2X1 U46999 ( .A(u_mmu_dtlb_va_addr_q[28]), .B(n1870), .Y(n44928) );
  NAND2X1 U47000 ( .A(n44929), .B(n44928), .Y(n44930) );
  NOR2X1 U47001 ( .A(n44931), .B(n44930), .Y(n44932) );
  NAND2X1 U47002 ( .A(n44933), .B(n44932), .Y(n44934) );
  NOR2X1 U47003 ( .A(n44935), .B(n44934), .Y(n44943) );
  OR2X1 U47004 ( .A(u_mmu_store_q[1]), .B(u_mmu_store_q[0]), .Y(n44939) );
  NOR2X1 U47005 ( .A(n58194), .B(n37328), .Y(n44937) );
  NOR2X1 U47006 ( .A(n37327), .B(n58184), .Y(n44936) );
  NAND2X1 U47007 ( .A(n44937), .B(n44936), .Y(n44949) );
  INVX1 U47008 ( .A(n44949), .Y(n57377) );
  NAND2X1 U47009 ( .A(n8574), .B(n57377), .Y(n44938) );
  NOR2X1 U47010 ( .A(n44939), .B(n44938), .Y(n44942) );
  NAND2X1 U47011 ( .A(n37425), .B(n37329), .Y(n44940) );
  NOR2X1 U47012 ( .A(u_mmu_store_q[3]), .B(n44940), .Y(n44941) );
  NAND2X1 U47013 ( .A(n44942), .B(n44941), .Y(n57895) );
  INVX1 U47014 ( .A(n57895), .Y(n57893) );
  MX2X1 U47015 ( .A(n44944), .B(n44943), .S0(n57893), .Y(n44945) );
  NAND2X1 U47016 ( .A(u_mmu_dtlb_valid_q), .B(n44945), .Y(n58166) );
  INVX1 U47017 ( .A(n58166), .Y(n58176) );
  NAND2X1 U47018 ( .A(n58176), .B(n44073), .Y(n58189) );
  NOR2X1 U47019 ( .A(n44946), .B(n58189), .Y(n44948) );
  NAND2X1 U47020 ( .A(n8574), .B(n37425), .Y(n44947) );
  NAND2X1 U47021 ( .A(n44948), .B(n44947), .Y(n58218) );
  NAND2X1 U47022 ( .A(n37329), .B(n37430), .Y(n44952) );
  NOR2X1 U47023 ( .A(u_mmu_store_q[0]), .B(n44949), .Y(n44950) );
  NAND2X1 U47024 ( .A(n44950), .B(n37431), .Y(n44951) );
  NOR2X1 U47025 ( .A(n44952), .B(n44951), .Y(n44953) );
  NAND2X1 U47026 ( .A(n58218), .B(n58216), .Y(n58276) );
  INVX1 U47027 ( .A(n58276), .Y(n58278) );
  NAND2X1 U47028 ( .A(n42559), .B(n58278), .Y(n57427) );
  INVX1 U47029 ( .A(n57427), .Y(n72840) );
  OR2X1 U47030 ( .A(n1848), .B(n1891), .Y(n44956) );
  NAND2X1 U47031 ( .A(n44954), .B(n58164), .Y(n58822) );
  OR2X1 U47032 ( .A(n35945), .B(n58822), .Y(n44955) );
  NOR2X1 U47033 ( .A(n44956), .B(n44955), .Y(n44958) );
  NOR2X1 U47034 ( .A(u_muldiv_div_busy_q), .B(u_muldiv_mult_busy_q), .Y(n44957) );
  NOR2X1 U47035 ( .A(n44958), .B(n44957), .Y(n50046) );
  NOR2X1 U47036 ( .A(n42685), .B(n42723), .Y(n44959) );
  INVX1 U47037 ( .A(n42853), .Y(n48370) );
  NAND2X1 U47038 ( .A(n42667), .B(n42792), .Y(n48585) );
  NAND2X1 U47039 ( .A(n40076), .B(n43017), .Y(n47624) );
  NOR2X1 U47040 ( .A(n24229), .B(n47624), .Y(n44961) );
  INVX1 U47041 ( .A(n42857), .Y(n58130) );
  NAND2X1 U47042 ( .A(n42758), .B(n48370), .Y(n45363) );
  NOR2X1 U47043 ( .A(n24275), .B(n45363), .Y(n44960) );
  NOR2X1 U47044 ( .A(n44961), .B(n44960), .Y(n44962) );
  NAND2X1 U47045 ( .A(n36207), .B(n44962), .Y(n44969) );
  NOR2X1 U47046 ( .A(opcode_opcode_w[17]), .B(n42728), .Y(n44963) );
  NAND2X1 U47047 ( .A(n44963), .B(n42727), .Y(n48560) );
  INVX1 U47048 ( .A(n24239), .Y(n45009) );
  NOR2X1 U47049 ( .A(n39800), .B(n45009), .Y(n44965) );
  NAND2X1 U47050 ( .A(n42667), .B(n42786), .Y(n48607) );
  INVX1 U47051 ( .A(n24125), .Y(n44976) );
  NOR2X1 U47052 ( .A(n47685), .B(n44976), .Y(n44964) );
  NOR2X1 U47053 ( .A(n44965), .B(n44964), .Y(n44967) );
  NAND2X1 U47054 ( .A(n24298), .B(n39137), .Y(n44966) );
  NAND2X1 U47055 ( .A(n44967), .B(n44966), .Y(n44968) );
  NOR2X1 U47056 ( .A(n44969), .B(n44968), .Y(n45002) );
  NAND2X1 U47057 ( .A(n42742), .B(n39669), .Y(n45347) );
  NAND2X1 U47058 ( .A(u_decode_scoreboard_q[21]), .B(n24263), .Y(n57439) );
  NOR2X1 U47059 ( .A(n42200), .B(n57439), .Y(n44972) );
  NOR2X1 U47060 ( .A(opcode_opcode_w[15]), .B(n42726), .Y(n44970) );
  INVX1 U47061 ( .A(n42860), .Y(n47674) );
  INVX1 U47062 ( .A(n42863), .Y(n46341) );
  NOR2X1 U47063 ( .A(n44972), .B(n44971), .Y(n44975) );
  NAND2X1 U47064 ( .A(mem_d_resp_tag_i[2]), .B(n44990), .Y(n45298) );
  INVX1 U47065 ( .A(n45298), .Y(n45162) );
  NAND2X1 U47066 ( .A(n45162), .B(mem_d_resp_tag_i[1]), .Y(n45105) );
  INVX1 U47067 ( .A(n45105), .Y(n73427) );
  NAND2X1 U47068 ( .A(n36009), .B(n73427), .Y(n24188) );
  NOR2X1 U47069 ( .A(n42200), .B(n37434), .Y(n44973) );
  NOR2X1 U47070 ( .A(n24188), .B(n44973), .Y(n44974) );
  NOR2X1 U47071 ( .A(n44975), .B(n44974), .Y(n44981) );
  NOR2X1 U47072 ( .A(n45009), .B(n42782), .Y(n44978) );
  NOR2X1 U47073 ( .A(n44976), .B(n42866), .Y(n44977) );
  NOR2X1 U47074 ( .A(n44978), .B(n44977), .Y(n44979) );
  NOR2X1 U47075 ( .A(n44979), .B(n38802), .Y(n44980) );
  NOR2X1 U47076 ( .A(n44981), .B(n44980), .Y(n44987) );
  INVX1 U47077 ( .A(n45025), .Y(n57515) );
  NAND2X1 U47078 ( .A(n45162), .B(n73556), .Y(n45039) );
  INVX1 U47079 ( .A(n45039), .Y(n73526) );
  NAND2X1 U47080 ( .A(n57515), .B(n73526), .Y(n58156) );
  NAND2X1 U47081 ( .A(u_decode_scoreboard_q[12]), .B(n58156), .Y(n57451) );
  INVX1 U47082 ( .A(n57451), .Y(n44985) );
  NOR2X1 U47083 ( .A(opcode_opcode_w[21]), .B(opcode_opcode_w[20]), .Y(n44982)
         );
  INVX1 U47084 ( .A(n42868), .Y(n46216) );
  NOR2X1 U47085 ( .A(n42729), .B(n42722), .Y(n44983) );
  INVX1 U47086 ( .A(n42871), .Y(n48199) );
  NAND2X1 U47087 ( .A(n38364), .B(n43019), .Y(n45317) );
  NAND2X1 U47088 ( .A(n45245), .B(n45317), .Y(n44984) );
  NAND2X1 U47089 ( .A(n44985), .B(n44984), .Y(n44986) );
  NAND2X1 U47090 ( .A(n44987), .B(n44986), .Y(n45000) );
  NOR2X1 U47091 ( .A(n42687), .B(n42730), .Y(n44988) );
  NAND2X1 U47092 ( .A(n44988), .B(n42722), .Y(n48611) );
  INVX1 U47093 ( .A(n45168), .Y(n58254) );
  INVX1 U47094 ( .A(n46007), .Y(n47422) );
  NOR2X1 U47095 ( .A(n43070), .B(n47422), .Y(n44989) );
  NAND2X1 U47096 ( .A(n44990), .B(mem_d_resp_tag_i[0]), .Y(n45292) );
  NAND2X1 U47097 ( .A(n40841), .B(n57519), .Y(n24170) );
  NAND2X1 U47098 ( .A(u_decode_scoreboard_q[3]), .B(n24170), .Y(n57416) );
  NOR2X1 U47099 ( .A(n44989), .B(n57416), .Y(n44993) );
  NAND2X1 U47100 ( .A(n42793), .B(n42662), .Y(n48595) );
  INVX1 U47101 ( .A(n48595), .Y(n48372) );
  NOR2X1 U47102 ( .A(n43060), .B(n40404), .Y(n44991) );
  NAND2X1 U47103 ( .A(mem_d_resp_tag_i[4]), .B(n44990), .Y(n45299) );
  INVX1 U47104 ( .A(n45299), .Y(n73527) );
  NAND2X1 U47105 ( .A(n40938), .B(n57519), .Y(n24283) );
  NAND2X1 U47106 ( .A(u_decode_scoreboard_q[19]), .B(n24283), .Y(n57423) );
  NOR2X1 U47107 ( .A(n44991), .B(n57423), .Y(n44992) );
  NOR2X1 U47108 ( .A(n44993), .B(n44992), .Y(n44998) );
  NAND2X1 U47109 ( .A(n73427), .B(n40938), .Y(n24247) );
  NAND2X1 U47110 ( .A(u_decode_scoreboard_q[23]), .B(n24247), .Y(n57431) );
  INVX1 U47111 ( .A(n57431), .Y(n44996) );
  INVX1 U47112 ( .A(n46326), .Y(n46183) );
  NOR2X1 U47113 ( .A(n42731), .B(n42725), .Y(n44994) );
  NAND2X1 U47114 ( .A(n49587), .B(n47636), .Y(n44995) );
  NAND2X1 U47115 ( .A(n44996), .B(n44995), .Y(n44997) );
  NAND2X1 U47116 ( .A(n44998), .B(n44997), .Y(n44999) );
  NOR2X1 U47117 ( .A(n45000), .B(n44999), .Y(n45001) );
  NAND2X1 U47118 ( .A(opcode_opcode_w[10]), .B(n54586), .Y(n45046) );
  INVX1 U47119 ( .A(n45046), .Y(n45026) );
  NAND2X1 U47120 ( .A(opcode_opcode_w[7]), .B(n45026), .Y(n58537) );
  INVX1 U47121 ( .A(n58537), .Y(n57472) );
  NAND2X1 U47122 ( .A(n24117), .B(n57472), .Y(n45004) );
  NAND2X1 U47123 ( .A(opcode_opcode_w[11]), .B(n54447), .Y(n45047) );
  INVX1 U47124 ( .A(n45047), .Y(n45024) );
  NAND2X1 U47125 ( .A(opcode_opcode_w[7]), .B(n45024), .Y(n58525) );
  INVX1 U47126 ( .A(n58525), .Y(n57438) );
  NAND2X1 U47127 ( .A(n57438), .B(n24298), .Y(n45003) );
  NAND2X1 U47128 ( .A(n45004), .B(n45003), .Y(n45008) );
  NAND2X1 U47129 ( .A(n45024), .B(n50700), .Y(n58523) );
  INVX1 U47130 ( .A(n58523), .Y(n57541) );
  NAND2X1 U47131 ( .A(n24306), .B(n57541), .Y(n45006) );
  NAND2X1 U47132 ( .A(n45026), .B(n50700), .Y(n58534) );
  INVX1 U47133 ( .A(n58534), .Y(n57456) );
  NAND2X1 U47134 ( .A(n57456), .B(n24125), .Y(n45005) );
  NAND2X1 U47135 ( .A(n45006), .B(n45005), .Y(n45007) );
  NOR2X1 U47136 ( .A(n45008), .B(n45007), .Y(n45017) );
  NAND2X1 U47137 ( .A(opcode_opcode_w[11]), .B(opcode_opcode_w[10]), .Y(n45053) );
  INVX1 U47138 ( .A(n45053), .Y(n45010) );
  NAND2X1 U47139 ( .A(n45010), .B(n50700), .Y(n58529) );
  NOR2X1 U47140 ( .A(n45009), .B(n58529), .Y(n45015) );
  NAND2X1 U47141 ( .A(n45010), .B(opcode_opcode_w[7]), .Y(n57479) );
  INVX1 U47142 ( .A(n57479), .Y(n58531) );
  INVX1 U47143 ( .A(n24229), .Y(n45011) );
  NAND2X1 U47144 ( .A(n58531), .B(n45011), .Y(n45013) );
  NAND2X1 U47145 ( .A(n54586), .B(n54447), .Y(n45052) );
  INVX1 U47146 ( .A(n45052), .Y(n45018) );
  NAND2X1 U47147 ( .A(n45018), .B(opcode_opcode_w[7]), .Y(n57419) );
  INVX1 U47148 ( .A(n57419), .Y(n58527) );
  INVX1 U47149 ( .A(n24275), .Y(n45143) );
  NAND2X1 U47150 ( .A(n58527), .B(n45143), .Y(n45012) );
  NAND2X1 U47151 ( .A(n45013), .B(n45012), .Y(n45014) );
  NOR2X1 U47152 ( .A(n45015), .B(n45014), .Y(n45016) );
  NAND2X1 U47153 ( .A(n45017), .B(n45016), .Y(n45062) );
  INVX1 U47154 ( .A(n58529), .Y(n57493) );
  NAND2X1 U47155 ( .A(u_decode_scoreboard_q[28]), .B(n57493), .Y(n45020) );
  NAND2X1 U47156 ( .A(n45018), .B(n50700), .Y(n57505) );
  INVX1 U47157 ( .A(n57505), .Y(n57535) );
  NAND2X1 U47158 ( .A(u_decode_scoreboard_q[4]), .B(n57535), .Y(n45019) );
  NAND2X1 U47159 ( .A(n45020), .B(n45019), .Y(n45035) );
  INVX1 U47160 ( .A(n45035), .Y(n45023) );
  NAND2X1 U47161 ( .A(n36009), .B(n45052), .Y(n45022) );
  NAND2X1 U47162 ( .A(n57534), .B(n45053), .Y(n45021) );
  NAND2X1 U47163 ( .A(n45022), .B(n45021), .Y(n45092) );
  NOR2X1 U47164 ( .A(n45023), .B(n45092), .Y(n45044) );
  NAND2X1 U47165 ( .A(n36227), .B(n73527), .Y(n57499) );
  NAND2X1 U47166 ( .A(n45024), .B(n57499), .Y(n45028) );
  NAND2X1 U47167 ( .A(n45026), .B(n45025), .Y(n45027) );
  NAND2X1 U47168 ( .A(n45028), .B(n45027), .Y(n45096) );
  NAND2X1 U47169 ( .A(u_decode_scoreboard_q[20]), .B(n57541), .Y(n45030) );
  NAND2X1 U47170 ( .A(n57456), .B(u_decode_scoreboard_q[12]), .Y(n45029) );
  NAND2X1 U47171 ( .A(n45030), .B(n45029), .Y(n45036) );
  NAND2X1 U47172 ( .A(n45096), .B(n45036), .Y(n45042) );
  NAND2X1 U47173 ( .A(n57472), .B(u_decode_scoreboard_q[13]), .Y(n45032) );
  NAND2X1 U47174 ( .A(n57438), .B(u_decode_scoreboard_q[21]), .Y(n45031) );
  NAND2X1 U47175 ( .A(n45032), .B(n45031), .Y(n45045) );
  NAND2X1 U47176 ( .A(n58531), .B(u_decode_scoreboard_q[29]), .Y(n45034) );
  NAND2X1 U47177 ( .A(u_decode_scoreboard_q[5]), .B(n58527), .Y(n45033) );
  NAND2X1 U47178 ( .A(n45034), .B(n45033), .Y(n45051) );
  NOR2X1 U47179 ( .A(n45045), .B(n45051), .Y(n45038) );
  NOR2X1 U47180 ( .A(n45036), .B(n45035), .Y(n45037) );
  NAND2X1 U47181 ( .A(n45038), .B(n45037), .Y(n45040) );
  NAND2X1 U47182 ( .A(n45040), .B(n45039), .Y(n45041) );
  NAND2X1 U47183 ( .A(n45042), .B(n45041), .Y(n45043) );
  NOR2X1 U47184 ( .A(n45044), .B(n45043), .Y(n45060) );
  INVX1 U47185 ( .A(n45045), .Y(n45050) );
  NAND2X1 U47186 ( .A(n40938), .B(n45046), .Y(n45049) );
  NAND2X1 U47187 ( .A(n40937), .B(n45047), .Y(n45048) );
  NAND2X1 U47188 ( .A(n45049), .B(n45048), .Y(n45112) );
  NOR2X1 U47189 ( .A(n45050), .B(n45112), .Y(n45058) );
  INVX1 U47190 ( .A(n45051), .Y(n45056) );
  NAND2X1 U47191 ( .A(n35997), .B(n45052), .Y(n45055) );
  NAND2X1 U47192 ( .A(n40841), .B(n45053), .Y(n45054) );
  NAND2X1 U47193 ( .A(n45055), .B(n45054), .Y(n45115) );
  NOR2X1 U47194 ( .A(n45056), .B(n45115), .Y(n45057) );
  NOR2X1 U47195 ( .A(n45058), .B(n45057), .Y(n45059) );
  NAND2X1 U47196 ( .A(n45060), .B(n45059), .Y(n45061) );
  MX2X1 U47197 ( .A(n45062), .B(n45061), .S0(opcode_opcode_w[9]), .Y(n45124)
         );
  NAND2X1 U47198 ( .A(u_decode_scoreboard_q[11]), .B(n57472), .Y(n45064) );
  NAND2X1 U47199 ( .A(n57438), .B(u_decode_scoreboard_q[19]), .Y(n45063) );
  NAND2X1 U47200 ( .A(n45064), .B(n45063), .Y(n45072) );
  INVX1 U47201 ( .A(n45072), .Y(n45065) );
  NOR2X1 U47202 ( .A(n45065), .B(n45112), .Y(n45081) );
  NAND2X1 U47203 ( .A(u_decode_scoreboard_q[18]), .B(n57541), .Y(n45067) );
  NAND2X1 U47204 ( .A(u_decode_scoreboard_q[10]), .B(n57456), .Y(n45066) );
  NAND2X1 U47205 ( .A(n45067), .B(n45066), .Y(n45073) );
  NAND2X1 U47206 ( .A(n45073), .B(n45096), .Y(n45079) );
  NAND2X1 U47207 ( .A(n58531), .B(u_decode_scoreboard_q[27]), .Y(n45069) );
  NAND2X1 U47208 ( .A(n58527), .B(u_decode_scoreboard_q[3]), .Y(n45068) );
  NAND2X1 U47209 ( .A(n45069), .B(n45068), .Y(n45082) );
  NAND2X1 U47210 ( .A(u_decode_scoreboard_q[26]), .B(n57493), .Y(n45071) );
  NAND2X1 U47211 ( .A(u_decode_scoreboard_q[2]), .B(n57535), .Y(n45070) );
  NAND2X1 U47212 ( .A(n45071), .B(n45070), .Y(n45084) );
  NOR2X1 U47213 ( .A(n45082), .B(n45084), .Y(n45075) );
  NOR2X1 U47214 ( .A(n45073), .B(n45072), .Y(n45074) );
  NAND2X1 U47215 ( .A(n45075), .B(n45074), .Y(n45077) );
  NAND2X1 U47216 ( .A(n45077), .B(n45076), .Y(n45078) );
  NAND2X1 U47217 ( .A(n45079), .B(n45078), .Y(n45080) );
  NOR2X1 U47218 ( .A(n45081), .B(n45080), .Y(n45089) );
  INVX1 U47219 ( .A(n45082), .Y(n45083) );
  NOR2X1 U47220 ( .A(n45083), .B(n45115), .Y(n45087) );
  INVX1 U47221 ( .A(n45084), .Y(n45085) );
  NOR2X1 U47222 ( .A(n45085), .B(n45092), .Y(n45086) );
  NOR2X1 U47223 ( .A(n45087), .B(n45086), .Y(n45088) );
  NAND2X1 U47224 ( .A(n45089), .B(n45088), .Y(n45122) );
  NAND2X1 U47225 ( .A(n57493), .B(u_decode_scoreboard_q[30]), .Y(n45091) );
  NAND2X1 U47226 ( .A(u_decode_scoreboard_q[6]), .B(n57535), .Y(n45090) );
  NAND2X1 U47227 ( .A(n45091), .B(n45090), .Y(n45101) );
  INVX1 U47228 ( .A(n45101), .Y(n45093) );
  NOR2X1 U47229 ( .A(n45093), .B(n45092), .Y(n45110) );
  NAND2X1 U47230 ( .A(u_decode_scoreboard_q[22]), .B(n57541), .Y(n45095) );
  NAND2X1 U47231 ( .A(n57456), .B(u_decode_scoreboard_q[14]), .Y(n45094) );
  NAND2X1 U47232 ( .A(n45095), .B(n45094), .Y(n45102) );
  NAND2X1 U47233 ( .A(n45102), .B(n45096), .Y(n45108) );
  NAND2X1 U47234 ( .A(n57472), .B(u_decode_scoreboard_q[15]), .Y(n45098) );
  NAND2X1 U47235 ( .A(n57438), .B(u_decode_scoreboard_q[23]), .Y(n45097) );
  NAND2X1 U47236 ( .A(n45098), .B(n45097), .Y(n45111) );
  NAND2X1 U47237 ( .A(u_decode_scoreboard_q[31]), .B(n58531), .Y(n45100) );
  NAND2X1 U47238 ( .A(u_decode_scoreboard_q[7]), .B(n58527), .Y(n45099) );
  NAND2X1 U47239 ( .A(n45100), .B(n45099), .Y(n45114) );
  NOR2X1 U47240 ( .A(n45111), .B(n45114), .Y(n45104) );
  NOR2X1 U47241 ( .A(n45102), .B(n45101), .Y(n45103) );
  NAND2X1 U47242 ( .A(n45104), .B(n45103), .Y(n45106) );
  NAND2X1 U47243 ( .A(n45106), .B(n45105), .Y(n45107) );
  NAND2X1 U47244 ( .A(n45108), .B(n45107), .Y(n45109) );
  NOR2X1 U47245 ( .A(n45110), .B(n45109), .Y(n45120) );
  INVX1 U47246 ( .A(n45111), .Y(n45113) );
  NOR2X1 U47247 ( .A(n45113), .B(n45112), .Y(n45118) );
  INVX1 U47248 ( .A(n45114), .Y(n45116) );
  NOR2X1 U47249 ( .A(n45116), .B(n45115), .Y(n45117) );
  NOR2X1 U47250 ( .A(n45118), .B(n45117), .Y(n45119) );
  NAND2X1 U47251 ( .A(n45120), .B(n45119), .Y(n45121) );
  MX2X1 U47252 ( .A(n45122), .B(n45121), .S0(opcode_opcode_w[9]), .Y(n45123)
         );
  MX2X1 U47253 ( .A(n45124), .B(n45123), .S0(opcode_opcode_w[8]), .Y(n45125)
         );
  OR2X1 U47254 ( .A(n36228), .B(n45125), .Y(n45126) );
  NOR2X1 U47255 ( .A(n36191), .B(n45126), .Y(n45129) );
  OR2X1 U47256 ( .A(n35999), .B(n36175), .Y(n45127) );
  NOR2X1 U47257 ( .A(n35970), .B(n45127), .Y(n45128) );
  NAND2X1 U47258 ( .A(n45129), .B(n45128), .Y(n45154) );
  INVX1 U47259 ( .A(n49594), .Y(n49674) );
  NOR2X1 U47260 ( .A(n43051), .B(n40519), .Y(n45130) );
  NAND2X1 U47261 ( .A(n35997), .B(n73526), .Y(n24203) );
  NAND2X1 U47262 ( .A(u_decode_scoreboard_q[29]), .B(n24203), .Y(n57467) );
  NOR2X1 U47263 ( .A(n45130), .B(n57467), .Y(n45138) );
  NAND2X1 U47264 ( .A(n40937), .B(n73427), .Y(n24316) );
  NAND2X1 U47265 ( .A(u_decode_scoreboard_q[15]), .B(n24316), .Y(n57462) );
  INVX1 U47266 ( .A(n57462), .Y(n45132) );
  NAND2X1 U47267 ( .A(n42682), .B(n47625), .Y(n45131) );
  NAND2X1 U47268 ( .A(n45132), .B(n45131), .Y(n45136) );
  NAND2X1 U47269 ( .A(n57515), .B(n73427), .Y(n24328) );
  NAND2X1 U47270 ( .A(u_decode_scoreboard_q[14]), .B(n24328), .Y(n57457) );
  INVX1 U47271 ( .A(n57457), .Y(n45134) );
  NAND2X1 U47272 ( .A(n47674), .B(n43019), .Y(n45324) );
  NAND2X1 U47273 ( .A(n45244), .B(n45324), .Y(n45133) );
  NAND2X1 U47274 ( .A(n45134), .B(n45133), .Y(n45135) );
  NAND2X1 U47275 ( .A(n45136), .B(n45135), .Y(n45137) );
  NOR2X1 U47276 ( .A(n45138), .B(n45137), .Y(n45152) );
  NOR2X1 U47277 ( .A(n43071), .B(n45614), .Y(n45139) );
  NAND2X1 U47278 ( .A(n35997), .B(n57519), .Y(n24217) );
  NAND2X1 U47279 ( .A(u_decode_scoreboard_q[27]), .B(n24217), .Y(n57478) );
  NOR2X1 U47280 ( .A(n45139), .B(n57478), .Y(n45150) );
  INVX1 U47281 ( .A(n58469), .Y(n51983) );
  INVX1 U47282 ( .A(n24298), .Y(n45140) );
  NOR2X1 U47283 ( .A(n45140), .B(n40509), .Y(n45142) );
  NOR2X1 U47284 ( .A(n24229), .B(n42782), .Y(n45141) );
  NOR2X1 U47285 ( .A(n45142), .B(n45141), .Y(n45145) );
  NAND2X1 U47286 ( .A(n42771), .B(n45143), .Y(n45144) );
  NAND2X1 U47287 ( .A(n45145), .B(n45144), .Y(n45146) );
  NAND2X1 U47288 ( .A(n38537), .B(n45146), .Y(n45148) );
  NAND2X1 U47289 ( .A(n40937), .B(n73526), .Y(n24336) );
  NAND2X1 U47290 ( .A(u_decode_scoreboard_q[13]), .B(n24336), .Y(n57473) );
  NAND2X1 U47291 ( .A(n42743), .B(n42673), .Y(n45350) );
  NAND2X1 U47292 ( .A(n45148), .B(n45147), .Y(n45149) );
  NOR2X1 U47293 ( .A(n45150), .B(n45149), .Y(n45151) );
  NAND2X1 U47294 ( .A(n45152), .B(n45151), .Y(n45153) );
  OR2X1 U47295 ( .A(n50046), .B(n50045), .Y(n45156) );
  NAND2X1 U47296 ( .A(u_decode_valid_q), .B(n8696), .Y(n45155) );
  NOR2X1 U47297 ( .A(n45156), .B(n45155), .Y(n50530) );
  NAND2X1 U47298 ( .A(n72840), .B(n50530), .Y(n57362) );
  INVX1 U47299 ( .A(n57362), .Y(n57351) );
  NAND2X1 U47300 ( .A(n58183), .B(n37448), .Y(n45157) );
  NOR2X1 U47301 ( .A(n44257), .B(n440), .Y(n45158) );
  NAND2X1 U47302 ( .A(n44073), .B(n58166), .Y(n52001) );
  NAND2X1 U47303 ( .A(n45158), .B(n52001), .Y(n45159) );
  NAND2X1 U47304 ( .A(n45160), .B(n57377), .Y(n45161) );
  NAND2X1 U47305 ( .A(n42441), .B(n45161), .Y(n28934) );
  INVX1 U47306 ( .A(n42872), .Y(n54897) );
  XNOR2X1 U47307 ( .A(opcode_opcode_w[22]), .B(n45162), .Y(n45173) );
  INVX1 U47308 ( .A(n45173), .Y(n45165) );
  NAND2X1 U47309 ( .A(opcode_opcode_w[20]), .B(n73557), .Y(n45174) );
  XNOR2X1 U47310 ( .A(opcode_opcode_w[23]), .B(n45163), .Y(n45175) );
  NAND2X1 U47311 ( .A(n45174), .B(n45175), .Y(n45164) );
  NOR2X1 U47312 ( .A(opcode_opcode_w[21]), .B(n73556), .Y(n45167) );
  NOR2X1 U47313 ( .A(opcode_opcode_w[20]), .B(n45292), .Y(n45166) );
  NAND2X1 U47314 ( .A(n35922), .B(n57534), .Y(n45293) );
  NOR2X1 U47315 ( .A(n45168), .B(n40508), .Y(n45169) );
  NAND2X1 U47316 ( .A(n45169), .B(n2942), .Y(n45170) );
  NOR2X1 U47317 ( .A(n42231), .B(n45170), .Y(n45171) );
  XNOR2X1 U47318 ( .A(writeback_exec_idx_w[4]), .B(opcode_opcode_w[24]), .Y(
        n45276) );
  XNOR2X1 U47319 ( .A(opcode_opcode_w[23]), .B(writeback_exec_idx_w[3]), .Y(
        n45534) );
  NAND2X1 U47320 ( .A(n45171), .B(n42705), .Y(n45180) );
  NOR2X1 U47321 ( .A(n40579), .B(n38637), .Y(n45172) );
  NAND2X1 U47322 ( .A(n45172), .B(n45534), .Y(n45181) );
  INVX1 U47323 ( .A(n45277), .Y(n45446) );
  NAND2X1 U47324 ( .A(n45520), .B(n39501), .Y(n45176) );
  NOR2X1 U47325 ( .A(n42230), .B(n46009), .Y(n45178) );
  INVX1 U47326 ( .A(n58820), .Y(n58458) );
  NOR2X1 U47327 ( .A(n57608), .B(n37074), .Y(n45177) );
  NAND2X1 U47328 ( .A(n45178), .B(n45177), .Y(n45179) );
  NAND2X1 U47329 ( .A(n45180), .B(n45179), .Y(n60948) );
  INVX1 U47330 ( .A(n60948), .Y(n61190) );
  NAND2X1 U47331 ( .A(n45276), .B(n45533), .Y(n45255) );
  NOR2X1 U47332 ( .A(n45277), .B(n45255), .Y(n45182) );
  NOR2X1 U47333 ( .A(n46009), .B(n45182), .Y(n45184) );
  NAND2X1 U47334 ( .A(n46216), .B(n58254), .Y(n46577) );
  NOR2X1 U47335 ( .A(n46577), .B(n37067), .Y(n45183) );
  NAND2X1 U47336 ( .A(n45184), .B(n45183), .Y(n45191) );
  NAND2X1 U47337 ( .A(n46054), .B(n58254), .Y(n45185) );
  NAND2X1 U47338 ( .A(n42771), .B(n58254), .Y(n45186) );
  NOR2X1 U47339 ( .A(n42230), .B(n45187), .Y(n45189) );
  NAND2X1 U47340 ( .A(n45189), .B(n40152), .Y(n45190) );
  NAND2X1 U47341 ( .A(n45191), .B(n45190), .Y(n60949) );
  INVX1 U47342 ( .A(n60949), .Y(n61189) );
  INVX1 U47343 ( .A(n46366), .Y(n61188) );
  NOR2X1 U47344 ( .A(n45193), .B(n45192), .Y(n45198) );
  NAND2X1 U47345 ( .A(n2943), .B(n40523), .Y(n45194) );
  NOR2X1 U47346 ( .A(n40508), .B(n45194), .Y(n45195) );
  NOR2X1 U47347 ( .A(n45196), .B(n45195), .Y(n45197) );
  NAND2X1 U47348 ( .A(n45198), .B(n45197), .Y(n45218) );
  NAND2X1 U47349 ( .A(opcode_opcode_w[23]), .B(opcode_opcode_w[24]), .Y(n45199) );
  NOR2X1 U47350 ( .A(n36795), .B(n42783), .Y(n45202) );
  NAND2X1 U47351 ( .A(n42749), .B(n42760), .Y(n45200) );
  NOR2X1 U47352 ( .A(n36797), .B(n45200), .Y(n45201) );
  NOR2X1 U47353 ( .A(n45202), .B(n45201), .Y(n45203) );
  NOR2X1 U47354 ( .A(n45203), .B(n38823), .Y(n45206) );
  NAND2X1 U47355 ( .A(n2944), .B(n38947), .Y(n45204) );
  NOR2X1 U47356 ( .A(n40510), .B(n45204), .Y(n45205) );
  NOR2X1 U47357 ( .A(n45206), .B(n45205), .Y(n45216) );
  NOR2X1 U47358 ( .A(n40454), .B(n42747), .Y(n45207) );
  NAND2X1 U47359 ( .A(n45207), .B(n2925), .Y(n45208) );
  NOR2X1 U47360 ( .A(n42881), .B(n45208), .Y(n45214) );
  NAND2X1 U47361 ( .A(n45209), .B(n38947), .Y(n45212) );
  NAND2X1 U47362 ( .A(n42516), .B(n45210), .Y(n45211) );
  NAND2X1 U47363 ( .A(n45212), .B(n45211), .Y(n45213) );
  NOR2X1 U47364 ( .A(n45214), .B(n45213), .Y(n45215) );
  NAND2X1 U47365 ( .A(n45216), .B(n45215), .Y(n45217) );
  NAND2X1 U47366 ( .A(n40453), .B(n36599), .Y(n45220) );
  NAND2X1 U47367 ( .A(n2923), .B(n39115), .Y(n45219) );
  NOR2X1 U47368 ( .A(n45220), .B(n45219), .Y(n45221) );
  NAND2X1 U47369 ( .A(n45221), .B(n46054), .Y(n45227) );
  NAND2X1 U47370 ( .A(n36599), .B(n42749), .Y(n45222) );
  NOR2X1 U47371 ( .A(n39116), .B(n45222), .Y(n45225) );
  NAND2X1 U47372 ( .A(n40453), .B(n42760), .Y(n45223) );
  NOR2X1 U47373 ( .A(n36796), .B(n45223), .Y(n45224) );
  NAND2X1 U47374 ( .A(n45225), .B(n45224), .Y(n45226) );
  NAND2X1 U47375 ( .A(n45227), .B(n45226), .Y(n45228) );
  NOR2X1 U47376 ( .A(n45229), .B(n45228), .Y(n45239) );
  NOR2X1 U47377 ( .A(n1799), .B(n39116), .Y(n45231) );
  NOR2X1 U47378 ( .A(n2945), .B(n39115), .Y(n45230) );
  NOR2X1 U47379 ( .A(n45231), .B(n45230), .Y(n45233) );
  NOR2X1 U47380 ( .A(n38919), .B(n42762), .Y(n45232) );
  NAND2X1 U47381 ( .A(n45233), .B(n45232), .Y(n45234) );
  NOR2X1 U47382 ( .A(n40507), .B(n45234), .Y(n45237) );
  NAND2X1 U47383 ( .A(n2941), .B(n42516), .Y(n45235) );
  NOR2X1 U47384 ( .A(n40511), .B(n45235), .Y(n45236) );
  NOR2X1 U47385 ( .A(n45237), .B(n45236), .Y(n45238) );
  NAND2X1 U47386 ( .A(n45239), .B(n45238), .Y(n45249) );
  NOR2X1 U47387 ( .A(n42747), .B(n42760), .Y(n45240) );
  NAND2X1 U47388 ( .A(n45240), .B(n2933), .Y(n45241) );
  NOR2X1 U47389 ( .A(n42875), .B(n45241), .Y(n45243) );
  NOR2X1 U47390 ( .A(n36843), .B(n45244), .Y(n45247) );
  NAND2X1 U47391 ( .A(n40523), .B(n46049), .Y(n45245) );
  NAND2X1 U47392 ( .A(n61188), .B(n61187), .Y(n63821) );
  NAND2X1 U47393 ( .A(n58458), .B(n46216), .Y(n45250) );
  NOR2X1 U47394 ( .A(n36818), .B(n45250), .Y(n45253) );
  NAND2X1 U47395 ( .A(n58458), .B(n46341), .Y(n45251) );
  NOR2X1 U47396 ( .A(n36819), .B(n45251), .Y(n45252) );
  NOR2X1 U47397 ( .A(n45253), .B(n45252), .Y(n45254) );
  NOR2X1 U47398 ( .A(n42231), .B(n45254), .Y(n45256) );
  NAND2X1 U47399 ( .A(n50802), .B(n50720), .Y(n50792) );
  NAND2X1 U47400 ( .A(n50824), .B(n39766), .Y(n45262) );
  NOR2X1 U47401 ( .A(n50792), .B(n45262), .Y(n45258) );
  OR2X1 U47402 ( .A(writeback_exec_idx_w[4]), .B(opcode_opcode_w[24]), .Y(
        n45257) );
  NOR2X1 U47403 ( .A(n45258), .B(n45257), .Y(n45530) );
  NOR2X1 U47404 ( .A(n42498), .B(n45530), .Y(n45259) );
  NAND2X1 U47405 ( .A(n45267), .B(n45266), .Y(n45531) );
  NOR2X1 U47406 ( .A(n45259), .B(n45531), .Y(n45260) );
  NAND2X1 U47407 ( .A(n45534), .B(n45533), .Y(n45271) );
  NOR2X1 U47408 ( .A(writeback_exec_idx_w[1]), .B(writeback_exec_idx_w[2]), 
        .Y(n45263) );
  NAND2X1 U47409 ( .A(n45264), .B(n45263), .Y(n45265) );
  NAND2X1 U47410 ( .A(n45266), .B(n45265), .Y(n45536) );
  XNOR2X1 U47411 ( .A(writeback_exec_idx_w[4]), .B(n42748), .Y(n45268) );
  NAND2X1 U47412 ( .A(n45268), .B(n45267), .Y(n45537) );
  INVX1 U47413 ( .A(n45537), .Y(n45269) );
  NAND2X1 U47414 ( .A(n36620), .B(n45269), .Y(n45270) );
  NOR2X1 U47415 ( .A(n45271), .B(n45270), .Y(n45274) );
  INVX1 U47416 ( .A(mem_d_data_rd_i[31]), .Y(n45272) );
  NAND2X1 U47417 ( .A(n40935), .B(n45272), .Y(n45273) );
  NOR2X1 U47418 ( .A(n45274), .B(n43279), .Y(n45275) );
  NAND2X1 U47419 ( .A(n45275), .B(n46024), .Y(n45290) );
  NAND2X1 U47420 ( .A(n45172), .B(n45534), .Y(n45277) );
  NOR2X1 U47421 ( .A(n45181), .B(n38807), .Y(n45278) );
  NOR2X1 U47422 ( .A(n42231), .B(n45278), .Y(n45288) );
  NAND2X1 U47423 ( .A(n2940), .B(n51983), .Y(n45279) );
  NOR2X1 U47424 ( .A(n40507), .B(n45279), .Y(n45282) );
  NAND2X1 U47425 ( .A(n51983), .B(n42770), .Y(n45280) );
  NOR2X1 U47426 ( .A(n36832), .B(n45280), .Y(n45281) );
  NOR2X1 U47427 ( .A(n45282), .B(n45281), .Y(n45286) );
  NOR2X1 U47428 ( .A(n45284), .B(n45283), .Y(n45285) );
  NAND2X1 U47429 ( .A(n45286), .B(n45285), .Y(n45287) );
  NAND2X1 U47430 ( .A(n45288), .B(n45287), .Y(n45289) );
  OR2X1 U47431 ( .A(n63823), .B(n45291), .Y(n72348) );
  XOR2X1 U47432 ( .A(n42723), .B(mem_d_resp_tag_i[1]), .Y(n45296) );
  MX2X1 U47433 ( .A(n45292), .B(mem_d_resp_tag_i[0]), .S0(n42729), .Y(n45294)
         );
  NAND2X1 U47434 ( .A(n45294), .B(n45293), .Y(n45295) );
  NOR2X1 U47435 ( .A(n45296), .B(n45295), .Y(n45311) );
  XNOR2X1 U47436 ( .A(n45297), .B(n42668), .Y(n45303) );
  XOR2X1 U47437 ( .A(n45298), .B(n42686), .Y(n45301) );
  XOR2X1 U47438 ( .A(n45299), .B(n42794), .Y(n45300) );
  NAND2X1 U47439 ( .A(n45301), .B(n45300), .Y(n45302) );
  NOR2X1 U47440 ( .A(n45303), .B(n45302), .Y(n45310) );
  XNOR2X1 U47441 ( .A(writeback_exec_idx_w[4]), .B(n42792), .Y(n45307) );
  NAND2X1 U47442 ( .A(n42787), .B(n39766), .Y(n45304) );
  NOR2X1 U47443 ( .A(n50792), .B(n45304), .Y(n45305) );
  NAND2X1 U47444 ( .A(n45305), .B(n50824), .Y(n45306) );
  NAND2X1 U47445 ( .A(n45307), .B(n45306), .Y(n48105) );
  NOR2X1 U47446 ( .A(n43279), .B(n43455), .Y(n45309) );
  INVX1 U47447 ( .A(writeback_exec_value_w[31]), .Y(n57234) );
  NAND2X1 U47448 ( .A(n39210), .B(n39612), .Y(n49806) );
  NOR2X1 U47449 ( .A(n43282), .B(n43023), .Y(n45308) );
  NAND2X1 U47450 ( .A(n45311), .B(n45310), .Y(n62905) );
  NAND2X1 U47451 ( .A(n42377), .B(n39612), .Y(n45314) );
  NAND2X1 U47452 ( .A(n62905), .B(n45314), .Y(n64082) );
  INVX1 U47453 ( .A(n64082), .Y(n59145) );
  NAND2X1 U47454 ( .A(n2945), .B(n43363), .Y(n45316) );
  NAND2X1 U47455 ( .A(n38413), .B(n2920), .Y(n45315) );
  NAND2X1 U47456 ( .A(n45316), .B(n45315), .Y(n45321) );
  NAND2X1 U47457 ( .A(n38402), .B(n2927), .Y(n45319) );
  NAND2X1 U47458 ( .A(n43027), .B(n2935), .Y(n45318) );
  NAND2X1 U47459 ( .A(n45319), .B(n45318), .Y(n45320) );
  NOR2X1 U47460 ( .A(n45321), .B(n45320), .Y(n45330) );
  NAND2X1 U47461 ( .A(n2917), .B(n43031), .Y(n45323) );
  NAND2X1 U47462 ( .A(n43032), .B(n2922), .Y(n45322) );
  NAND2X1 U47463 ( .A(n45323), .B(n45322), .Y(n45328) );
  NAND2X1 U47464 ( .A(n43036), .B(n2937), .Y(n45326) );
  NAND2X1 U47465 ( .A(n43351), .B(n2929), .Y(n45325) );
  NAND2X1 U47466 ( .A(n45326), .B(n45325), .Y(n45327) );
  NOR2X1 U47467 ( .A(n45328), .B(n45327), .Y(n45329) );
  NAND2X1 U47468 ( .A(n45330), .B(n45329), .Y(n45346) );
  INVX1 U47469 ( .A(n42879), .Y(n48205) );
  NAND2X1 U47470 ( .A(n43355), .B(n2933), .Y(n45332) );
  NAND2X1 U47471 ( .A(n2931), .B(n43040), .Y(n45331) );
  NAND2X1 U47472 ( .A(n45332), .B(n45331), .Y(n45336) );
  NAND2X1 U47473 ( .A(n1792), .B(n39805), .Y(n45334) );
  NAND2X1 U47474 ( .A(n39584), .B(n40018), .Y(n57609) );
  NAND2X1 U47475 ( .A(n43042), .B(n2939), .Y(n45333) );
  NAND2X1 U47476 ( .A(n45334), .B(n45333), .Y(n45335) );
  NOR2X1 U47477 ( .A(n45336), .B(n45335), .Y(n45344) );
  NAND2X1 U47478 ( .A(n38390), .B(n2943), .Y(n45338) );
  NAND2X1 U47479 ( .A(n43345), .B(n2918), .Y(n45337) );
  NAND2X1 U47480 ( .A(n45338), .B(n45337), .Y(n45342) );
  NAND2X1 U47481 ( .A(n43338), .B(n2925), .Y(n45340) );
  NAND2X1 U47482 ( .A(n43365), .B(n2941), .Y(n45339) );
  NAND2X1 U47483 ( .A(n45340), .B(n45339), .Y(n45341) );
  NOR2X1 U47484 ( .A(n45342), .B(n45341), .Y(n45343) );
  NAND2X1 U47485 ( .A(n45344), .B(n45343), .Y(n45345) );
  NOR2X1 U47486 ( .A(n45346), .B(n45345), .Y(n45379) );
  NAND2X1 U47487 ( .A(n43044), .B(n2938), .Y(n45349) );
  NAND2X1 U47488 ( .A(n43047), .B(n2944), .Y(n45348) );
  NAND2X1 U47489 ( .A(n45349), .B(n45348), .Y(n45354) );
  INVX1 U47490 ( .A(n45350), .Y(n49841) );
  NAND2X1 U47491 ( .A(n43049), .B(n2936), .Y(n45352) );
  NAND2X1 U47492 ( .A(n43051), .B(n2921), .Y(n45351) );
  NAND2X1 U47493 ( .A(n45352), .B(n45351), .Y(n45353) );
  NOR2X1 U47494 ( .A(n45354), .B(n45353), .Y(n45360) );
  NOR2X1 U47495 ( .A(n36796), .B(n43370), .Y(n45358) );
  NAND2X1 U47496 ( .A(n42735), .B(n43018), .Y(n57625) );
  NAND2X1 U47497 ( .A(n43054), .B(n2923), .Y(n45356) );
  NAND2X1 U47498 ( .A(n1799), .B(n43058), .Y(n45355) );
  NAND2X1 U47499 ( .A(n45356), .B(n45355), .Y(n45357) );
  NOR2X1 U47500 ( .A(n45358), .B(n45357), .Y(n45359) );
  NAND2X1 U47501 ( .A(n45360), .B(n45359), .Y(n45377) );
  NAND2X1 U47502 ( .A(n43060), .B(n2942), .Y(n45362) );
  NAND2X1 U47503 ( .A(n2940), .B(n39139), .Y(n45361) );
  NAND2X1 U47504 ( .A(n45362), .B(n45361), .Y(n45367) );
  NAND2X1 U47505 ( .A(n40076), .B(n43019), .Y(n57604) );
  NAND2X1 U47506 ( .A(n43063), .B(n2932), .Y(n45365) );
  NAND2X1 U47507 ( .A(n2924), .B(n43068), .Y(n45364) );
  NAND2X1 U47508 ( .A(n45365), .B(n45364), .Y(n45366) );
  NOR2X1 U47509 ( .A(n45367), .B(n45366), .Y(n45375) );
  NAND2X1 U47510 ( .A(n42742), .B(n42757), .Y(n47637) );
  NAND2X1 U47511 ( .A(n43372), .B(n2928), .Y(n45369) );
  NAND2X1 U47512 ( .A(n40448), .B(n43019), .Y(n47621) );
  NAND2X1 U47513 ( .A(n43350), .B(n2934), .Y(n45368) );
  NAND2X1 U47514 ( .A(n45369), .B(n45368), .Y(n45373) );
  NAND2X1 U47515 ( .A(n43070), .B(n2926), .Y(n45371) );
  NAND2X1 U47516 ( .A(n43071), .B(n2919), .Y(n45370) );
  NAND2X1 U47517 ( .A(n45371), .B(n45370), .Y(n45372) );
  NOR2X1 U47518 ( .A(n45373), .B(n45372), .Y(n45374) );
  NAND2X1 U47519 ( .A(n45375), .B(n45374), .Y(n45376) );
  NOR2X1 U47520 ( .A(n45377), .B(n45376), .Y(n45378) );
  NAND2X1 U47521 ( .A(n45379), .B(n45378), .Y(n45380) );
  NAND2X1 U47522 ( .A(n43611), .B(n44054), .Y(n49885) );
  INVX1 U47523 ( .A(n49885), .Y(n58158) );
  INVX1 U47524 ( .A(mem_d_data_rd_i[29]), .Y(n45381) );
  NAND2X1 U47525 ( .A(n40935), .B(n45381), .Y(n45382) );
  NOR2X1 U47526 ( .A(n43455), .B(n43223), .Y(n45384) );
  NOR2X1 U47527 ( .A(n43022), .B(n43226), .Y(n45383) );
  NAND2X1 U47528 ( .A(n3011), .B(n43363), .Y(n45386) );
  NAND2X1 U47529 ( .A(n2986), .B(n38409), .Y(n45385) );
  NAND2X1 U47530 ( .A(n45386), .B(n45385), .Y(n45390) );
  NAND2X1 U47531 ( .A(n2993), .B(n38401), .Y(n45388) );
  NAND2X1 U47532 ( .A(n3001), .B(n43027), .Y(n45387) );
  NAND2X1 U47533 ( .A(n45388), .B(n45387), .Y(n45389) );
  NOR2X1 U47534 ( .A(n45390), .B(n45389), .Y(n45398) );
  NAND2X1 U47535 ( .A(n2983), .B(n43031), .Y(n45392) );
  NAND2X1 U47536 ( .A(n2988), .B(n43032), .Y(n45391) );
  NAND2X1 U47537 ( .A(n45392), .B(n45391), .Y(n45396) );
  NAND2X1 U47538 ( .A(n3003), .B(n43036), .Y(n45394) );
  NAND2X1 U47539 ( .A(n2995), .B(n43351), .Y(n45393) );
  NAND2X1 U47540 ( .A(n45394), .B(n45393), .Y(n45395) );
  NOR2X1 U47541 ( .A(n45396), .B(n45395), .Y(n45397) );
  NAND2X1 U47542 ( .A(n45398), .B(n45397), .Y(n45414) );
  NAND2X1 U47543 ( .A(n2999), .B(n43354), .Y(n45400) );
  NAND2X1 U47544 ( .A(n2997), .B(n43040), .Y(n45399) );
  NAND2X1 U47545 ( .A(n45400), .B(n45399), .Y(n45404) );
  NAND2X1 U47546 ( .A(n1800), .B(n39803), .Y(n45402) );
  NAND2X1 U47547 ( .A(n3005), .B(n43042), .Y(n45401) );
  NAND2X1 U47548 ( .A(n45402), .B(n45401), .Y(n45403) );
  NOR2X1 U47549 ( .A(n45404), .B(n45403), .Y(n45412) );
  NAND2X1 U47550 ( .A(n3009), .B(n38389), .Y(n45406) );
  NAND2X1 U47551 ( .A(n2984), .B(n43345), .Y(n45405) );
  NAND2X1 U47552 ( .A(n45406), .B(n45405), .Y(n45410) );
  NAND2X1 U47553 ( .A(n2991), .B(n43338), .Y(n45408) );
  NAND2X1 U47554 ( .A(n3007), .B(n43365), .Y(n45407) );
  NAND2X1 U47555 ( .A(n45408), .B(n45407), .Y(n45409) );
  NOR2X1 U47556 ( .A(n45410), .B(n45409), .Y(n45411) );
  NAND2X1 U47557 ( .A(n45412), .B(n45411), .Y(n45413) );
  NOR2X1 U47558 ( .A(n45414), .B(n45413), .Y(n45444) );
  NAND2X1 U47559 ( .A(n3004), .B(n43044), .Y(n45416) );
  NAND2X1 U47560 ( .A(n3010), .B(n43047), .Y(n45415) );
  NAND2X1 U47561 ( .A(n45416), .B(n45415), .Y(n45420) );
  NAND2X1 U47562 ( .A(n3002), .B(n43049), .Y(n45418) );
  NAND2X1 U47563 ( .A(n2987), .B(n43051), .Y(n45417) );
  NAND2X1 U47564 ( .A(n45418), .B(n45417), .Y(n45419) );
  NOR2X1 U47565 ( .A(n45420), .B(n45419), .Y(n45426) );
  NOR2X1 U47566 ( .A(n43371), .B(n37324), .Y(n45424) );
  NAND2X1 U47567 ( .A(n2989), .B(n43054), .Y(n45422) );
  NAND2X1 U47568 ( .A(n1802), .B(n43058), .Y(n45421) );
  NAND2X1 U47569 ( .A(n45422), .B(n45421), .Y(n45423) );
  NOR2X1 U47570 ( .A(n45424), .B(n45423), .Y(n45425) );
  NAND2X1 U47571 ( .A(n45426), .B(n45425), .Y(n45442) );
  NAND2X1 U47572 ( .A(n3008), .B(n43060), .Y(n45428) );
  NAND2X1 U47573 ( .A(n3006), .B(n39135), .Y(n45427) );
  NAND2X1 U47574 ( .A(n45428), .B(n45427), .Y(n45432) );
  NAND2X1 U47575 ( .A(n2998), .B(n43063), .Y(n45430) );
  NAND2X1 U47576 ( .A(n2990), .B(n43068), .Y(n45429) );
  NAND2X1 U47577 ( .A(n45430), .B(n45429), .Y(n45431) );
  NOR2X1 U47578 ( .A(n45432), .B(n45431), .Y(n45440) );
  NAND2X1 U47579 ( .A(n2994), .B(n43372), .Y(n45434) );
  NAND2X1 U47580 ( .A(n3000), .B(n43349), .Y(n45433) );
  NAND2X1 U47581 ( .A(n45434), .B(n45433), .Y(n45438) );
  NAND2X1 U47582 ( .A(n2992), .B(n43070), .Y(n45436) );
  NAND2X1 U47583 ( .A(n2985), .B(n43071), .Y(n45435) );
  NAND2X1 U47584 ( .A(n45436), .B(n45435), .Y(n45437) );
  NOR2X1 U47585 ( .A(n45438), .B(n45437), .Y(n45439) );
  NAND2X1 U47586 ( .A(n45440), .B(n45439), .Y(n45441) );
  NOR2X1 U47587 ( .A(n45442), .B(n45441), .Y(n45443) );
  NAND2X1 U47588 ( .A(n45444), .B(n45443), .Y(n45445) );
  INVX1 U47589 ( .A(n46372), .Y(n46979) );
  NAND2X1 U47590 ( .A(n2990), .B(n46979), .Y(n45448) );
  NAND2X1 U47591 ( .A(n45176), .B(n45710), .Y(n45447) );
  NOR2X1 U47592 ( .A(n45448), .B(n45447), .Y(n45451) );
  INVX1 U47593 ( .A(n57608), .Y(n46741) );
  NAND2X1 U47594 ( .A(n3005), .B(n46741), .Y(n45449) );
  NOR2X1 U47595 ( .A(n45451), .B(n45450), .Y(n45455) );
  NOR2X1 U47596 ( .A(n46236), .B(n37029), .Y(n45452) );
  NAND2X1 U47597 ( .A(n45453), .B(n45452), .Y(n45454) );
  NAND2X1 U47598 ( .A(n45455), .B(n45454), .Y(n45463) );
  NOR2X1 U47599 ( .A(n46009), .B(n38846), .Y(n45457) );
  NOR2X1 U47600 ( .A(n46570), .B(n37034), .Y(n45456) );
  NAND2X1 U47601 ( .A(n45457), .B(n45456), .Y(n45461) );
  INVX1 U47602 ( .A(n46014), .Y(n46235) );
  NOR2X1 U47603 ( .A(n45521), .B(n46024), .Y(n45459) );
  NOR2X1 U47604 ( .A(n46007), .B(n37037), .Y(n45458) );
  NAND2X1 U47605 ( .A(n45459), .B(n45458), .Y(n45460) );
  NAND2X1 U47606 ( .A(n45461), .B(n45460), .Y(n45462) );
  NAND2X1 U47607 ( .A(n2986), .B(n42785), .Y(n45464) );
  NOR2X1 U47608 ( .A(n38822), .B(n45464), .Y(n45471) );
  NOR2X1 U47609 ( .A(n42867), .B(n39195), .Y(n45465) );
  NAND2X1 U47610 ( .A(n45465), .B(n3002), .Y(n45469) );
  NOR2X1 U47611 ( .A(n46927), .B(n45466), .Y(n45467) );
  NAND2X1 U47612 ( .A(n45467), .B(n40513), .Y(n45468) );
  NAND2X1 U47613 ( .A(n45469), .B(n45468), .Y(n45470) );
  NOR2X1 U47614 ( .A(n45471), .B(n45470), .Y(n45482) );
  NOR2X1 U47615 ( .A(n40534), .B(n39809), .Y(n45472) );
  NAND2X1 U47616 ( .A(n45472), .B(n2989), .Y(n45474) );
  NAND2X1 U47617 ( .A(n45662), .B(n3004), .Y(n45473) );
  NAND2X1 U47618 ( .A(n45474), .B(n45473), .Y(n45480) );
  NOR2X1 U47619 ( .A(n42765), .B(n40534), .Y(n45475) );
  NAND2X1 U47620 ( .A(n45475), .B(n2996), .Y(n45478) );
  NOR2X1 U47621 ( .A(n40866), .B(n39196), .Y(n45476) );
  NAND2X1 U47622 ( .A(n45476), .B(n2994), .Y(n45477) );
  NAND2X1 U47623 ( .A(n45478), .B(n45477), .Y(n45479) );
  NOR2X1 U47624 ( .A(n45480), .B(n45479), .Y(n45481) );
  NAND2X1 U47625 ( .A(n45482), .B(n45481), .Y(n45506) );
  NOR2X1 U47626 ( .A(n40529), .B(n45483), .Y(n45484) );
  NAND2X1 U47627 ( .A(n45484), .B(n40513), .Y(n45486) );
  NAND2X1 U47628 ( .A(n45754), .B(n3011), .Y(n45485) );
  NAND2X1 U47629 ( .A(n45486), .B(n45485), .Y(n45492) );
  NOR2X1 U47630 ( .A(n42767), .B(n42695), .Y(n45487) );
  NAND2X1 U47631 ( .A(n45487), .B(n2995), .Y(n45490) );
  NOR2X1 U47632 ( .A(n39809), .B(n39195), .Y(n45488) );
  NAND2X1 U47633 ( .A(n45488), .B(n2987), .Y(n45489) );
  NAND2X1 U47634 ( .A(n45490), .B(n45489), .Y(n45491) );
  NOR2X1 U47635 ( .A(n45492), .B(n45491), .Y(n45504) );
  NOR2X1 U47636 ( .A(n42868), .B(n40529), .Y(n45493) );
  NAND2X1 U47637 ( .A(n45493), .B(n3001), .Y(n45496) );
  NAND2X1 U47638 ( .A(n45494), .B(n42883), .Y(n45495) );
  NAND2X1 U47639 ( .A(n45496), .B(n45495), .Y(n45502) );
  NOR2X1 U47640 ( .A(n42766), .B(n40529), .Y(n45497) );
  NAND2X1 U47641 ( .A(n45497), .B(n2993), .Y(n45500) );
  NAND2X1 U47642 ( .A(n45498), .B(n42882), .Y(n45499) );
  NAND2X1 U47643 ( .A(n45500), .B(n45499), .Y(n45501) );
  NOR2X1 U47644 ( .A(n45502), .B(n45501), .Y(n45503) );
  NAND2X1 U47645 ( .A(n45504), .B(n45503), .Y(n45505) );
  NOR2X1 U47646 ( .A(n45506), .B(n45505), .Y(n45518) );
  NOR2X1 U47647 ( .A(n36841), .B(n49665), .Y(n45510) );
  NAND2X1 U47648 ( .A(n42883), .B(n42785), .Y(n45508) );
  NOR2X1 U47649 ( .A(n36848), .B(n45508), .Y(n45509) );
  NOR2X1 U47650 ( .A(n45510), .B(n45509), .Y(n45512) );
  NAND2X1 U47651 ( .A(n42618), .B(n1802), .Y(n45511) );
  NAND2X1 U47652 ( .A(n45512), .B(n45511), .Y(n45516) );
  INVX1 U47653 ( .A(n45871), .Y(n49685) );
  NAND2X1 U47654 ( .A(n49685), .B(n3003), .Y(n45514) );
  NAND2X1 U47655 ( .A(n40248), .B(n2988), .Y(n45513) );
  NAND2X1 U47656 ( .A(n45514), .B(n45513), .Y(n45515) );
  NOR2X1 U47657 ( .A(n45516), .B(n45515), .Y(n45517) );
  NAND2X1 U47658 ( .A(n45518), .B(n45517), .Y(n45519) );
  INVX1 U47659 ( .A(n42691), .Y(n45521) );
  INVX1 U47660 ( .A(n40685), .Y(n45922) );
  NOR2X1 U47661 ( .A(n46231), .B(n36935), .Y(n45523) );
  NOR2X1 U47662 ( .A(n46207), .B(n36940), .Y(n45524) );
  NOR2X1 U47663 ( .A(n38846), .B(n46009), .Y(n45527) );
  NOR2X1 U47664 ( .A(n57605), .B(n37045), .Y(n45526) );
  NAND2X1 U47665 ( .A(n45527), .B(n45526), .Y(n45528) );
  NAND2X1 U47666 ( .A(n45529), .B(n45528), .Y(n45542) );
  NOR2X1 U47667 ( .A(n42498), .B(n45530), .Y(n45532) );
  NOR2X1 U47668 ( .A(n45532), .B(n45531), .Y(n45535) );
  NAND2X1 U47669 ( .A(n45535), .B(n42373), .Y(n49715) );
  NAND2X1 U47670 ( .A(writeback_exec_value_w[29]), .B(n38805), .Y(n45540) );
  INVX1 U47671 ( .A(n38777), .Y(n46583) );
  NOR2X1 U47672 ( .A(n46583), .B(n43225), .Y(n45538) );
  NAND2X1 U47673 ( .A(n45538), .B(n45922), .Y(n45539) );
  NAND2X1 U47674 ( .A(n45540), .B(n45539), .Y(n45541) );
  NAND2X1 U47675 ( .A(n44028), .B(n43500), .Y(n57684) );
  INVX1 U47676 ( .A(mem_d_data_rd_i[30]), .Y(n45543) );
  NAND2X1 U47677 ( .A(n40935), .B(n45543), .Y(n45544) );
  NOR2X1 U47678 ( .A(n43455), .B(n43229), .Y(n45546) );
  NOR2X1 U47679 ( .A(n43022), .B(n43232), .Y(n45545) );
  NAND2X1 U47680 ( .A(n2982), .B(n43362), .Y(n45548) );
  NAND2X1 U47681 ( .A(n2957), .B(n38410), .Y(n45547) );
  NAND2X1 U47682 ( .A(n45548), .B(n45547), .Y(n45552) );
  NAND2X1 U47683 ( .A(n2964), .B(n43343), .Y(n45550) );
  NAND2X1 U47684 ( .A(n2972), .B(n43027), .Y(n45549) );
  NAND2X1 U47685 ( .A(n45550), .B(n45549), .Y(n45551) );
  NOR2X1 U47686 ( .A(n45552), .B(n45551), .Y(n45560) );
  NAND2X1 U47687 ( .A(n2954), .B(n43030), .Y(n45554) );
  NAND2X1 U47688 ( .A(n2959), .B(n43032), .Y(n45553) );
  NAND2X1 U47689 ( .A(n45554), .B(n45553), .Y(n45558) );
  NAND2X1 U47690 ( .A(n2974), .B(n43036), .Y(n45556) );
  NAND2X1 U47691 ( .A(n2966), .B(n43351), .Y(n45555) );
  NAND2X1 U47692 ( .A(n45556), .B(n45555), .Y(n45557) );
  NOR2X1 U47693 ( .A(n45558), .B(n45557), .Y(n45559) );
  NAND2X1 U47694 ( .A(n45560), .B(n45559), .Y(n45576) );
  NAND2X1 U47695 ( .A(n2970), .B(n43356), .Y(n45562) );
  NAND2X1 U47696 ( .A(n2968), .B(n43039), .Y(n45561) );
  NAND2X1 U47697 ( .A(n45562), .B(n45561), .Y(n45566) );
  NAND2X1 U47698 ( .A(n1789), .B(n39804), .Y(n45564) );
  NAND2X1 U47699 ( .A(n2976), .B(n43042), .Y(n45563) );
  NAND2X1 U47700 ( .A(n45564), .B(n45563), .Y(n45565) );
  NOR2X1 U47701 ( .A(n45566), .B(n45565), .Y(n45574) );
  NAND2X1 U47702 ( .A(n2980), .B(n43359), .Y(n45568) );
  NAND2X1 U47703 ( .A(n2955), .B(n43345), .Y(n45567) );
  NAND2X1 U47704 ( .A(n45568), .B(n45567), .Y(n45572) );
  NAND2X1 U47705 ( .A(n2962), .B(n43338), .Y(n45570) );
  NAND2X1 U47706 ( .A(n2978), .B(n43365), .Y(n45569) );
  NAND2X1 U47707 ( .A(n45570), .B(n45569), .Y(n45571) );
  NOR2X1 U47708 ( .A(n45572), .B(n45571), .Y(n45573) );
  NAND2X1 U47709 ( .A(n45574), .B(n45573), .Y(n45575) );
  NOR2X1 U47710 ( .A(n45576), .B(n45575), .Y(n45606) );
  NAND2X1 U47711 ( .A(n2975), .B(n43044), .Y(n45578) );
  NAND2X1 U47712 ( .A(n2981), .B(n43047), .Y(n45577) );
  NAND2X1 U47713 ( .A(n45578), .B(n45577), .Y(n45582) );
  NAND2X1 U47714 ( .A(n2973), .B(n43049), .Y(n45580) );
  NAND2X1 U47715 ( .A(n2958), .B(n43051), .Y(n45579) );
  NAND2X1 U47716 ( .A(n45580), .B(n45579), .Y(n45581) );
  NOR2X1 U47717 ( .A(n45582), .B(n45581), .Y(n45588) );
  NOR2X1 U47718 ( .A(n43371), .B(n36823), .Y(n45586) );
  NAND2X1 U47719 ( .A(n2960), .B(n43054), .Y(n45584) );
  NAND2X1 U47720 ( .A(n1790), .B(n43057), .Y(n45583) );
  NAND2X1 U47721 ( .A(n45584), .B(n45583), .Y(n45585) );
  NOR2X1 U47722 ( .A(n45586), .B(n45585), .Y(n45587) );
  NAND2X1 U47723 ( .A(n45588), .B(n45587), .Y(n45604) );
  NAND2X1 U47724 ( .A(n2979), .B(n43060), .Y(n45590) );
  NAND2X1 U47725 ( .A(n2977), .B(n39136), .Y(n45589) );
  NAND2X1 U47726 ( .A(n45590), .B(n45589), .Y(n45594) );
  NAND2X1 U47727 ( .A(n2969), .B(n43063), .Y(n45592) );
  NAND2X1 U47728 ( .A(n2961), .B(n43067), .Y(n45591) );
  NAND2X1 U47729 ( .A(n45592), .B(n45591), .Y(n45593) );
  NOR2X1 U47730 ( .A(n45594), .B(n45593), .Y(n45602) );
  NAND2X1 U47731 ( .A(n2965), .B(n43372), .Y(n45596) );
  NAND2X1 U47732 ( .A(n2971), .B(n43349), .Y(n45595) );
  NAND2X1 U47733 ( .A(n45596), .B(n45595), .Y(n45600) );
  NAND2X1 U47734 ( .A(n2963), .B(n43070), .Y(n45598) );
  NAND2X1 U47735 ( .A(n2956), .B(n43071), .Y(n45597) );
  NAND2X1 U47736 ( .A(n45598), .B(n45597), .Y(n45599) );
  NOR2X1 U47737 ( .A(n45600), .B(n45599), .Y(n45601) );
  NAND2X1 U47738 ( .A(n45602), .B(n45601), .Y(n45603) );
  NOR2X1 U47739 ( .A(n45604), .B(n45603), .Y(n45605) );
  NAND2X1 U47740 ( .A(n45606), .B(n45605), .Y(n45607) );
  INVX1 U47741 ( .A(n45615), .Y(n45609) );
  NOR2X1 U47742 ( .A(n45609), .B(n45608), .Y(n45613) );
  INVX1 U47743 ( .A(n42691), .Y(n45612) );
  INVX1 U47744 ( .A(n46231), .Y(n45614) );
  NOR2X1 U47745 ( .A(n45616), .B(n45696), .Y(n45617) );
  NOR2X1 U47746 ( .A(n45618), .B(n45617), .Y(n45624) );
  NOR2X1 U47747 ( .A(n38662), .B(n38807), .Y(n45621) );
  NOR2X1 U47748 ( .A(n45621), .B(n45620), .Y(n45622) );
  NAND2X1 U47749 ( .A(n45622), .B(n40152), .Y(n45623) );
  NAND2X1 U47750 ( .A(n45624), .B(n45623), .Y(n45625) );
  NOR2X1 U47751 ( .A(n45626), .B(n45625), .Y(n60952) );
  NAND2X1 U47752 ( .A(n2980), .B(n40513), .Y(n45627) );
  NOR2X1 U47753 ( .A(n38821), .B(n45627), .Y(n45630) );
  NAND2X1 U47754 ( .A(n2981), .B(n39197), .Y(n45628) );
  NOR2X1 U47755 ( .A(n40511), .B(n45628), .Y(n45629) );
  NOR2X1 U47756 ( .A(n45630), .B(n45629), .Y(n45639) );
  NOR2X1 U47757 ( .A(n45631), .B(n40508), .Y(n45634) );
  NAND2X1 U47758 ( .A(n42759), .B(opcode_opcode_w[24]), .Y(n45632) );
  NOR2X1 U47759 ( .A(n36792), .B(n45632), .Y(n45633) );
  NOR2X1 U47760 ( .A(n45634), .B(n45633), .Y(n45636) );
  NAND2X1 U47761 ( .A(n2970), .B(n46049), .Y(n45635) );
  NAND2X1 U47762 ( .A(n45636), .B(n45635), .Y(n45637) );
  NAND2X1 U47763 ( .A(n38492), .B(n45637), .Y(n45638) );
  NAND2X1 U47764 ( .A(n45639), .B(n45638), .Y(n45650) );
  NAND2X1 U47765 ( .A(n42696), .B(n40512), .Y(n45640) );
  NOR2X1 U47766 ( .A(n36824), .B(n49677), .Y(n45642) );
  NOR2X1 U47767 ( .A(n45642), .B(n45641), .Y(n45648) );
  NAND2X1 U47768 ( .A(n45764), .B(n1790), .Y(n45644) );
  NAND2X1 U47769 ( .A(n45465), .B(n2973), .Y(n45643) );
  NAND2X1 U47770 ( .A(n45644), .B(n45643), .Y(n45645) );
  NOR2X1 U47771 ( .A(n45646), .B(n45645), .Y(n45647) );
  NAND2X1 U47772 ( .A(n45648), .B(n45647), .Y(n45649) );
  NOR2X1 U47773 ( .A(n45650), .B(n45649), .Y(n45677) );
  NAND2X1 U47774 ( .A(n46183), .B(n42773), .Y(n45651) );
  NOR2X1 U47775 ( .A(n36823), .B(n42895), .Y(n45653) );
  NOR2X1 U47776 ( .A(n45653), .B(n45652), .Y(n45658) );
  NAND2X1 U47777 ( .A(n38824), .B(n42773), .Y(n45654) );
  NOR2X1 U47778 ( .A(n36827), .B(n45654), .Y(n45655) );
  NOR2X1 U47779 ( .A(n45656), .B(n45655), .Y(n45657) );
  NAND2X1 U47780 ( .A(n45658), .B(n45657), .Y(n45675) );
  NOR2X1 U47781 ( .A(n42868), .B(n36793), .Y(n45660) );
  NOR2X1 U47782 ( .A(n39809), .B(n36794), .Y(n45659) );
  NOR2X1 U47783 ( .A(n45660), .B(n45659), .Y(n45661) );
  NOR2X1 U47784 ( .A(n45661), .B(n42693), .Y(n45667) );
  NOR2X1 U47785 ( .A(n40534), .B(n42866), .Y(n45662) );
  NAND2X1 U47786 ( .A(n45662), .B(n2975), .Y(n45665) );
  NOR2X1 U47787 ( .A(n45199), .B(n39196), .Y(n45663) );
  NAND2X1 U47788 ( .A(n45663), .B(n2958), .Y(n45664) );
  NAND2X1 U47789 ( .A(n45665), .B(n45664), .Y(n45666) );
  NOR2X1 U47790 ( .A(n45667), .B(n45666), .Y(n45673) );
  NAND2X1 U47791 ( .A(n2962), .B(n42772), .Y(n45668) );
  NOR2X1 U47792 ( .A(n42881), .B(n45668), .Y(n45671) );
  NAND2X1 U47793 ( .A(n38825), .B(n42676), .Y(n45669) );
  NOR2X1 U47794 ( .A(n36834), .B(n45669), .Y(n45670) );
  NOR2X1 U47795 ( .A(n45671), .B(n45670), .Y(n45672) );
  NAND2X1 U47796 ( .A(n45673), .B(n45672), .Y(n45674) );
  NOR2X1 U47797 ( .A(n45675), .B(n45674), .Y(n45676) );
  NAND2X1 U47798 ( .A(n45677), .B(n45676), .Y(n45678) );
  NAND2X1 U47799 ( .A(n61188), .B(n45678), .Y(n60951) );
  NAND2X1 U47800 ( .A(n2971), .B(n40447), .Y(n45680) );
  NAND2X1 U47801 ( .A(n45188), .B(n42692), .Y(n45679) );
  NOR2X1 U47802 ( .A(n45680), .B(n45679), .Y(n45684) );
  INVX1 U47803 ( .A(n46570), .Y(n46404) );
  NAND2X1 U47804 ( .A(n46404), .B(n2968), .Y(n45682) );
  NAND2X1 U47805 ( .A(n45710), .B(n45188), .Y(n45681) );
  NOR2X1 U47806 ( .A(n45682), .B(n45681), .Y(n45683) );
  OR2X1 U47807 ( .A(n45684), .B(n45683), .Y(n45692) );
  INVX1 U47808 ( .A(n46575), .Y(n46906) );
  NAND2X1 U47809 ( .A(n46906), .B(n1789), .Y(n45686) );
  NAND2X1 U47810 ( .A(n46019), .B(n45188), .Y(n45685) );
  NOR2X1 U47811 ( .A(n45686), .B(n45685), .Y(n45690) );
  NAND2X1 U47812 ( .A(n46979), .B(n2961), .Y(n45688) );
  NAND2X1 U47813 ( .A(n38441), .B(n45710), .Y(n45687) );
  NOR2X1 U47814 ( .A(n45688), .B(n45687), .Y(n45689) );
  OR2X1 U47815 ( .A(n45690), .B(n45689), .Y(n45691) );
  NOR2X1 U47816 ( .A(n45692), .B(n45691), .Y(n60950) );
  NAND2X1 U47817 ( .A(n37355), .B(n38777), .Y(n45693) );
  NOR2X1 U47818 ( .A(n40152), .B(n45693), .Y(n45695) );
  NOR2X1 U47819 ( .A(n43232), .B(n49715), .Y(n45694) );
  NAND2X1 U47820 ( .A(n40035), .B(n2969), .Y(n45697) );
  NAND2X1 U47821 ( .A(n45710), .B(n40398), .Y(n45696) );
  NOR2X1 U47822 ( .A(n45697), .B(n45696), .Y(n45701) );
  INVX1 U47823 ( .A(n46206), .Y(n46309) );
  NAND2X1 U47824 ( .A(n46309), .B(n2977), .Y(n45699) );
  NAND2X1 U47825 ( .A(n38441), .B(n42705), .Y(n45698) );
  NOR2X1 U47826 ( .A(n45699), .B(n45698), .Y(n45700) );
  NAND2X1 U47827 ( .A(n44051), .B(n39961), .Y(n57677) );
  NAND2X1 U47828 ( .A(n57684), .B(n57677), .Y(n49878) );
  NAND2X1 U47829 ( .A(n44811), .B(n49878), .Y(n45702) );
  NAND2X1 U47830 ( .A(n31124), .B(n45702), .Y(n49896) );
  NAND2X1 U47831 ( .A(n44059), .B(n43607), .Y(n58159) );
  NAND2X1 U47832 ( .A(n45704), .B(n44815), .Y(n49894) );
  INVX1 U47833 ( .A(n49894), .Y(n45705) );
  NOR2X1 U47834 ( .A(n45922), .B(n38846), .Y(n45707) );
  NOR2X1 U47835 ( .A(n46207), .B(n37054), .Y(n45706) );
  NAND2X1 U47836 ( .A(n45707), .B(n45706), .Y(n45708) );
  NAND2X1 U47837 ( .A(n45709), .B(n45708), .Y(n45717) );
  NOR2X1 U47838 ( .A(n57605), .B(n37046), .Y(n45711) );
  NAND2X1 U47839 ( .A(n45711), .B(n40499), .Y(n45715) );
  NOR2X1 U47840 ( .A(n46372), .B(n37053), .Y(n45713) );
  INVX1 U47841 ( .A(n42704), .Y(n46526) );
  NOR2X1 U47842 ( .A(n46009), .B(n45612), .Y(n45712) );
  NAND2X1 U47843 ( .A(n45713), .B(n45712), .Y(n45714) );
  NAND2X1 U47844 ( .A(n45715), .B(n45714), .Y(n45716) );
  NOR2X1 U47845 ( .A(n45717), .B(n45716), .Y(n45773) );
  INVX1 U47846 ( .A(n49699), .Y(n49621) );
  NOR2X1 U47847 ( .A(n42866), .B(n36803), .Y(n45718) );
  NAND2X1 U47848 ( .A(n45718), .B(n38824), .Y(n45721) );
  NOR2X1 U47849 ( .A(n42765), .B(n36804), .Y(n45719) );
  NAND2X1 U47850 ( .A(n45719), .B(n38824), .Y(n45720) );
  NAND2X1 U47851 ( .A(n45721), .B(n45720), .Y(n45727) );
  NOR2X1 U47852 ( .A(n42766), .B(n36806), .Y(n45722) );
  NAND2X1 U47853 ( .A(n45722), .B(n42882), .Y(n45725) );
  NOR2X1 U47854 ( .A(n42866), .B(n36809), .Y(n45723) );
  NAND2X1 U47855 ( .A(n45723), .B(n42882), .Y(n45724) );
  NAND2X1 U47856 ( .A(n45725), .B(n45724), .Y(n45726) );
  NOR2X1 U47857 ( .A(n45727), .B(n45726), .Y(n45738) );
  NOR2X1 U47858 ( .A(n42767), .B(n36805), .Y(n45729) );
  NOR2X1 U47859 ( .A(n45199), .B(n36808), .Y(n45728) );
  NOR2X1 U47860 ( .A(n45729), .B(n45728), .Y(n45730) );
  NOR2X1 U47861 ( .A(n45730), .B(n40534), .Y(n45736) );
  NOR2X1 U47862 ( .A(n45199), .B(n36807), .Y(n45731) );
  NAND2X1 U47863 ( .A(n45731), .B(n38825), .Y(n45734) );
  NOR2X1 U47864 ( .A(n39809), .B(n36811), .Y(n45732) );
  NAND2X1 U47865 ( .A(n45732), .B(n42883), .Y(n45733) );
  NAND2X1 U47866 ( .A(n45734), .B(n45733), .Y(n45735) );
  NOR2X1 U47867 ( .A(n45736), .B(n45735), .Y(n45737) );
  NAND2X1 U47868 ( .A(n45738), .B(n45737), .Y(n45751) );
  NAND2X1 U47869 ( .A(n39197), .B(n46049), .Y(n45739) );
  NOR2X1 U47870 ( .A(n36866), .B(n45739), .Y(n45741) );
  NOR2X1 U47871 ( .A(n45741), .B(n45740), .Y(n45749) );
  NAND2X1 U47872 ( .A(n39198), .B(n42785), .Y(n45742) );
  NOR2X1 U47873 ( .A(n36870), .B(n45742), .Y(n45747) );
  NAND2X1 U47874 ( .A(n46178), .B(n2216), .Y(n45745) );
  NOR2X1 U47875 ( .A(n40511), .B(n36813), .Y(n45743) );
  NAND2X1 U47876 ( .A(n45743), .B(n38824), .Y(n45744) );
  NAND2X1 U47877 ( .A(n45745), .B(n45744), .Y(n45746) );
  NOR2X1 U47878 ( .A(n45747), .B(n45746), .Y(n45748) );
  NAND2X1 U47879 ( .A(n45749), .B(n45748), .Y(n45750) );
  NOR2X1 U47880 ( .A(n45751), .B(n45750), .Y(n45770) );
  INVX1 U47881 ( .A(n42859), .Y(n47895) );
  NAND2X1 U47882 ( .A(n47895), .B(n2219), .Y(n45753) );
  NAND2X1 U47883 ( .A(n42679), .B(n2213), .Y(n45752) );
  NAND2X1 U47884 ( .A(n45753), .B(n45752), .Y(n45768) );
  NOR2X1 U47885 ( .A(n40508), .B(n42695), .Y(n45754) );
  NAND2X1 U47886 ( .A(n45754), .B(n2220), .Y(n45757) );
  NOR2X1 U47887 ( .A(n45200), .B(n42700), .Y(n45755) );
  NAND2X1 U47888 ( .A(n45755), .B(n2204), .Y(n45756) );
  NAND2X1 U47889 ( .A(n45757), .B(n45756), .Y(n45763) );
  NOR2X1 U47890 ( .A(n42700), .B(n42868), .Y(n45758) );
  NAND2X1 U47891 ( .A(n45758), .B(n2212), .Y(n45761) );
  NOR2X1 U47892 ( .A(n45199), .B(n42700), .Y(n45759) );
  NAND2X1 U47893 ( .A(n45759), .B(n2197), .Y(n45760) );
  NAND2X1 U47894 ( .A(n45761), .B(n45760), .Y(n45762) );
  NOR2X1 U47895 ( .A(n45763), .B(n45762), .Y(n45766) );
  NOR2X1 U47896 ( .A(n40510), .B(n40534), .Y(n45764) );
  NAND2X1 U47897 ( .A(n45764), .B(n1804), .Y(n45765) );
  NAND2X1 U47898 ( .A(n45766), .B(n45765), .Y(n45767) );
  NOR2X1 U47899 ( .A(n45768), .B(n45767), .Y(n45769) );
  NAND2X1 U47900 ( .A(n45770), .B(n45769), .Y(n45771) );
  NAND2X1 U47901 ( .A(n40490), .B(n45771), .Y(n45772) );
  NAND2X1 U47902 ( .A(n45773), .B(n45772), .Y(n60235) );
  NOR2X1 U47903 ( .A(n46575), .B(n37030), .Y(n45774) );
  NAND2X1 U47904 ( .A(n46019), .B(n42671), .Y(n46394) );
  NAND2X1 U47905 ( .A(n45774), .B(n38604), .Y(n45777) );
  NOR2X1 U47906 ( .A(n46231), .B(n37035), .Y(n45775) );
  NAND2X1 U47907 ( .A(n45775), .B(n38604), .Y(n45776) );
  NAND2X1 U47908 ( .A(n45777), .B(n45776), .Y(n45782) );
  NOR2X1 U47909 ( .A(n46007), .B(n37044), .Y(n45778) );
  NAND2X1 U47910 ( .A(n45778), .B(n42149), .Y(n45779) );
  NAND2X1 U47911 ( .A(n45780), .B(n45779), .Y(n45781) );
  NAND2X1 U47912 ( .A(n40935), .B(n373), .Y(n45783) );
  NAND2X1 U47913 ( .A(n45783), .B(n42876), .Y(n56124) );
  NAND2X1 U47914 ( .A(writeback_exec_value_w[28]), .B(n37976), .Y(n45784) );
  NAND2X1 U47915 ( .A(n45785), .B(n45784), .Y(n45793) );
  NOR2X1 U47916 ( .A(n46570), .B(n37042), .Y(n45786) );
  NAND2X1 U47917 ( .A(n45786), .B(n46412), .Y(n45791) );
  NAND2X1 U47918 ( .A(n2214), .B(n46741), .Y(n45788) );
  NAND2X1 U47919 ( .A(n2217), .B(n40404), .Y(n45787) );
  NAND2X1 U47920 ( .A(n45788), .B(n45787), .Y(n45789) );
  NAND2X1 U47921 ( .A(n46412), .B(n45789), .Y(n45790) );
  NAND2X1 U47922 ( .A(n45791), .B(n45790), .Y(n45792) );
  NOR2X1 U47923 ( .A(n43455), .B(n43217), .Y(n45795) );
  NOR2X1 U47924 ( .A(n43022), .B(n43220), .Y(n45794) );
  NAND2X1 U47925 ( .A(n2220), .B(n43362), .Y(n45797) );
  NAND2X1 U47926 ( .A(n2195), .B(n38408), .Y(n45796) );
  NAND2X1 U47927 ( .A(n45797), .B(n45796), .Y(n45801) );
  NAND2X1 U47928 ( .A(n2202), .B(n43342), .Y(n45799) );
  NAND2X1 U47929 ( .A(n2210), .B(n43027), .Y(n45798) );
  NAND2X1 U47930 ( .A(n45799), .B(n45798), .Y(n45800) );
  NOR2X1 U47931 ( .A(n45801), .B(n45800), .Y(n45809) );
  NAND2X1 U47932 ( .A(n2192), .B(n43030), .Y(n45803) );
  NAND2X1 U47933 ( .A(n2197), .B(n43032), .Y(n45802) );
  NAND2X1 U47934 ( .A(n45803), .B(n45802), .Y(n45807) );
  NAND2X1 U47935 ( .A(n2212), .B(n43036), .Y(n45805) );
  NAND2X1 U47936 ( .A(n2204), .B(n43351), .Y(n45804) );
  NAND2X1 U47937 ( .A(n45805), .B(n45804), .Y(n45806) );
  NOR2X1 U47938 ( .A(n45807), .B(n45806), .Y(n45808) );
  NAND2X1 U47939 ( .A(n45809), .B(n45808), .Y(n45825) );
  NAND2X1 U47940 ( .A(n2208), .B(n43356), .Y(n45811) );
  NAND2X1 U47941 ( .A(n2206), .B(n43039), .Y(n45810) );
  NAND2X1 U47942 ( .A(n45811), .B(n45810), .Y(n45815) );
  NAND2X1 U47943 ( .A(n1803), .B(n39802), .Y(n45813) );
  NAND2X1 U47944 ( .A(n2214), .B(n43042), .Y(n45812) );
  NAND2X1 U47945 ( .A(n45813), .B(n45812), .Y(n45814) );
  NOR2X1 U47946 ( .A(n45815), .B(n45814), .Y(n45823) );
  NAND2X1 U47947 ( .A(n2218), .B(n43358), .Y(n45817) );
  NAND2X1 U47948 ( .A(n2193), .B(n43345), .Y(n45816) );
  NAND2X1 U47949 ( .A(n45817), .B(n45816), .Y(n45821) );
  NAND2X1 U47950 ( .A(n2200), .B(n43338), .Y(n45819) );
  NAND2X1 U47951 ( .A(n2216), .B(n43365), .Y(n45818) );
  NAND2X1 U47952 ( .A(n45819), .B(n45818), .Y(n45820) );
  NOR2X1 U47953 ( .A(n45821), .B(n45820), .Y(n45822) );
  NAND2X1 U47954 ( .A(n45823), .B(n45822), .Y(n45824) );
  NOR2X1 U47955 ( .A(n45825), .B(n45824), .Y(n45855) );
  NAND2X1 U47956 ( .A(n2213), .B(n43044), .Y(n45827) );
  NAND2X1 U47957 ( .A(n2219), .B(n43047), .Y(n45826) );
  NAND2X1 U47958 ( .A(n45827), .B(n45826), .Y(n45831) );
  NAND2X1 U47959 ( .A(n2211), .B(n43049), .Y(n45829) );
  NAND2X1 U47960 ( .A(n2196), .B(n43051), .Y(n45828) );
  NAND2X1 U47961 ( .A(n45829), .B(n45828), .Y(n45830) );
  NOR2X1 U47962 ( .A(n45831), .B(n45830), .Y(n45837) );
  NOR2X1 U47963 ( .A(n43370), .B(n36805), .Y(n45835) );
  NAND2X1 U47964 ( .A(n2198), .B(n43054), .Y(n45833) );
  NAND2X1 U47965 ( .A(n1804), .B(n43057), .Y(n45832) );
  NAND2X1 U47966 ( .A(n45833), .B(n45832), .Y(n45834) );
  NOR2X1 U47967 ( .A(n45835), .B(n45834), .Y(n45836) );
  NAND2X1 U47968 ( .A(n45837), .B(n45836), .Y(n45853) );
  NAND2X1 U47969 ( .A(n2217), .B(n43060), .Y(n45839) );
  NAND2X1 U47970 ( .A(n2215), .B(n39134), .Y(n45838) );
  NAND2X1 U47971 ( .A(n45839), .B(n45838), .Y(n45843) );
  NAND2X1 U47972 ( .A(n2207), .B(n43063), .Y(n45841) );
  NAND2X1 U47973 ( .A(n2199), .B(n43067), .Y(n45840) );
  NAND2X1 U47974 ( .A(n45841), .B(n45840), .Y(n45842) );
  NOR2X1 U47975 ( .A(n45843), .B(n45842), .Y(n45851) );
  NAND2X1 U47976 ( .A(n2203), .B(n43372), .Y(n45845) );
  NAND2X1 U47977 ( .A(n2209), .B(n43350), .Y(n45844) );
  NAND2X1 U47978 ( .A(n45845), .B(n45844), .Y(n45849) );
  NAND2X1 U47979 ( .A(n2201), .B(n43070), .Y(n45847) );
  NAND2X1 U47980 ( .A(n2194), .B(n43071), .Y(n45846) );
  NAND2X1 U47981 ( .A(n45847), .B(n45846), .Y(n45848) );
  NOR2X1 U47982 ( .A(n45849), .B(n45848), .Y(n45850) );
  NAND2X1 U47983 ( .A(n45851), .B(n45850), .Y(n45852) );
  NOR2X1 U47984 ( .A(n45853), .B(n45852), .Y(n45854) );
  NAND2X1 U47985 ( .A(n45855), .B(n45854), .Y(n45856) );
  NAND2X1 U47986 ( .A(n43498), .B(n44016), .Y(n57695) );
  NOR2X1 U47987 ( .A(n46206), .B(n37019), .Y(n45857) );
  NAND2X1 U47988 ( .A(n45857), .B(n40590), .Y(n45860) );
  NOR2X1 U47989 ( .A(n46372), .B(n37021), .Y(n45858) );
  NAND2X1 U47990 ( .A(n45707), .B(n45858), .Y(n45859) );
  NAND2X1 U47991 ( .A(n45860), .B(n45859), .Y(n45866) );
  NOR2X1 U47992 ( .A(n57605), .B(n37023), .Y(n45861) );
  NAND2X1 U47993 ( .A(n45457), .B(n45861), .Y(n45864) );
  NOR2X1 U47994 ( .A(n46207), .B(n37020), .Y(n45862) );
  NAND2X1 U47995 ( .A(n45862), .B(n40499), .Y(n45863) );
  NAND2X1 U47996 ( .A(n45864), .B(n45863), .Y(n45865) );
  NOR2X1 U47997 ( .A(n36836), .B(n36609), .Y(n45869) );
  INVX1 U47998 ( .A(n2807), .Y(n45867) );
  NOR2X1 U47999 ( .A(n42682), .B(n45867), .Y(n45868) );
  NOR2X1 U48000 ( .A(n45869), .B(n45868), .Y(n45875) );
  NAND2X1 U48001 ( .A(n42699), .B(n39449), .Y(n45870) );
  NOR2X1 U48002 ( .A(n36837), .B(n45870), .Y(n45873) );
  NOR2X1 U48003 ( .A(n36839), .B(n45871), .Y(n45872) );
  NOR2X1 U48004 ( .A(n45873), .B(n45872), .Y(n45874) );
  NAND2X1 U48005 ( .A(n45875), .B(n45874), .Y(n45891) );
  NOR2X1 U48006 ( .A(n40509), .B(n38823), .Y(n45876) );
  NAND2X1 U48007 ( .A(n45876), .B(n2812), .Y(n45879) );
  NOR2X1 U48008 ( .A(n40866), .B(n36798), .Y(n45877) );
  NAND2X1 U48009 ( .A(n45877), .B(n42882), .Y(n45878) );
  NAND2X1 U48010 ( .A(n45879), .B(n45878), .Y(n45884) );
  NOR2X1 U48011 ( .A(n40511), .B(n42694), .Y(n45880) );
  NAND2X1 U48012 ( .A(n45880), .B(n2814), .Y(n45882) );
  NAND2X1 U48013 ( .A(n45475), .B(n2799), .Y(n45881) );
  NAND2X1 U48014 ( .A(n45882), .B(n45881), .Y(n45883) );
  NOR2X1 U48015 ( .A(n45884), .B(n45883), .Y(n45889) );
  NOR2X1 U48016 ( .A(n36840), .B(n42776), .Y(n45887) );
  INVX1 U48017 ( .A(n2804), .Y(n45885) );
  NOR2X1 U48018 ( .A(n45885), .B(n45245), .Y(n45886) );
  NOR2X1 U48019 ( .A(n45887), .B(n45886), .Y(n45888) );
  NAND2X1 U48020 ( .A(n45889), .B(n45888), .Y(n45890) );
  NOR2X1 U48021 ( .A(n42868), .B(n42881), .Y(n45892) );
  NAND2X1 U48022 ( .A(n45892), .B(n2802), .Y(n45893) );
  NAND2X1 U48023 ( .A(n45894), .B(n45893), .Y(n45899) );
  NOR2X1 U48024 ( .A(n46927), .B(n42867), .Y(n45895) );
  NAND2X1 U48025 ( .A(n45895), .B(n2805), .Y(n45897) );
  NAND2X1 U48026 ( .A(n46948), .B(n2810), .Y(n45896) );
  NAND2X1 U48027 ( .A(n45897), .B(n45896), .Y(n45898) );
  NOR2X1 U48028 ( .A(n45899), .B(n45898), .Y(n45905) );
  NAND2X1 U48029 ( .A(n2815), .B(n36665), .Y(n45900) );
  NOR2X1 U48030 ( .A(n40507), .B(n45900), .Y(n45903) );
  NAND2X1 U48031 ( .A(n2789), .B(n38824), .Y(n45901) );
  NOR2X1 U48032 ( .A(n45199), .B(n45901), .Y(n45902) );
  NOR2X1 U48033 ( .A(n45903), .B(n45902), .Y(n45904) );
  NAND2X1 U48034 ( .A(n45905), .B(n45904), .Y(n45915) );
  NOR2X1 U48035 ( .A(n36842), .B(n39654), .Y(n45907) );
  NOR2X1 U48036 ( .A(n36851), .B(n40907), .Y(n45906) );
  NOR2X1 U48037 ( .A(n45907), .B(n45906), .Y(n45913) );
  NAND2X1 U48038 ( .A(n38947), .B(n42770), .Y(n49604) );
  NOR2X1 U48039 ( .A(n36845), .B(n49604), .Y(n45911) );
  INVX1 U48040 ( .A(n2813), .Y(n45909) );
  NAND2X1 U48041 ( .A(n40593), .B(n40513), .Y(n45908) );
  NOR2X1 U48042 ( .A(n45909), .B(n45908), .Y(n45910) );
  NOR2X1 U48043 ( .A(n45911), .B(n45910), .Y(n45912) );
  NAND2X1 U48044 ( .A(n45913), .B(n45912), .Y(n45914) );
  NOR2X1 U48045 ( .A(n46570), .B(n37033), .Y(n45917) );
  NAND2X1 U48046 ( .A(n46412), .B(n45917), .Y(n45920) );
  NOR2X1 U48047 ( .A(n46231), .B(n37027), .Y(n45918) );
  NAND2X1 U48048 ( .A(n45918), .B(n38604), .Y(n45919) );
  NAND2X1 U48049 ( .A(n45920), .B(n45919), .Y(n45924) );
  NOR2X1 U48050 ( .A(n46007), .B(n37036), .Y(n45921) );
  NOR2X1 U48051 ( .A(n45924), .B(n45923), .Y(n45939) );
  NAND2X1 U48052 ( .A(n2808), .B(n46741), .Y(n45926) );
  NAND2X1 U48053 ( .A(n45610), .B(n45188), .Y(n45925) );
  NOR2X1 U48054 ( .A(n45926), .B(n45925), .Y(n45928) );
  NOR2X1 U48055 ( .A(n42645), .B(n43213), .Y(n45927) );
  NOR2X1 U48056 ( .A(n45928), .B(n45927), .Y(n45931) );
  NAND2X1 U48057 ( .A(n40935), .B(n384), .Y(n45929) );
  NAND2X1 U48058 ( .A(n45929), .B(n42877), .Y(n55947) );
  NAND2X1 U48059 ( .A(n45931), .B(n45930), .Y(n45937) );
  NOR2X1 U48060 ( .A(n46236), .B(n37025), .Y(n45932) );
  NAND2X1 U48061 ( .A(n45932), .B(n42146), .Y(n45935) );
  NOR2X1 U48062 ( .A(n46575), .B(n37031), .Y(n45933) );
  NAND2X1 U48063 ( .A(n45933), .B(n38604), .Y(n45934) );
  NAND2X1 U48064 ( .A(n45935), .B(n45934), .Y(n45936) );
  NOR2X1 U48065 ( .A(n45937), .B(n45936), .Y(n45938) );
  NAND2X1 U48066 ( .A(n38614), .B(n40574), .Y(n71033) );
  NAND2X1 U48067 ( .A(n40935), .B(n395), .Y(n45940) );
  NOR2X1 U48068 ( .A(n43455), .B(n43204), .Y(n45942) );
  NOR2X1 U48069 ( .A(n43022), .B(n43207), .Y(n45941) );
  NAND2X1 U48070 ( .A(n2647), .B(n43362), .Y(n45944) );
  NAND2X1 U48071 ( .A(n2622), .B(n38406), .Y(n45943) );
  NAND2X1 U48072 ( .A(n45944), .B(n45943), .Y(n45948) );
  NAND2X1 U48073 ( .A(n2629), .B(n43343), .Y(n45946) );
  NAND2X1 U48074 ( .A(n2637), .B(n43027), .Y(n45945) );
  NAND2X1 U48075 ( .A(n45946), .B(n45945), .Y(n45947) );
  NOR2X1 U48076 ( .A(n45948), .B(n45947), .Y(n45956) );
  NAND2X1 U48077 ( .A(n2619), .B(n43030), .Y(n45950) );
  NAND2X1 U48078 ( .A(n2624), .B(n43032), .Y(n45949) );
  NAND2X1 U48079 ( .A(n45950), .B(n45949), .Y(n45954) );
  NAND2X1 U48080 ( .A(n2639), .B(n43036), .Y(n45952) );
  NAND2X1 U48081 ( .A(n2631), .B(n43351), .Y(n45951) );
  NAND2X1 U48082 ( .A(n45952), .B(n45951), .Y(n45953) );
  NOR2X1 U48083 ( .A(n45954), .B(n45953), .Y(n45955) );
  NAND2X1 U48084 ( .A(n45956), .B(n45955), .Y(n45972) );
  NAND2X1 U48085 ( .A(n2635), .B(n43356), .Y(n45958) );
  NAND2X1 U48086 ( .A(n2633), .B(n43039), .Y(n45957) );
  NAND2X1 U48087 ( .A(n45958), .B(n45957), .Y(n45962) );
  NAND2X1 U48088 ( .A(n1820), .B(n39808), .Y(n45960) );
  NAND2X1 U48089 ( .A(n2641), .B(n43042), .Y(n45959) );
  NAND2X1 U48090 ( .A(n45960), .B(n45959), .Y(n45961) );
  NOR2X1 U48091 ( .A(n45962), .B(n45961), .Y(n45970) );
  NAND2X1 U48092 ( .A(n2645), .B(n43359), .Y(n45964) );
  NAND2X1 U48093 ( .A(n2620), .B(n43345), .Y(n45963) );
  NAND2X1 U48094 ( .A(n45964), .B(n45963), .Y(n45968) );
  NAND2X1 U48095 ( .A(n2627), .B(n43338), .Y(n45966) );
  NAND2X1 U48096 ( .A(n2643), .B(n43365), .Y(n45965) );
  NAND2X1 U48097 ( .A(n45966), .B(n45965), .Y(n45967) );
  NOR2X1 U48098 ( .A(n45968), .B(n45967), .Y(n45969) );
  NAND2X1 U48099 ( .A(n45970), .B(n45969), .Y(n45971) );
  NOR2X1 U48100 ( .A(n45972), .B(n45971), .Y(n46003) );
  NAND2X1 U48101 ( .A(n2640), .B(n43044), .Y(n45974) );
  NAND2X1 U48102 ( .A(n2646), .B(n43047), .Y(n45973) );
  NAND2X1 U48103 ( .A(n45974), .B(n45973), .Y(n45978) );
  NAND2X1 U48104 ( .A(n2638), .B(n43049), .Y(n45976) );
  NAND2X1 U48105 ( .A(n2623), .B(n43051), .Y(n45975) );
  NAND2X1 U48106 ( .A(n45976), .B(n45975), .Y(n45977) );
  NOR2X1 U48107 ( .A(n45978), .B(n45977), .Y(n45985) );
  INVX1 U48108 ( .A(n2632), .Y(n45979) );
  NOR2X1 U48109 ( .A(n43370), .B(n45979), .Y(n45983) );
  NAND2X1 U48110 ( .A(n2625), .B(n43054), .Y(n45981) );
  NAND2X1 U48111 ( .A(n2648), .B(n43057), .Y(n45980) );
  NAND2X1 U48112 ( .A(n45981), .B(n45980), .Y(n45982) );
  NOR2X1 U48113 ( .A(n45983), .B(n45982), .Y(n45984) );
  NAND2X1 U48114 ( .A(n45985), .B(n45984), .Y(n46001) );
  NAND2X1 U48115 ( .A(n2644), .B(n43060), .Y(n45987) );
  NAND2X1 U48116 ( .A(n2642), .B(n39132), .Y(n45986) );
  NAND2X1 U48117 ( .A(n45987), .B(n45986), .Y(n45991) );
  NAND2X1 U48118 ( .A(n2634), .B(n43063), .Y(n45989) );
  NAND2X1 U48119 ( .A(n2626), .B(n43067), .Y(n45988) );
  NAND2X1 U48120 ( .A(n45989), .B(n45988), .Y(n45990) );
  NOR2X1 U48121 ( .A(n45991), .B(n45990), .Y(n45999) );
  NAND2X1 U48122 ( .A(n2630), .B(n43372), .Y(n45993) );
  NAND2X1 U48123 ( .A(n2636), .B(n43350), .Y(n45992) );
  NAND2X1 U48124 ( .A(n45993), .B(n45992), .Y(n45997) );
  NAND2X1 U48125 ( .A(n2628), .B(n43070), .Y(n45995) );
  NAND2X1 U48126 ( .A(n2621), .B(n43071), .Y(n45994) );
  NAND2X1 U48127 ( .A(n45995), .B(n45994), .Y(n45996) );
  NOR2X1 U48128 ( .A(n45997), .B(n45996), .Y(n45998) );
  NAND2X1 U48129 ( .A(n45999), .B(n45998), .Y(n46000) );
  NOR2X1 U48130 ( .A(n46001), .B(n46000), .Y(n46002) );
  NAND2X1 U48131 ( .A(n46003), .B(n46002), .Y(n46004) );
  NAND2X1 U48132 ( .A(n2642), .B(n46309), .Y(n46005) );
  OR2X1 U48133 ( .A(n46006), .B(n46005), .Y(n46012) );
  INVX1 U48134 ( .A(n40685), .Y(n46009) );
  NOR2X1 U48135 ( .A(n46009), .B(n46008), .Y(n46010) );
  NAND2X1 U48136 ( .A(n46010), .B(n42704), .Y(n46011) );
  NAND2X1 U48137 ( .A(n46012), .B(n46011), .Y(n46016) );
  NAND2X1 U48138 ( .A(n2634), .B(n40035), .Y(n46013) );
  NOR2X1 U48139 ( .A(n46016), .B(n46015), .Y(n59887) );
  INVX1 U48140 ( .A(n46236), .Y(n46017) );
  NAND2X1 U48141 ( .A(n2644), .B(n46017), .Y(n46018) );
  NOR2X1 U48142 ( .A(n46018), .B(n46394), .Y(n46022) );
  NOR2X1 U48143 ( .A(n46020), .B(n46394), .Y(n46021) );
  NOR2X1 U48144 ( .A(n46022), .B(n46021), .Y(n46027) );
  INVX1 U48145 ( .A(n40685), .Y(n46024) );
  OR2X1 U48146 ( .A(n46235), .B(n57608), .Y(n46023) );
  NOR2X1 U48147 ( .A(n46024), .B(n46023), .Y(n46025) );
  NAND2X1 U48148 ( .A(n2641), .B(n46025), .Y(n46026) );
  NAND2X1 U48149 ( .A(n46027), .B(n46026), .Y(n46069) );
  NAND2X1 U48150 ( .A(n2640), .B(n42678), .Y(n46029) );
  NAND2X1 U48151 ( .A(n46029), .B(n46028), .Y(n46040) );
  OR2X1 U48152 ( .A(n40507), .B(n40534), .Y(n46030) );
  NOR2X1 U48153 ( .A(n36800), .B(n46030), .Y(n46034) );
  OR2X1 U48154 ( .A(n40510), .B(n39196), .Y(n46031) );
  NOR2X1 U48155 ( .A(n46032), .B(n46031), .Y(n46033) );
  NOR2X1 U48156 ( .A(n46034), .B(n46033), .Y(n46038) );
  NOR2X1 U48157 ( .A(n46036), .B(n46035), .Y(n46037) );
  NAND2X1 U48158 ( .A(n46038), .B(n46037), .Y(n46039) );
  NOR2X1 U48159 ( .A(n46040), .B(n46039), .Y(n46044) );
  NOR2X1 U48160 ( .A(n46042), .B(n46041), .Y(n46043) );
  NOR2X1 U48161 ( .A(n38752), .B(n36817), .Y(n46048) );
  NAND2X1 U48162 ( .A(n45876), .B(n2645), .Y(n46046) );
  NAND2X1 U48163 ( .A(n46418), .B(n2643), .Y(n46045) );
  NAND2X1 U48164 ( .A(n46046), .B(n46045), .Y(n46047) );
  OR2X1 U48165 ( .A(n46048), .B(n46047), .Y(n46059) );
  INVX1 U48166 ( .A(n42867), .Y(n46049) );
  NAND2X1 U48167 ( .A(n2635), .B(n42676), .Y(n46050) );
  NOR2X1 U48168 ( .A(n36608), .B(n46050), .Y(n46051) );
  NAND2X1 U48169 ( .A(n2637), .B(n42676), .Y(n46053) );
  NOR2X1 U48170 ( .A(n38821), .B(n46053), .Y(n46057) );
  INVX1 U48171 ( .A(n42863), .Y(n46054) );
  NAND2X1 U48172 ( .A(n2620), .B(n36759), .Y(n46055) );
  NOR2X1 U48173 ( .A(n42875), .B(n46055), .Y(n46056) );
  NOR2X1 U48174 ( .A(n46059), .B(n46058), .Y(n46064) );
  OR2X1 U48175 ( .A(n39809), .B(n42700), .Y(n46060) );
  NOR2X1 U48176 ( .A(n36868), .B(n46060), .Y(n46062) );
  NOR2X1 U48177 ( .A(n46062), .B(n46061), .Y(n46063) );
  NAND2X1 U48178 ( .A(n46064), .B(n46063), .Y(n46065) );
  NAND2X1 U48179 ( .A(n42884), .B(n46065), .Y(n46066) );
  NAND2X1 U48180 ( .A(n46067), .B(n46066), .Y(n46068) );
  NOR2X1 U48181 ( .A(n46069), .B(n46068), .Y(n59886) );
  NOR2X1 U48182 ( .A(n46372), .B(n37022), .Y(n46071) );
  NOR2X1 U48183 ( .A(n38473), .B(n46235), .Y(n46070) );
  NAND2X1 U48184 ( .A(n46071), .B(n46070), .Y(n46075) );
  NAND2X1 U48185 ( .A(n46404), .B(n45610), .Y(n46072) );
  NOR2X1 U48186 ( .A(n46024), .B(n46072), .Y(n46073) );
  NAND2X1 U48187 ( .A(n46073), .B(n2633), .Y(n46074) );
  NAND2X1 U48188 ( .A(n46075), .B(n46074), .Y(n46082) );
  NOR2X1 U48189 ( .A(n42645), .B(n43209), .Y(n46078) );
  NAND2X1 U48190 ( .A(n46009), .B(n46367), .Y(n46076) );
  NOR2X1 U48191 ( .A(n43204), .B(n46076), .Y(n46077) );
  NOR2X1 U48192 ( .A(n46078), .B(n46077), .Y(n46080) );
  NAND2X1 U48193 ( .A(n46395), .B(n1820), .Y(n46079) );
  NAND2X1 U48194 ( .A(n46080), .B(n46079), .Y(n46081) );
  NAND2X1 U48195 ( .A(n2622), .B(n38824), .Y(n46083) );
  NOR2X1 U48196 ( .A(n42782), .B(n46083), .Y(n46089) );
  NOR2X1 U48197 ( .A(n38823), .B(n36846), .Y(n46084) );
  NAND2X1 U48198 ( .A(n46084), .B(n42770), .Y(n46087) );
  NOR2X1 U48199 ( .A(n36608), .B(n36852), .Y(n46085) );
  NAND2X1 U48200 ( .A(n46085), .B(n42771), .Y(n46086) );
  NAND2X1 U48201 ( .A(n46087), .B(n46086), .Y(n46088) );
  NOR2X1 U48202 ( .A(n46089), .B(n46088), .Y(n46090) );
  NOR2X1 U48203 ( .A(n46090), .B(n42885), .Y(n46092) );
  INVX1 U48204 ( .A(n46207), .Y(n46736) );
  NAND2X1 U48205 ( .A(n45707), .B(n46736), .Y(n46312) );
  NOR2X1 U48206 ( .A(n46312), .B(n37108), .Y(n46091) );
  NAND2X1 U48207 ( .A(n42221), .B(n40253), .Y(n70671) );
  NAND2X1 U48208 ( .A(n44006), .B(n43486), .Y(n57680) );
  INVX1 U48209 ( .A(mem_d_data_rd_i[25]), .Y(n46093) );
  NAND2X1 U48210 ( .A(n40935), .B(n46093), .Y(n46094) );
  NOR2X1 U48211 ( .A(n43454), .B(n43199), .Y(n46096) );
  NOR2X1 U48212 ( .A(n43022), .B(n43202), .Y(n46095) );
  NAND2X1 U48213 ( .A(n2847), .B(n43362), .Y(n46098) );
  NAND2X1 U48214 ( .A(n2822), .B(n38413), .Y(n46097) );
  NAND2X1 U48215 ( .A(n46098), .B(n46097), .Y(n46102) );
  NAND2X1 U48216 ( .A(n2829), .B(n38402), .Y(n46100) );
  NAND2X1 U48217 ( .A(n2837), .B(n43027), .Y(n46099) );
  NAND2X1 U48218 ( .A(n46100), .B(n46099), .Y(n46101) );
  NOR2X1 U48219 ( .A(n46102), .B(n46101), .Y(n46110) );
  NAND2X1 U48220 ( .A(n2819), .B(n43030), .Y(n46104) );
  NAND2X1 U48221 ( .A(n2824), .B(n43033), .Y(n46103) );
  NAND2X1 U48222 ( .A(n46104), .B(n46103), .Y(n46108) );
  NAND2X1 U48223 ( .A(n2839), .B(n43036), .Y(n46106) );
  NAND2X1 U48224 ( .A(n2831), .B(n43351), .Y(n46105) );
  NAND2X1 U48225 ( .A(n46106), .B(n46105), .Y(n46107) );
  NOR2X1 U48226 ( .A(n46108), .B(n46107), .Y(n46109) );
  NAND2X1 U48227 ( .A(n46110), .B(n46109), .Y(n46126) );
  NAND2X1 U48228 ( .A(n2835), .B(n43354), .Y(n46112) );
  NAND2X1 U48229 ( .A(n2833), .B(n43039), .Y(n46111) );
  NAND2X1 U48230 ( .A(n46112), .B(n46111), .Y(n46116) );
  NAND2X1 U48231 ( .A(n1810), .B(n39808), .Y(n46114) );
  NAND2X1 U48232 ( .A(n2841), .B(n43042), .Y(n46113) );
  NAND2X1 U48233 ( .A(n46114), .B(n46113), .Y(n46115) );
  NOR2X1 U48234 ( .A(n46116), .B(n46115), .Y(n46124) );
  NAND2X1 U48235 ( .A(n2845), .B(n38390), .Y(n46118) );
  NAND2X1 U48236 ( .A(n2820), .B(n43345), .Y(n46117) );
  NAND2X1 U48237 ( .A(n46118), .B(n46117), .Y(n46122) );
  NAND2X1 U48238 ( .A(n2827), .B(n43338), .Y(n46120) );
  NAND2X1 U48239 ( .A(n2843), .B(n43365), .Y(n46119) );
  NAND2X1 U48240 ( .A(n46120), .B(n46119), .Y(n46121) );
  NOR2X1 U48241 ( .A(n46122), .B(n46121), .Y(n46123) );
  NAND2X1 U48242 ( .A(n46124), .B(n46123), .Y(n46125) );
  NOR2X1 U48243 ( .A(n46126), .B(n46125), .Y(n46156) );
  NAND2X1 U48244 ( .A(n2840), .B(n43044), .Y(n46128) );
  NAND2X1 U48245 ( .A(n2846), .B(n43047), .Y(n46127) );
  NAND2X1 U48246 ( .A(n46128), .B(n46127), .Y(n46132) );
  NAND2X1 U48247 ( .A(n2838), .B(n43049), .Y(n46130) );
  NAND2X1 U48248 ( .A(n2823), .B(n43052), .Y(n46129) );
  NAND2X1 U48249 ( .A(n46130), .B(n46129), .Y(n46131) );
  NOR2X1 U48250 ( .A(n46132), .B(n46131), .Y(n46138) );
  NOR2X1 U48251 ( .A(n43371), .B(n37322), .Y(n46136) );
  NAND2X1 U48252 ( .A(n2825), .B(n43054), .Y(n46134) );
  NAND2X1 U48253 ( .A(n2848), .B(n43057), .Y(n46133) );
  NAND2X1 U48254 ( .A(n46134), .B(n46133), .Y(n46135) );
  NOR2X1 U48255 ( .A(n46136), .B(n46135), .Y(n46137) );
  NAND2X1 U48256 ( .A(n46138), .B(n46137), .Y(n46154) );
  NAND2X1 U48257 ( .A(n2844), .B(n43061), .Y(n46140) );
  NAND2X1 U48258 ( .A(n2842), .B(n39139), .Y(n46139) );
  NAND2X1 U48259 ( .A(n46140), .B(n46139), .Y(n46144) );
  NAND2X1 U48260 ( .A(n2834), .B(n43063), .Y(n46142) );
  NAND2X1 U48261 ( .A(n2826), .B(n43067), .Y(n46141) );
  NAND2X1 U48262 ( .A(n46142), .B(n46141), .Y(n46143) );
  NOR2X1 U48263 ( .A(n46144), .B(n46143), .Y(n46152) );
  NAND2X1 U48264 ( .A(n2830), .B(n43372), .Y(n46146) );
  NAND2X1 U48265 ( .A(n2836), .B(n43349), .Y(n46145) );
  NAND2X1 U48266 ( .A(n46146), .B(n46145), .Y(n46150) );
  NAND2X1 U48267 ( .A(n2828), .B(n43069), .Y(n46148) );
  NAND2X1 U48268 ( .A(n2821), .B(n43072), .Y(n46147) );
  NAND2X1 U48269 ( .A(n46148), .B(n46147), .Y(n46149) );
  NOR2X1 U48270 ( .A(n46150), .B(n46149), .Y(n46151) );
  NAND2X1 U48271 ( .A(n46152), .B(n46151), .Y(n46153) );
  NOR2X1 U48272 ( .A(n46154), .B(n46153), .Y(n46155) );
  NAND2X1 U48273 ( .A(n46156), .B(n46155), .Y(n46157) );
  NAND2X1 U48274 ( .A(n2838), .B(n42625), .Y(n46158) );
  NAND2X1 U48275 ( .A(n46159), .B(n46158), .Y(n46164) );
  INVX1 U48276 ( .A(n38213), .Y(n46160) );
  NAND2X1 U48277 ( .A(n2846), .B(n46160), .Y(n46161) );
  NAND2X1 U48278 ( .A(n46162), .B(n46161), .Y(n46163) );
  NOR2X1 U48279 ( .A(n46164), .B(n46163), .Y(n46173) );
  NAND2X1 U48280 ( .A(n2829), .B(n38740), .Y(n46166) );
  NAND2X1 U48281 ( .A(n2837), .B(n40424), .Y(n46165) );
  NAND2X1 U48282 ( .A(n46166), .B(n46165), .Y(n46171) );
  NOR2X1 U48283 ( .A(n40509), .B(n38821), .Y(n46167) );
  NAND2X1 U48284 ( .A(n2845), .B(n46167), .Y(n46168) );
  NAND2X1 U48285 ( .A(n46169), .B(n46168), .Y(n46170) );
  NOR2X1 U48286 ( .A(n46171), .B(n46170), .Y(n46172) );
  NAND2X1 U48287 ( .A(n46173), .B(n46172), .Y(n46204) );
  INVX1 U48288 ( .A(n49610), .Y(n46174) );
  NAND2X1 U48289 ( .A(n2827), .B(n46174), .Y(n46176) );
  NAND2X1 U48290 ( .A(n2820), .B(n38710), .Y(n46175) );
  NAND2X1 U48291 ( .A(n46176), .B(n46175), .Y(n46182) );
  INVX1 U48292 ( .A(n49605), .Y(n46177) );
  NAND2X1 U48293 ( .A(n2835), .B(n57615), .Y(n46180) );
  NOR2X1 U48294 ( .A(n40510), .B(n36608), .Y(n46178) );
  NAND2X1 U48295 ( .A(n2843), .B(n46178), .Y(n46179) );
  NAND2X1 U48296 ( .A(n46180), .B(n46179), .Y(n46181) );
  NOR2X1 U48297 ( .A(n46182), .B(n46181), .Y(n46202) );
  INVX1 U48298 ( .A(n2832), .Y(n46184) );
  NOR2X1 U48299 ( .A(n46184), .B(n45651), .Y(n46186) );
  NOR2X1 U48300 ( .A(n42891), .B(n36830), .Y(n46185) );
  NOR2X1 U48301 ( .A(n46186), .B(n46185), .Y(n46190) );
  NOR2X1 U48302 ( .A(n42684), .B(n36833), .Y(n46188) );
  NOR2X1 U48303 ( .A(n46188), .B(n46187), .Y(n46189) );
  NAND2X1 U48304 ( .A(n46190), .B(n46189), .Y(n46200) );
  NOR2X1 U48305 ( .A(n42646), .B(n36831), .Y(n46193) );
  OR2X1 U48306 ( .A(n40509), .B(n42695), .Y(n46191) );
  NOR2X1 U48307 ( .A(n36829), .B(n46191), .Y(n46192) );
  NOR2X1 U48308 ( .A(n46193), .B(n46192), .Y(n46198) );
  NOR2X1 U48309 ( .A(n40328), .B(n42700), .Y(n46196) );
  OR2X1 U48310 ( .A(n42765), .B(n42700), .Y(n46194) );
  NOR2X1 U48311 ( .A(n36835), .B(n46194), .Y(n46195) );
  NOR2X1 U48312 ( .A(n46196), .B(n46195), .Y(n46197) );
  NAND2X1 U48313 ( .A(n46198), .B(n46197), .Y(n46199) );
  NOR2X1 U48314 ( .A(n46200), .B(n46199), .Y(n46201) );
  NAND2X1 U48315 ( .A(n46202), .B(n46201), .Y(n46203) );
  NOR2X1 U48316 ( .A(n46204), .B(n46203), .Y(n46205) );
  NOR2X1 U48317 ( .A(n46205), .B(n42886), .Y(n46215) );
  NOR2X1 U48318 ( .A(n43199), .B(n42898), .Y(n46213) );
  NOR2X1 U48319 ( .A(n46206), .B(n37017), .Y(n46209) );
  NOR2X1 U48320 ( .A(n46207), .B(n37018), .Y(n46208) );
  NOR2X1 U48321 ( .A(n46209), .B(n46208), .Y(n46211) );
  NAND2X1 U48322 ( .A(n42692), .B(n40152), .Y(n46210) );
  NOR2X1 U48323 ( .A(n46211), .B(n46210), .Y(n46212) );
  NAND2X1 U48324 ( .A(n38604), .B(n46906), .Y(n46382) );
  NOR2X1 U48325 ( .A(n46215), .B(n46214), .Y(n59224) );
  NOR2X1 U48326 ( .A(n49715), .B(n43203), .Y(n46221) );
  NAND2X1 U48327 ( .A(n2834), .B(n46049), .Y(n46217) );
  NOR2X1 U48328 ( .A(n38464), .B(n46217), .Y(n46218) );
  NAND2X1 U48329 ( .A(n46218), .B(n38441), .Y(n46219) );
  NOR2X1 U48330 ( .A(n46526), .B(n46219), .Y(n46220) );
  NOR2X1 U48331 ( .A(n46221), .B(n46220), .Y(n46224) );
  NOR2X1 U48332 ( .A(n57608), .B(n46210), .Y(n46222) );
  NAND2X1 U48333 ( .A(n46222), .B(n2841), .Y(n46223) );
  NAND2X1 U48334 ( .A(n46224), .B(n46223), .Y(n46229) );
  INVX1 U48335 ( .A(n49630), .Y(n49719) );
  NOR2X1 U48336 ( .A(n46577), .B(n46210), .Y(n46225) );
  NAND2X1 U48337 ( .A(n46225), .B(n2836), .Y(n46226) );
  NAND2X1 U48338 ( .A(n46227), .B(n46226), .Y(n46228) );
  NOR2X1 U48339 ( .A(n46228), .B(n46229), .Y(n46243) );
  NOR2X1 U48340 ( .A(n46372), .B(n45681), .Y(n46230) );
  NAND2X1 U48341 ( .A(n46230), .B(n2826), .Y(n46234) );
  NOR2X1 U48342 ( .A(n46231), .B(n46394), .Y(n46232) );
  NAND2X1 U48343 ( .A(n46232), .B(n2821), .Y(n46233) );
  NAND2X1 U48344 ( .A(n46234), .B(n46233), .Y(n46241) );
  NAND2X1 U48345 ( .A(n40531), .B(n2828), .Y(n46239) );
  NOR2X1 U48346 ( .A(n46236), .B(n37071), .Y(n46237) );
  NAND2X1 U48347 ( .A(n46237), .B(n42146), .Y(n46238) );
  NAND2X1 U48348 ( .A(n46238), .B(n46239), .Y(n46240) );
  NOR2X1 U48349 ( .A(n46241), .B(n46240), .Y(n46242) );
  NAND2X1 U48350 ( .A(n59224), .B(n42347), .Y(n70371) );
  NAND2X1 U48351 ( .A(n43996), .B(n43484), .Y(n57717) );
  INVX1 U48352 ( .A(mem_d_data_rd_i[24]), .Y(n46244) );
  NAND2X1 U48353 ( .A(n40935), .B(n46244), .Y(n46245) );
  NOR2X1 U48354 ( .A(n43454), .B(n43194), .Y(n46247) );
  NOR2X1 U48355 ( .A(n43022), .B(n43197), .Y(n46246) );
  NAND2X1 U48356 ( .A(n2880), .B(n43362), .Y(n46249) );
  NAND2X1 U48357 ( .A(n2855), .B(n38413), .Y(n46248) );
  NAND2X1 U48358 ( .A(n46249), .B(n46248), .Y(n46253) );
  NAND2X1 U48359 ( .A(n2862), .B(n38401), .Y(n46251) );
  NAND2X1 U48360 ( .A(n2870), .B(n43027), .Y(n46250) );
  NAND2X1 U48361 ( .A(n46251), .B(n46250), .Y(n46252) );
  NOR2X1 U48362 ( .A(n46253), .B(n46252), .Y(n46261) );
  NAND2X1 U48363 ( .A(n2852), .B(n43030), .Y(n46255) );
  NAND2X1 U48364 ( .A(n2857), .B(n43032), .Y(n46254) );
  NAND2X1 U48365 ( .A(n46255), .B(n46254), .Y(n46259) );
  NAND2X1 U48366 ( .A(n2872), .B(n43036), .Y(n46257) );
  NAND2X1 U48367 ( .A(n2864), .B(n43352), .Y(n46256) );
  NAND2X1 U48368 ( .A(n46257), .B(n46256), .Y(n46258) );
  NOR2X1 U48369 ( .A(n46259), .B(n46258), .Y(n46260) );
  NAND2X1 U48370 ( .A(n46261), .B(n46260), .Y(n46277) );
  NAND2X1 U48371 ( .A(n2868), .B(n43356), .Y(n46263) );
  NAND2X1 U48372 ( .A(n2866), .B(n43039), .Y(n46262) );
  NAND2X1 U48373 ( .A(n46263), .B(n46262), .Y(n46267) );
  NAND2X1 U48374 ( .A(n1809), .B(n39808), .Y(n46265) );
  NAND2X1 U48375 ( .A(n2874), .B(n43042), .Y(n46264) );
  NAND2X1 U48376 ( .A(n46265), .B(n46264), .Y(n46266) );
  NOR2X1 U48377 ( .A(n46267), .B(n46266), .Y(n46275) );
  NAND2X1 U48378 ( .A(n2878), .B(n38389), .Y(n46269) );
  NAND2X1 U48379 ( .A(n2853), .B(n43346), .Y(n46268) );
  NAND2X1 U48380 ( .A(n46269), .B(n46268), .Y(n46273) );
  NAND2X1 U48381 ( .A(n2860), .B(n43339), .Y(n46271) );
  NAND2X1 U48382 ( .A(n2876), .B(n43366), .Y(n46270) );
  NAND2X1 U48383 ( .A(n46271), .B(n46270), .Y(n46272) );
  NOR2X1 U48384 ( .A(n46273), .B(n46272), .Y(n46274) );
  NAND2X1 U48385 ( .A(n46275), .B(n46274), .Y(n46276) );
  NOR2X1 U48386 ( .A(n46277), .B(n46276), .Y(n46307) );
  NAND2X1 U48387 ( .A(n2873), .B(n43044), .Y(n46279) );
  NAND2X1 U48388 ( .A(n2879), .B(n43047), .Y(n46278) );
  NAND2X1 U48389 ( .A(n46279), .B(n46278), .Y(n46283) );
  NAND2X1 U48390 ( .A(n2871), .B(n43049), .Y(n46281) );
  NAND2X1 U48391 ( .A(n2856), .B(n43051), .Y(n46280) );
  NAND2X1 U48392 ( .A(n46281), .B(n46280), .Y(n46282) );
  NOR2X1 U48393 ( .A(n46283), .B(n46282), .Y(n46289) );
  NOR2X1 U48394 ( .A(n43370), .B(n37321), .Y(n46287) );
  NAND2X1 U48395 ( .A(n2858), .B(n43054), .Y(n46285) );
  NAND2X1 U48396 ( .A(n2881), .B(n43057), .Y(n46284) );
  NAND2X1 U48397 ( .A(n46285), .B(n46284), .Y(n46286) );
  NOR2X1 U48398 ( .A(n46287), .B(n46286), .Y(n46288) );
  NAND2X1 U48399 ( .A(n46289), .B(n46288), .Y(n46305) );
  NAND2X1 U48400 ( .A(n2877), .B(n43060), .Y(n46291) );
  NAND2X1 U48401 ( .A(n2875), .B(n39139), .Y(n46290) );
  NAND2X1 U48402 ( .A(n46291), .B(n46290), .Y(n46295) );
  NAND2X1 U48403 ( .A(n2867), .B(n43063), .Y(n46293) );
  NAND2X1 U48404 ( .A(n2859), .B(n43067), .Y(n46292) );
  NAND2X1 U48405 ( .A(n46293), .B(n46292), .Y(n46294) );
  NOR2X1 U48406 ( .A(n46295), .B(n46294), .Y(n46303) );
  NAND2X1 U48407 ( .A(n2863), .B(n38528), .Y(n46297) );
  NAND2X1 U48408 ( .A(n2869), .B(n43350), .Y(n46296) );
  NAND2X1 U48409 ( .A(n46297), .B(n46296), .Y(n46301) );
  NAND2X1 U48410 ( .A(n2861), .B(n43070), .Y(n46299) );
  NAND2X1 U48411 ( .A(n2854), .B(n43071), .Y(n46298) );
  NAND2X1 U48412 ( .A(n46299), .B(n46298), .Y(n46300) );
  NOR2X1 U48413 ( .A(n46301), .B(n46300), .Y(n46302) );
  NAND2X1 U48414 ( .A(n46303), .B(n46302), .Y(n46304) );
  NOR2X1 U48415 ( .A(n46305), .B(n46304), .Y(n46306) );
  NAND2X1 U48416 ( .A(n46307), .B(n46306), .Y(n46308) );
  NAND2X1 U48417 ( .A(n43988), .B(n43995), .Y(n57713) );
  INVX1 U48418 ( .A(n57713), .Y(n46392) );
  NAND2X1 U48419 ( .A(n46572), .B(n2867), .Y(n46311) );
  NAND2X1 U48420 ( .A(n2875), .B(n40521), .Y(n46310) );
  NAND2X1 U48421 ( .A(n46311), .B(n46310), .Y(n46316) );
  NAND2X1 U48422 ( .A(n46314), .B(n46313), .Y(n46315) );
  NOR2X1 U48423 ( .A(n46316), .B(n46315), .Y(n46363) );
  NOR2X1 U48424 ( .A(n40427), .B(n36985), .Y(n46318) );
  NOR2X1 U48425 ( .A(n42776), .B(n37001), .Y(n46317) );
  NOR2X1 U48426 ( .A(n46318), .B(n46317), .Y(n46322) );
  NOR2X1 U48427 ( .A(n39654), .B(n36997), .Y(n46320) );
  NOR2X1 U48428 ( .A(n49604), .B(n37012), .Y(n46319) );
  NOR2X1 U48429 ( .A(n46320), .B(n46319), .Y(n46321) );
  NAND2X1 U48430 ( .A(n46322), .B(n46321), .Y(n46340) );
  NOR2X1 U48431 ( .A(n45199), .B(n38822), .Y(n46323) );
  NAND2X1 U48432 ( .A(n46323), .B(n2855), .Y(n46325) );
  NAND2X1 U48433 ( .A(n49577), .B(n2879), .Y(n46324) );
  NAND2X1 U48434 ( .A(n46325), .B(n46324), .Y(n46330) );
  NAND2X1 U48435 ( .A(n45472), .B(n2858), .Y(n46328) );
  NAND2X1 U48436 ( .A(n45475), .B(n2865), .Y(n46327) );
  NAND2X1 U48437 ( .A(n46328), .B(n46327), .Y(n46329) );
  NOR2X1 U48438 ( .A(n46330), .B(n46329), .Y(n46338) );
  NOR2X1 U48439 ( .A(n42628), .B(n37010), .Y(n46336) );
  NOR2X1 U48440 ( .A(n42768), .B(n36825), .Y(n46331) );
  NAND2X1 U48441 ( .A(n46331), .B(n38609), .Y(n46334) );
  NOR2X1 U48442 ( .A(n42866), .B(n36826), .Y(n46332) );
  NAND2X1 U48443 ( .A(n46332), .B(n38492), .Y(n46333) );
  NAND2X1 U48444 ( .A(n46334), .B(n46333), .Y(n46335) );
  NOR2X1 U48445 ( .A(n46336), .B(n46335), .Y(n46337) );
  NAND2X1 U48446 ( .A(n46338), .B(n46337), .Y(n46339) );
  NOR2X1 U48447 ( .A(n46340), .B(n46339), .Y(n46361) );
  NOR2X1 U48448 ( .A(n49599), .B(n36957), .Y(n46343) );
  NOR2X1 U48449 ( .A(n36975), .B(n42646), .Y(n46342) );
  NOR2X1 U48450 ( .A(n46343), .B(n46342), .Y(n46347) );
  NOR2X1 U48451 ( .A(n42623), .B(n36980), .Y(n46345) );
  NOR2X1 U48452 ( .A(n45244), .B(n36992), .Y(n46344) );
  NOR2X1 U48453 ( .A(n46345), .B(n46344), .Y(n46346) );
  NAND2X1 U48454 ( .A(n46347), .B(n46346), .Y(n46359) );
  NOR2X1 U48455 ( .A(n42684), .B(n36983), .Y(n46353) );
  NOR2X1 U48456 ( .A(n40507), .B(n36821), .Y(n46348) );
  NAND2X1 U48457 ( .A(n46348), .B(n38609), .Y(n46351) );
  NOR2X1 U48458 ( .A(n45199), .B(n36822), .Y(n46349) );
  NAND2X1 U48459 ( .A(n46349), .B(n38492), .Y(n46350) );
  NAND2X1 U48460 ( .A(n46351), .B(n46350), .Y(n46352) );
  NOR2X1 U48461 ( .A(n46353), .B(n46352), .Y(n46357) );
  NOR2X1 U48462 ( .A(n49677), .B(n36998), .Y(n46355) );
  NOR2X1 U48463 ( .A(n42905), .B(n37013), .Y(n46354) );
  NOR2X1 U48464 ( .A(n46355), .B(n46354), .Y(n46356) );
  NAND2X1 U48465 ( .A(n46357), .B(n46356), .Y(n46358) );
  NOR2X1 U48466 ( .A(n46359), .B(n46358), .Y(n46360) );
  NAND2X1 U48467 ( .A(n46363), .B(n46362), .Y(n46364) );
  NAND2X1 U48468 ( .A(n42692), .B(n38441), .Y(n46366) );
  NAND2X1 U48469 ( .A(n2874), .B(n46741), .Y(n46365) );
  NOR2X1 U48470 ( .A(n46366), .B(n46365), .Y(n46376) );
  NOR2X1 U48471 ( .A(n49715), .B(n43198), .Y(n46370) );
  NAND2X1 U48472 ( .A(n38473), .B(n46367), .Y(n46368) );
  NOR2X1 U48473 ( .A(n43194), .B(n46368), .Y(n46369) );
  NOR2X1 U48474 ( .A(n46370), .B(n46369), .Y(n46374) );
  NAND2X1 U48475 ( .A(n45610), .B(n45176), .Y(n46371) );
  NOR2X1 U48476 ( .A(n46372), .B(n46371), .Y(n49705) );
  NAND2X1 U48477 ( .A(n2859), .B(n49705), .Y(n46373) );
  NAND2X1 U48478 ( .A(n46374), .B(n46373), .Y(n46375) );
  NOR2X1 U48479 ( .A(n46376), .B(n46375), .Y(n46388) );
  NAND2X1 U48480 ( .A(n2869), .B(n40447), .Y(n46377) );
  NOR2X1 U48481 ( .A(n46726), .B(n46377), .Y(n46379) );
  NOR2X1 U48482 ( .A(n46379), .B(n46378), .Y(n46381) );
  NAND2X1 U48483 ( .A(n2854), .B(n40432), .Y(n46380) );
  NAND2X1 U48484 ( .A(n46381), .B(n46380), .Y(n46386) );
  NAND2X1 U48485 ( .A(n46384), .B(n46383), .Y(n46385) );
  NOR2X1 U48486 ( .A(n46386), .B(n46385), .Y(n46387) );
  NAND2X1 U48487 ( .A(n46388), .B(n46387), .Y(n46389) );
  NAND2X1 U48488 ( .A(n43996), .B(n43478), .Y(n46391) );
  NAND2X1 U48489 ( .A(n43988), .B(n38313), .Y(n46390) );
  NAND2X1 U48490 ( .A(n46391), .B(n46390), .Y(n57716) );
  NOR2X1 U48491 ( .A(n46392), .B(n57716), .Y(n46393) );
  NAND2X1 U48492 ( .A(n43477), .B(n43483), .Y(n57714) );
  NAND2X1 U48493 ( .A(n46393), .B(n57714), .Y(n49803) );
  NAND2X1 U48494 ( .A(n42146), .B(n40404), .Y(n49625) );
  NOR2X1 U48495 ( .A(n37111), .B(n40862), .Y(n46397) );
  NOR2X1 U48496 ( .A(n46575), .B(n46394), .Y(n46395) );
  NOR2X1 U48497 ( .A(n37107), .B(n49624), .Y(n46403) );
  INVX1 U48498 ( .A(mem_d_data_rd_i[23]), .Y(n46398) );
  NAND2X1 U48499 ( .A(n40935), .B(n46398), .Y(n46399) );
  NAND2X1 U48500 ( .A(n46399), .B(n42878), .Y(n53889) );
  NAND2X1 U48501 ( .A(writeback_exec_value_w[23]), .B(n37976), .Y(n46400) );
  NAND2X1 U48502 ( .A(n46401), .B(n46400), .Y(n46402) );
  NOR2X1 U48503 ( .A(n46403), .B(n46402), .Y(n46409) );
  NAND2X1 U48504 ( .A(n42705), .B(n40152), .Y(n46569) );
  NAND2X1 U48505 ( .A(n2467), .B(n46404), .Y(n46405) );
  NOR2X1 U48506 ( .A(n46569), .B(n46405), .Y(n46406) );
  NOR2X1 U48507 ( .A(n46407), .B(n46406), .Y(n46408) );
  NAND2X1 U48508 ( .A(n46409), .B(n46408), .Y(n59148) );
  NOR2X1 U48509 ( .A(n59149), .B(n59148), .Y(n46458) );
  NAND2X1 U48510 ( .A(n49705), .B(n2459), .Y(n46411) );
  NAND2X1 U48511 ( .A(n46411), .B(n46410), .Y(n46417) );
  NAND2X1 U48512 ( .A(n2462), .B(n40531), .Y(n46415) );
  NOR2X1 U48513 ( .A(n57608), .B(n37096), .Y(n46413) );
  NOR2X1 U48514 ( .A(n46024), .B(n46235), .Y(n46412) );
  NAND2X1 U48515 ( .A(n46413), .B(n45712), .Y(n46414) );
  NAND2X1 U48516 ( .A(n46415), .B(n46414), .Y(n46416) );
  NOR2X1 U48517 ( .A(n36938), .B(n49599), .Y(n46422) );
  INVX1 U48518 ( .A(n42894), .Y(n57621) );
  NAND2X1 U48519 ( .A(n2456), .B(n38844), .Y(n46420) );
  NOR2X1 U48520 ( .A(n40479), .B(n36600), .Y(n46418) );
  NAND2X1 U48521 ( .A(n46418), .B(n2477), .Y(n46419) );
  NAND2X1 U48522 ( .A(n46420), .B(n46419), .Y(n46421) );
  NOR2X1 U48523 ( .A(n46422), .B(n46421), .Y(n46426) );
  NOR2X1 U48524 ( .A(n49604), .B(n36952), .Y(n46424) );
  NOR2X1 U48525 ( .A(n42615), .B(n36968), .Y(n46423) );
  NOR2X1 U48526 ( .A(n46424), .B(n46423), .Y(n46425) );
  NAND2X1 U48527 ( .A(n46426), .B(n46425), .Y(n46436) );
  NOR2X1 U48528 ( .A(n42741), .B(n36955), .Y(n46430) );
  INVX1 U48529 ( .A(n42892), .Y(n49611) );
  NAND2X1 U48530 ( .A(n2460), .B(n36610), .Y(n46427) );
  NAND2X1 U48531 ( .A(n46428), .B(n46427), .Y(n46429) );
  NOR2X1 U48532 ( .A(n46430), .B(n46429), .Y(n46434) );
  NOR2X1 U48533 ( .A(n38712), .B(n36970), .Y(n46432) );
  NOR2X1 U48534 ( .A(n42776), .B(n36984), .Y(n46431) );
  NOR2X1 U48535 ( .A(n46432), .B(n46431), .Y(n46433) );
  NAND2X1 U48536 ( .A(n46434), .B(n46433), .Y(n46435) );
  NOR2X1 U48537 ( .A(n46436), .B(n46435), .Y(n46456) );
  NOR2X1 U48538 ( .A(n42858), .B(n36950), .Y(n46440) );
  NAND2X1 U48539 ( .A(n2474), .B(n42678), .Y(n46438) );
  NAND2X1 U48540 ( .A(n2458), .B(n40249), .Y(n46437) );
  NAND2X1 U48541 ( .A(n46438), .B(n46437), .Y(n46439) );
  NOR2X1 U48542 ( .A(n46440), .B(n46439), .Y(n46444) );
  NOR2X1 U48543 ( .A(n45244), .B(n36958), .Y(n46442) );
  NOR2X1 U48544 ( .A(n40427), .B(n36978), .Y(n46441) );
  NOR2X1 U48545 ( .A(n46442), .B(n46441), .Y(n46443) );
  NAND2X1 U48546 ( .A(n46444), .B(n46443), .Y(n46454) );
  NOR2X1 U48547 ( .A(n36946), .B(n42906), .Y(n46448) );
  NAND2X1 U48548 ( .A(n2457), .B(n49674), .Y(n46446) );
  NAND2X1 U48549 ( .A(n2472), .B(n42625), .Y(n46445) );
  NAND2X1 U48550 ( .A(n46446), .B(n46445), .Y(n46447) );
  NOR2X1 U48551 ( .A(n46448), .B(n46447), .Y(n46452) );
  NOR2X1 U48552 ( .A(n36951), .B(n42902), .Y(n46450) );
  NOR2X1 U48553 ( .A(n42622), .B(n36995), .Y(n46449) );
  NOR2X1 U48554 ( .A(n46450), .B(n46449), .Y(n46451) );
  NAND2X1 U48555 ( .A(n46452), .B(n46451), .Y(n46453) );
  NOR2X1 U48556 ( .A(n46454), .B(n46453), .Y(n46455) );
  NAND2X1 U48557 ( .A(n46456), .B(n46455), .Y(n46457) );
  INVX1 U48558 ( .A(n59147), .Y(n59120) );
  NAND2X1 U48559 ( .A(n46458), .B(n59120), .Y(n72803) );
  INVX1 U48560 ( .A(mem_d_data_rd_i[22]), .Y(n46459) );
  NAND2X1 U48561 ( .A(n40935), .B(n46459), .Y(n46460) );
  NAND2X1 U48562 ( .A(n46460), .B(n42876), .Y(n53762) );
  NOR2X1 U48563 ( .A(n43454), .B(n43182), .Y(n46462) );
  NOR2X1 U48564 ( .A(n43022), .B(n43185), .Y(n46461) );
  NAND2X1 U48565 ( .A(n2513), .B(n43362), .Y(n46464) );
  NAND2X1 U48566 ( .A(n2488), .B(n38411), .Y(n46463) );
  NAND2X1 U48567 ( .A(n46464), .B(n46463), .Y(n46468) );
  NAND2X1 U48568 ( .A(n2495), .B(n43344), .Y(n46466) );
  NAND2X1 U48569 ( .A(n2503), .B(n43027), .Y(n46465) );
  NAND2X1 U48570 ( .A(n46466), .B(n46465), .Y(n46467) );
  NOR2X1 U48571 ( .A(n46468), .B(n46467), .Y(n46476) );
  NAND2X1 U48572 ( .A(n2485), .B(n43030), .Y(n46470) );
  NAND2X1 U48573 ( .A(n2490), .B(n43032), .Y(n46469) );
  NAND2X1 U48574 ( .A(n46470), .B(n46469), .Y(n46474) );
  NAND2X1 U48575 ( .A(n2505), .B(n43036), .Y(n46472) );
  NAND2X1 U48576 ( .A(n2497), .B(n43351), .Y(n46471) );
  NAND2X1 U48577 ( .A(n46472), .B(n46471), .Y(n46473) );
  NOR2X1 U48578 ( .A(n46474), .B(n46473), .Y(n46475) );
  NAND2X1 U48579 ( .A(n46476), .B(n46475), .Y(n46492) );
  NAND2X1 U48580 ( .A(n2501), .B(n43354), .Y(n46478) );
  NAND2X1 U48581 ( .A(n2499), .B(n43039), .Y(n46477) );
  NAND2X1 U48582 ( .A(n46478), .B(n46477), .Y(n46482) );
  NAND2X1 U48583 ( .A(n1824), .B(n39808), .Y(n46480) );
  NAND2X1 U48584 ( .A(n2507), .B(n43042), .Y(n46479) );
  NAND2X1 U48585 ( .A(n46480), .B(n46479), .Y(n46481) );
  NOR2X1 U48586 ( .A(n46482), .B(n46481), .Y(n46490) );
  NAND2X1 U48587 ( .A(n2511), .B(n43360), .Y(n46484) );
  NAND2X1 U48588 ( .A(n2486), .B(n43345), .Y(n46483) );
  NAND2X1 U48589 ( .A(n46484), .B(n46483), .Y(n46488) );
  NAND2X1 U48590 ( .A(n2493), .B(n43338), .Y(n46486) );
  NAND2X1 U48591 ( .A(n2509), .B(n43365), .Y(n46485) );
  NAND2X1 U48592 ( .A(n46486), .B(n46485), .Y(n46487) );
  NOR2X1 U48593 ( .A(n46488), .B(n46487), .Y(n46489) );
  NAND2X1 U48594 ( .A(n46490), .B(n46489), .Y(n46491) );
  NOR2X1 U48595 ( .A(n46492), .B(n46491), .Y(n46522) );
  NAND2X1 U48596 ( .A(n2506), .B(n43044), .Y(n46494) );
  NAND2X1 U48597 ( .A(n2512), .B(n43047), .Y(n46493) );
  NAND2X1 U48598 ( .A(n46494), .B(n46493), .Y(n46498) );
  NAND2X1 U48599 ( .A(n2504), .B(n43049), .Y(n46496) );
  NAND2X1 U48600 ( .A(n2489), .B(n43051), .Y(n46495) );
  NAND2X1 U48601 ( .A(n46496), .B(n46495), .Y(n46497) );
  NOR2X1 U48602 ( .A(n46498), .B(n46497), .Y(n46504) );
  NOR2X1 U48603 ( .A(n43370), .B(n37317), .Y(n46502) );
  NAND2X1 U48604 ( .A(n2492), .B(n43054), .Y(n46500) );
  NAND2X1 U48605 ( .A(n2514), .B(n43057), .Y(n46499) );
  NAND2X1 U48606 ( .A(n46500), .B(n46499), .Y(n46501) );
  NOR2X1 U48607 ( .A(n46502), .B(n46501), .Y(n46503) );
  NAND2X1 U48608 ( .A(n46504), .B(n46503), .Y(n46520) );
  NAND2X1 U48609 ( .A(n2510), .B(n43060), .Y(n46506) );
  NAND2X1 U48610 ( .A(n2508), .B(n39137), .Y(n46505) );
  NAND2X1 U48611 ( .A(n46506), .B(n46505), .Y(n46510) );
  NAND2X1 U48612 ( .A(n2500), .B(n43063), .Y(n46508) );
  NAND2X1 U48613 ( .A(n2491), .B(n43067), .Y(n46507) );
  NAND2X1 U48614 ( .A(n46508), .B(n46507), .Y(n46509) );
  NOR2X1 U48615 ( .A(n46510), .B(n46509), .Y(n46518) );
  NAND2X1 U48616 ( .A(n2496), .B(n43372), .Y(n46512) );
  NAND2X1 U48617 ( .A(n2502), .B(n43350), .Y(n46511) );
  NAND2X1 U48618 ( .A(n46512), .B(n46511), .Y(n46516) );
  NAND2X1 U48619 ( .A(n2494), .B(n43070), .Y(n46514) );
  NAND2X1 U48620 ( .A(n2487), .B(n43071), .Y(n46513) );
  NAND2X1 U48621 ( .A(n46514), .B(n46513), .Y(n46515) );
  NOR2X1 U48622 ( .A(n46516), .B(n46515), .Y(n46517) );
  NAND2X1 U48623 ( .A(n46518), .B(n46517), .Y(n46519) );
  NOR2X1 U48624 ( .A(n46520), .B(n46519), .Y(n46521) );
  NAND2X1 U48625 ( .A(n46522), .B(n46521), .Y(n46523) );
  NOR2X1 U48626 ( .A(n43778), .B(n43945), .Y(n46654) );
  NAND2X1 U48627 ( .A(n2491), .B(n49705), .Y(n46525) );
  NAND2X1 U48628 ( .A(n2487), .B(n40432), .Y(n46524) );
  NAND2X1 U48629 ( .A(n46525), .B(n46524), .Y(n46530) );
  NAND2X1 U48630 ( .A(n2494), .B(n40531), .Y(n46528) );
  NAND2X1 U48631 ( .A(n42830), .B(n2507), .Y(n46527) );
  NAND2X1 U48632 ( .A(n46528), .B(n46527), .Y(n46529) );
  NAND2X1 U48633 ( .A(n2495), .B(n42779), .Y(n46532) );
  NAND2X1 U48634 ( .A(n2486), .B(n38708), .Y(n46531) );
  NAND2X1 U48635 ( .A(n46532), .B(n46531), .Y(n46536) );
  INVX1 U48636 ( .A(n42904), .Y(n57617) );
  NAND2X1 U48637 ( .A(n2511), .B(n42223), .Y(n46534) );
  INVX1 U48638 ( .A(n45640), .Y(n57619) );
  NAND2X1 U48639 ( .A(n2513), .B(n42147), .Y(n46533) );
  NAND2X1 U48640 ( .A(n46534), .B(n46533), .Y(n46535) );
  NOR2X1 U48641 ( .A(n46536), .B(n46535), .Y(n46540) );
  NOR2X1 U48642 ( .A(n42647), .B(n36989), .Y(n46538) );
  NOR2X1 U48643 ( .A(n42859), .B(n37002), .Y(n46537) );
  NOR2X1 U48644 ( .A(n46538), .B(n46537), .Y(n46539) );
  NAND2X1 U48645 ( .A(n46540), .B(n46539), .Y(n46548) );
  NOR2X1 U48646 ( .A(n49587), .B(n36996), .Y(n46542) );
  NOR2X1 U48647 ( .A(n49610), .B(n37005), .Y(n46541) );
  NOR2X1 U48648 ( .A(n46542), .B(n46541), .Y(n46546) );
  NOR2X1 U48649 ( .A(n42893), .B(n37011), .Y(n46543) );
  NOR2X1 U48650 ( .A(n46544), .B(n46543), .Y(n46545) );
  NAND2X1 U48651 ( .A(n46546), .B(n46545), .Y(n46547) );
  NOR2X1 U48652 ( .A(n46548), .B(n46547), .Y(n46567) );
  NAND2X1 U48653 ( .A(n2498), .B(n42821), .Y(n46550) );
  NAND2X1 U48654 ( .A(n2492), .B(n49611), .Y(n46549) );
  NAND2X1 U48655 ( .A(n46550), .B(n46549), .Y(n46553) );
  NAND2X1 U48656 ( .A(n2506), .B(n42678), .Y(n46551) );
  INVX1 U48657 ( .A(n49599), .Y(n57613) );
  NAND2X1 U48658 ( .A(n46551), .B(n42475), .Y(n46552) );
  NOR2X1 U48659 ( .A(n46553), .B(n46552), .Y(n46557) );
  NOR2X1 U48660 ( .A(n49604), .B(n37000), .Y(n46555) );
  NOR2X1 U48661 ( .A(n42616), .B(n37009), .Y(n46554) );
  NOR2X1 U48662 ( .A(n46555), .B(n46554), .Y(n46556) );
  NAND2X1 U48663 ( .A(n46557), .B(n46556), .Y(n46565) );
  NOR2X1 U48664 ( .A(n42628), .B(n37003), .Y(n46559) );
  NOR2X1 U48665 ( .A(n39654), .B(n37014), .Y(n46558) );
  NOR2X1 U48666 ( .A(n46559), .B(n46558), .Y(n46563) );
  NOR2X1 U48667 ( .A(n45244), .B(n37008), .Y(n46561) );
  NOR2X1 U48668 ( .A(n40428), .B(n37016), .Y(n46560) );
  NOR2X1 U48669 ( .A(n46561), .B(n46560), .Y(n46562) );
  NAND2X1 U48670 ( .A(n46563), .B(n46562), .Y(n46564) );
  NOR2X1 U48671 ( .A(n46565), .B(n46564), .Y(n46566) );
  NAND2X1 U48672 ( .A(n46567), .B(n46566), .Y(n46568) );
  NOR2X1 U48673 ( .A(n46570), .B(n46569), .Y(n46571) );
  NAND2X1 U48674 ( .A(n46571), .B(n2499), .Y(n46574) );
  NOR2X1 U48675 ( .A(n57605), .B(n45681), .Y(n46572) );
  NAND2X1 U48676 ( .A(n46572), .B(n2500), .Y(n46573) );
  NAND2X1 U48677 ( .A(n46574), .B(n46573), .Y(n46582) );
  NOR2X1 U48678 ( .A(n46575), .B(n37098), .Y(n46576) );
  NAND2X1 U48679 ( .A(n46576), .B(n38604), .Y(n46580) );
  NOR2X1 U48680 ( .A(n46577), .B(n46726), .Y(n46578) );
  NAND2X1 U48681 ( .A(n46578), .B(n2502), .Y(n46579) );
  NAND2X1 U48682 ( .A(n46580), .B(n46579), .Y(n46581) );
  NOR2X1 U48683 ( .A(n42908), .B(n37151), .Y(n46587) );
  NAND2X1 U48684 ( .A(writeback_exec_value_w[22]), .B(n37976), .Y(n46584) );
  NAND2X1 U48685 ( .A(n42838), .B(n36621), .Y(n72811) );
  NAND2X1 U48686 ( .A(n43796), .B(n43775), .Y(n46653) );
  NOR2X1 U48687 ( .A(n43454), .B(n43188), .Y(n46589) );
  NOR2X1 U48688 ( .A(n43022), .B(n43191), .Y(n46588) );
  NAND2X1 U48689 ( .A(n2481), .B(n43362), .Y(n46591) );
  NAND2X1 U48690 ( .A(n2456), .B(n38412), .Y(n46590) );
  NAND2X1 U48691 ( .A(n46591), .B(n46590), .Y(n46595) );
  NAND2X1 U48692 ( .A(n2463), .B(n43342), .Y(n46593) );
  NAND2X1 U48693 ( .A(n2471), .B(n43027), .Y(n46592) );
  NAND2X1 U48694 ( .A(n46593), .B(n46592), .Y(n46594) );
  NOR2X1 U48695 ( .A(n46595), .B(n46594), .Y(n46603) );
  NAND2X1 U48696 ( .A(n2453), .B(n43030), .Y(n46597) );
  NAND2X1 U48697 ( .A(n2458), .B(n43032), .Y(n46596) );
  NAND2X1 U48698 ( .A(n46597), .B(n46596), .Y(n46601) );
  NAND2X1 U48699 ( .A(n2473), .B(n43036), .Y(n46599) );
  NAND2X1 U48700 ( .A(n2465), .B(n43351), .Y(n46598) );
  NAND2X1 U48701 ( .A(n46599), .B(n46598), .Y(n46600) );
  NOR2X1 U48702 ( .A(n46601), .B(n46600), .Y(n46602) );
  NAND2X1 U48703 ( .A(n46603), .B(n46602), .Y(n46619) );
  NAND2X1 U48704 ( .A(n2469), .B(n43355), .Y(n46605) );
  NAND2X1 U48705 ( .A(n2467), .B(n43039), .Y(n46604) );
  NAND2X1 U48706 ( .A(n46605), .B(n46604), .Y(n46609) );
  NAND2X1 U48707 ( .A(n1825), .B(n39808), .Y(n46607) );
  NAND2X1 U48708 ( .A(n2475), .B(n43042), .Y(n46606) );
  NAND2X1 U48709 ( .A(n46607), .B(n46606), .Y(n46608) );
  NOR2X1 U48710 ( .A(n46609), .B(n46608), .Y(n46617) );
  NAND2X1 U48711 ( .A(n2479), .B(n43358), .Y(n46611) );
  NAND2X1 U48712 ( .A(n2454), .B(n43345), .Y(n46610) );
  NAND2X1 U48713 ( .A(n46611), .B(n46610), .Y(n46615) );
  NAND2X1 U48714 ( .A(n2461), .B(n43338), .Y(n46613) );
  NAND2X1 U48715 ( .A(n2477), .B(n43365), .Y(n46612) );
  NAND2X1 U48716 ( .A(n46613), .B(n46612), .Y(n46614) );
  NOR2X1 U48717 ( .A(n46615), .B(n46614), .Y(n46616) );
  NAND2X1 U48718 ( .A(n46617), .B(n46616), .Y(n46618) );
  NOR2X1 U48719 ( .A(n46619), .B(n46618), .Y(n46650) );
  NAND2X1 U48720 ( .A(n2474), .B(n43044), .Y(n46621) );
  NAND2X1 U48721 ( .A(n2480), .B(n43047), .Y(n46620) );
  NAND2X1 U48722 ( .A(n46621), .B(n46620), .Y(n46625) );
  NAND2X1 U48723 ( .A(n2472), .B(n43049), .Y(n46623) );
  NAND2X1 U48724 ( .A(n2457), .B(n43051), .Y(n46622) );
  NAND2X1 U48725 ( .A(n46623), .B(n46622), .Y(n46624) );
  NOR2X1 U48726 ( .A(n46625), .B(n46624), .Y(n46632) );
  NOR2X1 U48727 ( .A(n43371), .B(n46626), .Y(n46630) );
  NAND2X1 U48728 ( .A(n2460), .B(n43054), .Y(n46628) );
  NAND2X1 U48729 ( .A(n2482), .B(n43057), .Y(n46627) );
  NAND2X1 U48730 ( .A(n46628), .B(n46627), .Y(n46629) );
  NOR2X1 U48731 ( .A(n46630), .B(n46629), .Y(n46631) );
  NAND2X1 U48732 ( .A(n46632), .B(n46631), .Y(n46648) );
  NAND2X1 U48733 ( .A(n2478), .B(n43060), .Y(n46634) );
  NAND2X1 U48734 ( .A(n2476), .B(n39138), .Y(n46633) );
  NAND2X1 U48735 ( .A(n46634), .B(n46633), .Y(n46638) );
  NAND2X1 U48736 ( .A(n2468), .B(n43063), .Y(n46636) );
  NAND2X1 U48737 ( .A(n2459), .B(n43067), .Y(n46635) );
  NAND2X1 U48738 ( .A(n46636), .B(n46635), .Y(n46637) );
  NOR2X1 U48739 ( .A(n46638), .B(n46637), .Y(n46646) );
  NAND2X1 U48740 ( .A(n2464), .B(n43372), .Y(n46640) );
  NAND2X1 U48741 ( .A(n2470), .B(n43349), .Y(n46639) );
  NAND2X1 U48742 ( .A(n46640), .B(n46639), .Y(n46644) );
  NAND2X1 U48743 ( .A(n2462), .B(n43070), .Y(n46642) );
  NAND2X1 U48744 ( .A(n2455), .B(n43071), .Y(n46641) );
  NAND2X1 U48745 ( .A(n46642), .B(n46641), .Y(n46643) );
  NOR2X1 U48746 ( .A(n46644), .B(n46643), .Y(n46645) );
  NAND2X1 U48747 ( .A(n46646), .B(n46645), .Y(n46647) );
  NOR2X1 U48748 ( .A(n46648), .B(n46647), .Y(n46649) );
  NAND2X1 U48749 ( .A(n46650), .B(n46649), .Y(n46651) );
  NAND2X1 U48750 ( .A(n43949), .B(n43979), .Y(n46652) );
  NAND2X1 U48751 ( .A(n46653), .B(n46652), .Y(n57730) );
  NOR2X1 U48752 ( .A(n46654), .B(n57730), .Y(n46656) );
  NAND2X1 U48753 ( .A(n43978), .B(n43795), .Y(n46655) );
  NAND2X1 U48754 ( .A(n46656), .B(n46655), .Y(n49800) );
  NAND2X1 U48755 ( .A(n43949), .B(n43795), .Y(n46786) );
  INVX1 U48756 ( .A(mem_d_data_rd_i[21]), .Y(n73548) );
  NAND2X1 U48757 ( .A(n40935), .B(n73548), .Y(n46657) );
  NOR2X1 U48758 ( .A(n43454), .B(n43176), .Y(n46659) );
  NOR2X1 U48759 ( .A(n43022), .B(n43179), .Y(n46658) );
  NOR2X1 U48760 ( .A(n46659), .B(n46658), .Y(n46723) );
  NAND2X1 U48761 ( .A(n2579), .B(n43362), .Y(n46661) );
  NAND2X1 U48762 ( .A(n2554), .B(n38410), .Y(n46660) );
  NAND2X1 U48763 ( .A(n46661), .B(n46660), .Y(n46665) );
  NAND2X1 U48764 ( .A(n2561), .B(n43343), .Y(n46663) );
  NAND2X1 U48765 ( .A(n2569), .B(n43027), .Y(n46662) );
  NAND2X1 U48766 ( .A(n46663), .B(n46662), .Y(n46664) );
  NOR2X1 U48767 ( .A(n46665), .B(n46664), .Y(n46673) );
  NAND2X1 U48768 ( .A(n2551), .B(n43030), .Y(n46667) );
  NAND2X1 U48769 ( .A(n2556), .B(n43032), .Y(n46666) );
  NAND2X1 U48770 ( .A(n46667), .B(n46666), .Y(n46671) );
  NAND2X1 U48771 ( .A(n2571), .B(n43036), .Y(n46669) );
  NAND2X1 U48772 ( .A(n2563), .B(n43351), .Y(n46668) );
  NAND2X1 U48773 ( .A(n46669), .B(n46668), .Y(n46670) );
  NOR2X1 U48774 ( .A(n46671), .B(n46670), .Y(n46672) );
  NAND2X1 U48775 ( .A(n46673), .B(n46672), .Y(n46689) );
  NAND2X1 U48776 ( .A(n2567), .B(n43356), .Y(n46675) );
  NAND2X1 U48777 ( .A(n2565), .B(n43039), .Y(n46674) );
  NAND2X1 U48778 ( .A(n46675), .B(n46674), .Y(n46679) );
  NAND2X1 U48779 ( .A(n1822), .B(n39807), .Y(n46677) );
  NAND2X1 U48780 ( .A(n2573), .B(n43042), .Y(n46676) );
  NAND2X1 U48781 ( .A(n46677), .B(n46676), .Y(n46678) );
  NOR2X1 U48782 ( .A(n46679), .B(n46678), .Y(n46687) );
  NAND2X1 U48783 ( .A(n2577), .B(n43359), .Y(n46681) );
  NAND2X1 U48784 ( .A(n2552), .B(n43345), .Y(n46680) );
  NAND2X1 U48785 ( .A(n46681), .B(n46680), .Y(n46685) );
  NAND2X1 U48786 ( .A(n2559), .B(n43338), .Y(n46683) );
  NAND2X1 U48787 ( .A(n2575), .B(n43365), .Y(n46682) );
  NAND2X1 U48788 ( .A(n46683), .B(n46682), .Y(n46684) );
  NOR2X1 U48789 ( .A(n46685), .B(n46684), .Y(n46686) );
  NAND2X1 U48790 ( .A(n46687), .B(n46686), .Y(n46688) );
  NOR2X1 U48791 ( .A(n46689), .B(n46688), .Y(n46720) );
  NAND2X1 U48792 ( .A(n2572), .B(n43044), .Y(n46691) );
  NAND2X1 U48793 ( .A(n2578), .B(n43047), .Y(n46690) );
  NAND2X1 U48794 ( .A(n46691), .B(n46690), .Y(n46695) );
  NAND2X1 U48795 ( .A(n2570), .B(n43049), .Y(n46693) );
  NAND2X1 U48796 ( .A(n2555), .B(n43051), .Y(n46692) );
  NAND2X1 U48797 ( .A(n46693), .B(n46692), .Y(n46694) );
  NOR2X1 U48798 ( .A(n46695), .B(n46694), .Y(n46702) );
  NOR2X1 U48799 ( .A(n43371), .B(n46696), .Y(n46700) );
  NAND2X1 U48800 ( .A(n2558), .B(n43054), .Y(n46698) );
  NAND2X1 U48801 ( .A(n2580), .B(n43057), .Y(n46697) );
  NAND2X1 U48802 ( .A(n46698), .B(n46697), .Y(n46699) );
  NOR2X1 U48803 ( .A(n46700), .B(n46699), .Y(n46701) );
  NAND2X1 U48804 ( .A(n46702), .B(n46701), .Y(n46718) );
  NAND2X1 U48805 ( .A(n2576), .B(n43060), .Y(n46704) );
  NAND2X1 U48806 ( .A(n2574), .B(n39136), .Y(n46703) );
  NAND2X1 U48807 ( .A(n46704), .B(n46703), .Y(n46708) );
  NAND2X1 U48808 ( .A(n2566), .B(n43063), .Y(n46706) );
  NAND2X1 U48809 ( .A(n2557), .B(n43067), .Y(n46705) );
  NAND2X1 U48810 ( .A(n46706), .B(n46705), .Y(n46707) );
  NOR2X1 U48811 ( .A(n46708), .B(n46707), .Y(n46716) );
  NAND2X1 U48812 ( .A(n2562), .B(n43372), .Y(n46710) );
  NAND2X1 U48813 ( .A(n2568), .B(n43349), .Y(n46709) );
  NAND2X1 U48814 ( .A(n46710), .B(n46709), .Y(n46714) );
  NAND2X1 U48815 ( .A(n2560), .B(n43070), .Y(n46712) );
  NAND2X1 U48816 ( .A(n2553), .B(n43071), .Y(n46711) );
  NAND2X1 U48817 ( .A(n46712), .B(n46711), .Y(n46713) );
  NOR2X1 U48818 ( .A(n46714), .B(n46713), .Y(n46715) );
  NAND2X1 U48819 ( .A(n46716), .B(n46715), .Y(n46717) );
  NOR2X1 U48820 ( .A(n46718), .B(n46717), .Y(n46719) );
  NAND2X1 U48821 ( .A(n46720), .B(n46719), .Y(n46721) );
  NAND2X1 U48822 ( .A(n42804), .B(n46721), .Y(n46722) );
  NAND2X1 U48823 ( .A(n46723), .B(n46722), .Y(n73254) );
  NOR2X1 U48824 ( .A(n40862), .B(n37136), .Y(n46724) );
  NOR2X1 U48825 ( .A(n46725), .B(n46724), .Y(n46731) );
  NAND2X1 U48826 ( .A(n36733), .B(n40447), .Y(n49710) );
  NOR2X1 U48827 ( .A(n37130), .B(n42909), .Y(n46729) );
  NAND2X1 U48828 ( .A(n38604), .B(n46906), .Y(n46727) );
  NOR2X1 U48829 ( .A(n37133), .B(n46727), .Y(n46728) );
  NOR2X1 U48830 ( .A(n46729), .B(n46728), .Y(n46730) );
  NAND2X1 U48831 ( .A(n46731), .B(n46730), .Y(n59127) );
  NOR2X1 U48832 ( .A(n42901), .B(n37137), .Y(n46735) );
  OR2X1 U48833 ( .A(n42898), .B(n43178), .Y(n46733) );
  NAND2X1 U48834 ( .A(writeback_exec_value_w[21]), .B(n37976), .Y(n46732) );
  NAND2X1 U48835 ( .A(n46733), .B(n46732), .Y(n46734) );
  NOR2X1 U48836 ( .A(n46735), .B(n46734), .Y(n46740) );
  NOR2X1 U48837 ( .A(n42900), .B(n37139), .Y(n46738) );
  NAND2X1 U48838 ( .A(n40499), .B(n46736), .Y(n49637) );
  NOR2X1 U48839 ( .A(n49637), .B(n37142), .Y(n46737) );
  NOR2X1 U48840 ( .A(n46738), .B(n46737), .Y(n46739) );
  NAND2X1 U48841 ( .A(n46740), .B(n46739), .Y(n59126) );
  NAND2X1 U48842 ( .A(n2557), .B(n49705), .Y(n46745) );
  NAND2X1 U48843 ( .A(n46741), .B(n45610), .Y(n46742) );
  NOR2X1 U48844 ( .A(n37095), .B(n46742), .Y(n46743) );
  NAND2X1 U48845 ( .A(n46743), .B(n40152), .Y(n46744) );
  NAND2X1 U48846 ( .A(n46745), .B(n46744), .Y(n46749) );
  NAND2X1 U48847 ( .A(n2553), .B(n40432), .Y(n46747) );
  NAND2X1 U48848 ( .A(n2560), .B(n40531), .Y(n46746) );
  NAND2X1 U48849 ( .A(n46747), .B(n46746), .Y(n46748) );
  NOR2X1 U48850 ( .A(n49599), .B(n36990), .Y(n46753) );
  NAND2X1 U48851 ( .A(n2554), .B(n38844), .Y(n46751) );
  NAND2X1 U48852 ( .A(n46178), .B(n2575), .Y(n46750) );
  NAND2X1 U48853 ( .A(n46751), .B(n46750), .Y(n46752) );
  NOR2X1 U48854 ( .A(n46753), .B(n46752), .Y(n46757) );
  NOR2X1 U48855 ( .A(n49604), .B(n36981), .Y(n46755) );
  NOR2X1 U48856 ( .A(n42616), .B(n36999), .Y(n46754) );
  NOR2X1 U48857 ( .A(n46755), .B(n46754), .Y(n46756) );
  NOR2X1 U48858 ( .A(n42741), .B(n36979), .Y(n46761) );
  NAND2X1 U48859 ( .A(n2558), .B(n36610), .Y(n46758) );
  NAND2X1 U48860 ( .A(n46759), .B(n46758), .Y(n46760) );
  NOR2X1 U48861 ( .A(n46761), .B(n46760), .Y(n46765) );
  NOR2X1 U48862 ( .A(n38712), .B(n36962), .Y(n46763) );
  NOR2X1 U48863 ( .A(n46763), .B(n46762), .Y(n46764) );
  NOR2X1 U48864 ( .A(n42683), .B(n36948), .Y(n46769) );
  NAND2X1 U48865 ( .A(n49577), .B(n2578), .Y(n46767) );
  NAND2X1 U48866 ( .A(n46767), .B(n46766), .Y(n46768) );
  NOR2X1 U48867 ( .A(n45244), .B(n36953), .Y(n46771) );
  NOR2X1 U48868 ( .A(n45245), .B(n36971), .Y(n46770) );
  NOR2X1 U48869 ( .A(n49587), .B(n36959), .Y(n46776) );
  NAND2X1 U48870 ( .A(n2577), .B(n42223), .Y(n46774) );
  NOR2X1 U48871 ( .A(n40509), .B(n42695), .Y(n46772) );
  NAND2X1 U48872 ( .A(n46772), .B(n2579), .Y(n46773) );
  NAND2X1 U48873 ( .A(n46774), .B(n46773), .Y(n46775) );
  NOR2X1 U48874 ( .A(n46776), .B(n46775), .Y(n46780) );
  NOR2X1 U48875 ( .A(n42628), .B(n36973), .Y(n46778) );
  NOR2X1 U48876 ( .A(n39654), .B(n36986), .Y(n46777) );
  NOR2X1 U48877 ( .A(n46778), .B(n46777), .Y(n46779) );
  NAND2X1 U48878 ( .A(n46780), .B(n46779), .Y(n46781) );
  NOR2X1 U48879 ( .A(n46782), .B(n46781), .Y(n46783) );
  NAND2X1 U48880 ( .A(n46784), .B(n46783), .Y(n46785) );
  NAND2X1 U48881 ( .A(n43939), .B(n42712), .Y(n57873) );
  NAND2X1 U48882 ( .A(n46786), .B(n57873), .Y(n57883) );
  INVX1 U48883 ( .A(n57883), .Y(n73436) );
  INVX1 U48884 ( .A(mem_d_data_rd_i[20]), .Y(n73549) );
  NAND2X1 U48885 ( .A(n40935), .B(n73549), .Y(n46787) );
  NOR2X1 U48886 ( .A(n43454), .B(n43171), .Y(n46789) );
  NOR2X1 U48887 ( .A(n43022), .B(n43174), .Y(n46788) );
  NAND2X1 U48888 ( .A(n2414), .B(n43362), .Y(n46791) );
  NAND2X1 U48889 ( .A(n2389), .B(n38413), .Y(n46790) );
  NAND2X1 U48890 ( .A(n46791), .B(n46790), .Y(n46795) );
  NAND2X1 U48891 ( .A(n2396), .B(n38402), .Y(n46793) );
  NAND2X1 U48892 ( .A(n2404), .B(n43027), .Y(n46792) );
  NAND2X1 U48893 ( .A(n46793), .B(n46792), .Y(n46794) );
  NOR2X1 U48894 ( .A(n46795), .B(n46794), .Y(n46803) );
  NAND2X1 U48895 ( .A(n2386), .B(n43030), .Y(n46797) );
  NAND2X1 U48896 ( .A(n2391), .B(n43032), .Y(n46796) );
  NAND2X1 U48897 ( .A(n46797), .B(n46796), .Y(n46801) );
  NAND2X1 U48898 ( .A(n2406), .B(n43036), .Y(n46799) );
  NAND2X1 U48899 ( .A(n2398), .B(n43351), .Y(n46798) );
  NAND2X1 U48900 ( .A(n46799), .B(n46798), .Y(n46800) );
  NOR2X1 U48901 ( .A(n46801), .B(n46800), .Y(n46802) );
  NAND2X1 U48902 ( .A(n46803), .B(n46802), .Y(n46819) );
  NAND2X1 U48903 ( .A(n2402), .B(n43355), .Y(n46805) );
  NAND2X1 U48904 ( .A(n2400), .B(n43039), .Y(n46804) );
  NAND2X1 U48905 ( .A(n46805), .B(n46804), .Y(n46809) );
  NAND2X1 U48906 ( .A(n1829), .B(n39806), .Y(n46807) );
  NAND2X1 U48907 ( .A(n2408), .B(n43042), .Y(n46806) );
  NAND2X1 U48908 ( .A(n46807), .B(n46806), .Y(n46808) );
  NOR2X1 U48909 ( .A(n46809), .B(n46808), .Y(n46817) );
  NAND2X1 U48910 ( .A(n2412), .B(n38390), .Y(n46811) );
  NAND2X1 U48911 ( .A(n2387), .B(n43345), .Y(n46810) );
  NAND2X1 U48912 ( .A(n46811), .B(n46810), .Y(n46815) );
  NAND2X1 U48913 ( .A(n2394), .B(n43338), .Y(n46813) );
  NAND2X1 U48914 ( .A(n2410), .B(n43365), .Y(n46812) );
  NAND2X1 U48915 ( .A(n46813), .B(n46812), .Y(n46814) );
  NOR2X1 U48916 ( .A(n46815), .B(n46814), .Y(n46816) );
  NAND2X1 U48917 ( .A(n46817), .B(n46816), .Y(n46818) );
  NOR2X1 U48918 ( .A(n46819), .B(n46818), .Y(n46849) );
  NAND2X1 U48919 ( .A(n2407), .B(n43044), .Y(n46821) );
  NAND2X1 U48920 ( .A(n2413), .B(n43047), .Y(n46820) );
  NAND2X1 U48921 ( .A(n46821), .B(n46820), .Y(n46825) );
  NAND2X1 U48922 ( .A(n2405), .B(n43049), .Y(n46823) );
  NAND2X1 U48923 ( .A(n2390), .B(n43051), .Y(n46822) );
  NAND2X1 U48924 ( .A(n46823), .B(n46822), .Y(n46824) );
  NOR2X1 U48925 ( .A(n46825), .B(n46824), .Y(n46831) );
  NOR2X1 U48926 ( .A(n43370), .B(n37316), .Y(n46829) );
  NAND2X1 U48927 ( .A(n2393), .B(n43054), .Y(n46827) );
  NAND2X1 U48928 ( .A(n2415), .B(n43057), .Y(n46826) );
  NAND2X1 U48929 ( .A(n46827), .B(n46826), .Y(n46828) );
  NOR2X1 U48930 ( .A(n46829), .B(n46828), .Y(n46830) );
  NAND2X1 U48931 ( .A(n46831), .B(n46830), .Y(n46847) );
  NAND2X1 U48932 ( .A(n2411), .B(n43060), .Y(n46833) );
  NAND2X1 U48933 ( .A(n2409), .B(n39139), .Y(n46832) );
  NAND2X1 U48934 ( .A(n46833), .B(n46832), .Y(n46837) );
  NAND2X1 U48935 ( .A(n2401), .B(n43063), .Y(n46835) );
  NAND2X1 U48936 ( .A(n2392), .B(n43067), .Y(n46834) );
  NAND2X1 U48937 ( .A(n46835), .B(n46834), .Y(n46836) );
  NOR2X1 U48938 ( .A(n46837), .B(n46836), .Y(n46845) );
  NAND2X1 U48939 ( .A(n2397), .B(n43372), .Y(n46839) );
  NAND2X1 U48940 ( .A(n2403), .B(n43350), .Y(n46838) );
  NAND2X1 U48941 ( .A(n46839), .B(n46838), .Y(n46843) );
  NAND2X1 U48942 ( .A(n2395), .B(n43070), .Y(n46841) );
  NAND2X1 U48943 ( .A(n2388), .B(n43071), .Y(n46840) );
  NAND2X1 U48944 ( .A(n46841), .B(n46840), .Y(n46842) );
  NOR2X1 U48945 ( .A(n46843), .B(n46842), .Y(n46844) );
  NAND2X1 U48946 ( .A(n46845), .B(n46844), .Y(n46846) );
  NOR2X1 U48947 ( .A(n46847), .B(n46846), .Y(n46848) );
  NAND2X1 U48948 ( .A(n46849), .B(n46848), .Y(n46850) );
  NAND2X1 U48949 ( .A(n43931), .B(n43939), .Y(n57869) );
  INVX1 U48950 ( .A(n57869), .Y(n58928) );
  NOR2X1 U48951 ( .A(n42910), .B(n37180), .Y(n46854) );
  NAND2X1 U48952 ( .A(n2392), .B(n49705), .Y(n46852) );
  NAND2X1 U48953 ( .A(n2408), .B(n42830), .Y(n46851) );
  NAND2X1 U48954 ( .A(n46852), .B(n46851), .Y(n46853) );
  NOR2X1 U48955 ( .A(n42893), .B(n37041), .Y(n46858) );
  NAND2X1 U48956 ( .A(n2398), .B(n40514), .Y(n46856) );
  NAND2X1 U48957 ( .A(n42882), .B(n40513), .Y(n49400) );
  NAND2X1 U48958 ( .A(n2410), .B(n38085), .Y(n46855) );
  NAND2X1 U48959 ( .A(n46856), .B(n46855), .Y(n46857) );
  NOR2X1 U48960 ( .A(n46858), .B(n46857), .Y(n46862) );
  NOR2X1 U48961 ( .A(n38752), .B(n37050), .Y(n46860) );
  NOR2X1 U48962 ( .A(n42616), .B(n37062), .Y(n46859) );
  NOR2X1 U48963 ( .A(n46860), .B(n46859), .Y(n46861) );
  NAND2X1 U48964 ( .A(n46862), .B(n46861), .Y(n46872) );
  NOR2X1 U48965 ( .A(n42741), .B(n37052), .Y(n46866) );
  NAND2X1 U48966 ( .A(n2399), .B(n42821), .Y(n46864) );
  NAND2X1 U48967 ( .A(n2393), .B(n36610), .Y(n46863) );
  NAND2X1 U48968 ( .A(n46864), .B(n46863), .Y(n46865) );
  NOR2X1 U48969 ( .A(n46866), .B(n46865), .Y(n46870) );
  NOR2X1 U48970 ( .A(n38712), .B(n37061), .Y(n46868) );
  NOR2X1 U48971 ( .A(n42776), .B(n37070), .Y(n46867) );
  NOR2X1 U48972 ( .A(n46868), .B(n46867), .Y(n46869) );
  NAND2X1 U48973 ( .A(n46870), .B(n46869), .Y(n46871) );
  NOR2X1 U48974 ( .A(n46872), .B(n46871), .Y(n46892) );
  NOR2X1 U48975 ( .A(n42683), .B(n37051), .Y(n46876) );
  NAND2X1 U48976 ( .A(n2413), .B(n47895), .Y(n46874) );
  NAND2X1 U48977 ( .A(n2391), .B(n40248), .Y(n46873) );
  NAND2X1 U48978 ( .A(n46874), .B(n46873), .Y(n46875) );
  NOR2X1 U48979 ( .A(n46876), .B(n46875), .Y(n46880) );
  NOR2X1 U48980 ( .A(n45244), .B(n37055), .Y(n46878) );
  NOR2X1 U48981 ( .A(n40427), .B(n37068), .Y(n46877) );
  NOR2X1 U48982 ( .A(n46878), .B(n46877), .Y(n46879) );
  NAND2X1 U48983 ( .A(n46880), .B(n46879), .Y(n46890) );
  NOR2X1 U48984 ( .A(n42905), .B(n37060), .Y(n46884) );
  NAND2X1 U48985 ( .A(n2415), .B(n42619), .Y(n46882) );
  NAND2X1 U48986 ( .A(n2414), .B(n42147), .Y(n46881) );
  NAND2X1 U48987 ( .A(n46882), .B(n46881), .Y(n46883) );
  NOR2X1 U48988 ( .A(n46884), .B(n46883), .Y(n46888) );
  NOR2X1 U48989 ( .A(n42628), .B(n37069), .Y(n46886) );
  NOR2X1 U48990 ( .A(n39654), .B(n37073), .Y(n46885) );
  NOR2X1 U48991 ( .A(n46886), .B(n46885), .Y(n46887) );
  NAND2X1 U48992 ( .A(n46888), .B(n46887), .Y(n46889) );
  NOR2X1 U48993 ( .A(n46890), .B(n46889), .Y(n46891) );
  NAND2X1 U48994 ( .A(n46892), .B(n46891), .Y(n46893) );
  INVX1 U48995 ( .A(n49625), .Y(n49648) );
  NAND2X1 U48996 ( .A(n2411), .B(n49648), .Y(n46896) );
  NAND2X1 U48997 ( .A(n2400), .B(n49719), .Y(n46895) );
  NAND2X1 U48998 ( .A(n46896), .B(n46895), .Y(n46902) );
  NOR2X1 U48999 ( .A(n49715), .B(n43175), .Y(n46898) );
  NOR2X1 U49000 ( .A(n42898), .B(n43173), .Y(n46897) );
  NOR2X1 U49001 ( .A(n46898), .B(n46897), .Y(n46900) );
  NAND2X1 U49002 ( .A(n2409), .B(n40521), .Y(n46899) );
  NAND2X1 U49003 ( .A(n46900), .B(n46899), .Y(n46901) );
  NOR2X1 U49004 ( .A(n46902), .B(n46901), .Y(n46914) );
  NOR2X1 U49005 ( .A(n37114), .B(n40517), .Y(n46905) );
  NOR2X1 U49006 ( .A(n46903), .B(n37118), .Y(n46904) );
  NOR2X1 U49007 ( .A(n46905), .B(n46904), .Y(n46908) );
  INVX1 U49008 ( .A(n46727), .Y(n49709) );
  NAND2X1 U49009 ( .A(n1829), .B(n49709), .Y(n46907) );
  NAND2X1 U49010 ( .A(n46908), .B(n46907), .Y(n46912) );
  NAND2X1 U49011 ( .A(n2401), .B(n41741), .Y(n46910) );
  INVX1 U49012 ( .A(n42911), .Y(n49706) );
  NAND2X1 U49013 ( .A(n2386), .B(n49706), .Y(n46909) );
  NAND2X1 U49014 ( .A(n46910), .B(n46909), .Y(n46911) );
  NOR2X1 U49015 ( .A(n46912), .B(n46911), .Y(n46913) );
  NAND2X1 U49016 ( .A(n46914), .B(n46913), .Y(n46915) );
  NAND2X1 U49017 ( .A(n43938), .B(n42659), .Y(n46917) );
  NAND2X1 U49018 ( .A(n43931), .B(n42712), .Y(n46916) );
  NAND2X1 U49019 ( .A(n46917), .B(n46916), .Y(n57872) );
  NOR2X1 U49020 ( .A(n58928), .B(n57872), .Y(n46918) );
  NAND2X1 U49021 ( .A(n42661), .B(n42711), .Y(n57870) );
  NAND2X1 U49022 ( .A(n46918), .B(n57870), .Y(n49797) );
  NOR2X1 U49023 ( .A(n42908), .B(n37150), .Y(n46920) );
  NOR2X1 U49024 ( .A(n38798), .B(n37156), .Y(n46919) );
  NOR2X1 U49025 ( .A(n46920), .B(n46919), .Y(n46922) );
  INVX1 U49026 ( .A(n49573), .Y(n49647) );
  NAND2X1 U49027 ( .A(n2887), .B(n42707), .Y(n46921) );
  NAND2X1 U49028 ( .A(n46922), .B(n46921), .Y(n46973) );
  NOR2X1 U49029 ( .A(n40847), .B(n37152), .Y(n46926) );
  NAND2X1 U49030 ( .A(n2908), .B(n40521), .Y(n46924) );
  NAND2X1 U49031 ( .A(n2907), .B(n42830), .Y(n46923) );
  NAND2X1 U49032 ( .A(n46924), .B(n46923), .Y(n46925) );
  NOR2X1 U49033 ( .A(n46926), .B(n46925), .Y(n46971) );
  NOR2X1 U49034 ( .A(n42683), .B(n36954), .Y(n46933) );
  NOR2X1 U49035 ( .A(n40510), .B(n46927), .Y(n46928) );
  NAND2X1 U49036 ( .A(n46928), .B(n2912), .Y(n46931) );
  NOR2X1 U49037 ( .A(n39809), .B(n42693), .Y(n46929) );
  NAND2X1 U49038 ( .A(n46929), .B(n2891), .Y(n46930) );
  NAND2X1 U49039 ( .A(n46931), .B(n46930), .Y(n46932) );
  NOR2X1 U49040 ( .A(n46933), .B(n46932), .Y(n46937) );
  NOR2X1 U49041 ( .A(n45244), .B(n36964), .Y(n46935) );
  NOR2X1 U49042 ( .A(n40427), .B(n36991), .Y(n46934) );
  NOR2X1 U49043 ( .A(n46935), .B(n46934), .Y(n46936) );
  NAND2X1 U49044 ( .A(n46937), .B(n46936), .Y(n46947) );
  NOR2X1 U49045 ( .A(n49587), .B(n36972), .Y(n46941) );
  NAND2X1 U49046 ( .A(n46167), .B(n2911), .Y(n46939) );
  NAND2X1 U49047 ( .A(n46772), .B(n2913), .Y(n46938) );
  NAND2X1 U49048 ( .A(n46939), .B(n46938), .Y(n46940) );
  NOR2X1 U49049 ( .A(n46941), .B(n46940), .Y(n46945) );
  NOR2X1 U49050 ( .A(n42629), .B(n36993), .Y(n46943) );
  NOR2X1 U49051 ( .A(n39654), .B(n37006), .Y(n46942) );
  NOR2X1 U49052 ( .A(n46943), .B(n46942), .Y(n46944) );
  NAND2X1 U49053 ( .A(n46945), .B(n46944), .Y(n46946) );
  NOR2X1 U49054 ( .A(n46947), .B(n46946), .Y(n46968) );
  NOR2X1 U49055 ( .A(n49599), .B(n36960), .Y(n46952) );
  NAND2X1 U49056 ( .A(n2888), .B(n57621), .Y(n46950) );
  NOR2X1 U49057 ( .A(n40511), .B(n36608), .Y(n46948) );
  NAND2X1 U49058 ( .A(n46948), .B(n2909), .Y(n46949) );
  NAND2X1 U49059 ( .A(n46950), .B(n46949), .Y(n46951) );
  NOR2X1 U49060 ( .A(n46952), .B(n46951), .Y(n46956) );
  NOR2X1 U49061 ( .A(n38752), .B(n36987), .Y(n46954) );
  NOR2X1 U49062 ( .A(n38701), .B(n37007), .Y(n46953) );
  NOR2X1 U49063 ( .A(n46954), .B(n46953), .Y(n46955) );
  NAND2X1 U49064 ( .A(n46956), .B(n46955), .Y(n46966) );
  NOR2X1 U49065 ( .A(n42741), .B(n36988), .Y(n46960) );
  NAND2X1 U49066 ( .A(n2898), .B(n42821), .Y(n46958) );
  NAND2X1 U49067 ( .A(n2892), .B(n49611), .Y(n46957) );
  NAND2X1 U49068 ( .A(n46958), .B(n46957), .Y(n46959) );
  NOR2X1 U49069 ( .A(n46960), .B(n46959), .Y(n46964) );
  NOR2X1 U49070 ( .A(n38711), .B(n37004), .Y(n46962) );
  NOR2X1 U49071 ( .A(n42775), .B(n37015), .Y(n46961) );
  NOR2X1 U49072 ( .A(n46962), .B(n46961), .Y(n46963) );
  NAND2X1 U49073 ( .A(n46964), .B(n46963), .Y(n46965) );
  NOR2X1 U49074 ( .A(n46966), .B(n46965), .Y(n46967) );
  NAND2X1 U49075 ( .A(n46968), .B(n46967), .Y(n46969) );
  NAND2X1 U49076 ( .A(n40490), .B(n46969), .Y(n46970) );
  NAND2X1 U49077 ( .A(n46971), .B(n46970), .Y(n46972) );
  INVX1 U49078 ( .A(mem_d_data_rd_i[17]), .Y(n73552) );
  NAND2X1 U49079 ( .A(n40935), .B(n73552), .Y(n46974) );
  NAND2X1 U49080 ( .A(writeback_exec_value_w[17]), .B(n43020), .Y(n46975) );
  NAND2X1 U49081 ( .A(n46976), .B(n46975), .Y(n46985) );
  NOR2X1 U49082 ( .A(n42909), .B(n37159), .Y(n46978) );
  NOR2X1 U49083 ( .A(n46727), .B(n37166), .Y(n46977) );
  NOR2X1 U49084 ( .A(n46978), .B(n46977), .Y(n46983) );
  NOR2X1 U49085 ( .A(n40855), .B(n37165), .Y(n46981) );
  NOR2X1 U49086 ( .A(n42917), .B(n37169), .Y(n46980) );
  NOR2X1 U49087 ( .A(n46981), .B(n46980), .Y(n46982) );
  NAND2X1 U49088 ( .A(n46983), .B(n46982), .Y(n46984) );
  NOR2X1 U49089 ( .A(n43454), .B(n43156), .Y(n46987) );
  NOR2X1 U49090 ( .A(n43022), .B(n43157), .Y(n46986) );
  NOR2X1 U49091 ( .A(n46987), .B(n46986), .Y(n47050) );
  NAND2X1 U49092 ( .A(n2913), .B(n43362), .Y(n46989) );
  NAND2X1 U49093 ( .A(n2888), .B(n38407), .Y(n46988) );
  NAND2X1 U49094 ( .A(n46989), .B(n46988), .Y(n46993) );
  NAND2X1 U49095 ( .A(n2895), .B(n43344), .Y(n46991) );
  NAND2X1 U49096 ( .A(n2903), .B(n43027), .Y(n46990) );
  NAND2X1 U49097 ( .A(n46991), .B(n46990), .Y(n46992) );
  NOR2X1 U49098 ( .A(n46993), .B(n46992), .Y(n47001) );
  NAND2X1 U49099 ( .A(n2885), .B(n43030), .Y(n46995) );
  NAND2X1 U49100 ( .A(n2891), .B(n43033), .Y(n46994) );
  NAND2X1 U49101 ( .A(n46995), .B(n46994), .Y(n46999) );
  NAND2X1 U49102 ( .A(n2905), .B(n43036), .Y(n46997) );
  NAND2X1 U49103 ( .A(n2897), .B(n43352), .Y(n46996) );
  NAND2X1 U49104 ( .A(n46997), .B(n46996), .Y(n46998) );
  NOR2X1 U49105 ( .A(n46999), .B(n46998), .Y(n47000) );
  NAND2X1 U49106 ( .A(n47001), .B(n47000), .Y(n47017) );
  NAND2X1 U49107 ( .A(n2901), .B(n43354), .Y(n47003) );
  NAND2X1 U49108 ( .A(n2899), .B(n43039), .Y(n47002) );
  NAND2X1 U49109 ( .A(n47003), .B(n47002), .Y(n47007) );
  NAND2X1 U49110 ( .A(n1808), .B(n39803), .Y(n47005) );
  NAND2X1 U49111 ( .A(n2907), .B(n43042), .Y(n47004) );
  NAND2X1 U49112 ( .A(n47005), .B(n47004), .Y(n47006) );
  NOR2X1 U49113 ( .A(n47007), .B(n47006), .Y(n47015) );
  NAND2X1 U49114 ( .A(n2911), .B(n43360), .Y(n47009) );
  NAND2X1 U49115 ( .A(n2886), .B(n43346), .Y(n47008) );
  NAND2X1 U49116 ( .A(n47009), .B(n47008), .Y(n47013) );
  NAND2X1 U49117 ( .A(n2893), .B(n43339), .Y(n47011) );
  NAND2X1 U49118 ( .A(n2909), .B(n43366), .Y(n47010) );
  NAND2X1 U49119 ( .A(n47011), .B(n47010), .Y(n47012) );
  NOR2X1 U49120 ( .A(n47013), .B(n47012), .Y(n47014) );
  NAND2X1 U49121 ( .A(n47015), .B(n47014), .Y(n47016) );
  NOR2X1 U49122 ( .A(n47017), .B(n47016), .Y(n47047) );
  NAND2X1 U49123 ( .A(n2906), .B(n43044), .Y(n47019) );
  NAND2X1 U49124 ( .A(n2912), .B(n43047), .Y(n47018) );
  NAND2X1 U49125 ( .A(n47019), .B(n47018), .Y(n47023) );
  NAND2X1 U49126 ( .A(n2904), .B(n43049), .Y(n47021) );
  NAND2X1 U49127 ( .A(n2889), .B(n43052), .Y(n47020) );
  NAND2X1 U49128 ( .A(n47021), .B(n47020), .Y(n47022) );
  NOR2X1 U49129 ( .A(n47023), .B(n47022), .Y(n47029) );
  NOR2X1 U49130 ( .A(n43371), .B(n37314), .Y(n47027) );
  NAND2X1 U49131 ( .A(n2892), .B(n43054), .Y(n47025) );
  NAND2X1 U49132 ( .A(n2914), .B(n43057), .Y(n47024) );
  NAND2X1 U49133 ( .A(n47025), .B(n47024), .Y(n47026) );
  NOR2X1 U49134 ( .A(n47027), .B(n47026), .Y(n47028) );
  NAND2X1 U49135 ( .A(n47029), .B(n47028), .Y(n47045) );
  NAND2X1 U49136 ( .A(n2910), .B(n43061), .Y(n47031) );
  NAND2X1 U49137 ( .A(n2908), .B(n39133), .Y(n47030) );
  NAND2X1 U49138 ( .A(n47031), .B(n47030), .Y(n47035) );
  NAND2X1 U49139 ( .A(n2900), .B(n43063), .Y(n47033) );
  NAND2X1 U49140 ( .A(n2890), .B(n43067), .Y(n47032) );
  NAND2X1 U49141 ( .A(n47033), .B(n47032), .Y(n47034) );
  NOR2X1 U49142 ( .A(n47035), .B(n47034), .Y(n47043) );
  NAND2X1 U49143 ( .A(n2896), .B(n38528), .Y(n47037) );
  NAND2X1 U49144 ( .A(n2902), .B(n43350), .Y(n47036) );
  NAND2X1 U49145 ( .A(n47037), .B(n47036), .Y(n47041) );
  NAND2X1 U49146 ( .A(n2894), .B(n43069), .Y(n47039) );
  NAND2X1 U49147 ( .A(n2887), .B(n43072), .Y(n47038) );
  NAND2X1 U49148 ( .A(n47039), .B(n47038), .Y(n47040) );
  NOR2X1 U49149 ( .A(n47041), .B(n47040), .Y(n47042) );
  NAND2X1 U49150 ( .A(n47043), .B(n47042), .Y(n47044) );
  NOR2X1 U49151 ( .A(n47045), .B(n47044), .Y(n47046) );
  NAND2X1 U49152 ( .A(n47047), .B(n47046), .Y(n47048) );
  NAND2X1 U49153 ( .A(n42806), .B(n47048), .Y(n47049) );
  NAND2X1 U49154 ( .A(n47050), .B(n47049), .Y(n73224) );
  NAND2X1 U49155 ( .A(n42642), .B(n43904), .Y(n57662) );
  INVX1 U49156 ( .A(n57662), .Y(n57833) );
  INVX1 U49157 ( .A(mem_d_data_rd_i[16]), .Y(n73553) );
  NAND2X1 U49158 ( .A(n40935), .B(n73553), .Y(n47051) );
  NOR2X1 U49159 ( .A(n43454), .B(n43148), .Y(n47053) );
  NOR2X1 U49160 ( .A(n43022), .B(n43151), .Y(n47052) );
  NOR2X1 U49161 ( .A(n47053), .B(n47052), .Y(n47116) );
  NAND2X1 U49162 ( .A(n2547), .B(n43362), .Y(n47055) );
  NAND2X1 U49163 ( .A(n2522), .B(n38413), .Y(n47054) );
  NAND2X1 U49164 ( .A(n47055), .B(n47054), .Y(n47059) );
  NAND2X1 U49165 ( .A(n2529), .B(n38402), .Y(n47057) );
  NAND2X1 U49166 ( .A(n2537), .B(n38602), .Y(n47056) );
  NAND2X1 U49167 ( .A(n47057), .B(n47056), .Y(n47058) );
  NOR2X1 U49168 ( .A(n47059), .B(n47058), .Y(n47067) );
  NAND2X1 U49169 ( .A(n2519), .B(n43030), .Y(n47061) );
  NAND2X1 U49170 ( .A(n2525), .B(n43033), .Y(n47060) );
  NAND2X1 U49171 ( .A(n47061), .B(n47060), .Y(n47065) );
  NAND2X1 U49172 ( .A(n2539), .B(n38534), .Y(n47063) );
  NAND2X1 U49173 ( .A(n2531), .B(n43352), .Y(n47062) );
  NAND2X1 U49174 ( .A(n47063), .B(n47062), .Y(n47064) );
  NOR2X1 U49175 ( .A(n47065), .B(n47064), .Y(n47066) );
  NAND2X1 U49176 ( .A(n47067), .B(n47066), .Y(n47083) );
  NAND2X1 U49177 ( .A(n2535), .B(n43354), .Y(n47069) );
  NAND2X1 U49178 ( .A(n2533), .B(n43039), .Y(n47068) );
  NAND2X1 U49179 ( .A(n47069), .B(n47068), .Y(n47073) );
  NAND2X1 U49180 ( .A(n1823), .B(n39802), .Y(n47071) );
  NAND2X1 U49181 ( .A(n2541), .B(n43043), .Y(n47070) );
  NAND2X1 U49182 ( .A(n47071), .B(n47070), .Y(n47072) );
  NOR2X1 U49183 ( .A(n47073), .B(n47072), .Y(n47081) );
  NAND2X1 U49184 ( .A(n2545), .B(n38390), .Y(n47075) );
  NAND2X1 U49185 ( .A(n2520), .B(n43346), .Y(n47074) );
  NAND2X1 U49186 ( .A(n47075), .B(n47074), .Y(n47079) );
  NAND2X1 U49187 ( .A(n2527), .B(n43339), .Y(n47077) );
  NAND2X1 U49188 ( .A(n2543), .B(n43366), .Y(n47076) );
  NAND2X1 U49189 ( .A(n47077), .B(n47076), .Y(n47078) );
  NOR2X1 U49190 ( .A(n47079), .B(n47078), .Y(n47080) );
  NAND2X1 U49191 ( .A(n47081), .B(n47080), .Y(n47082) );
  NOR2X1 U49192 ( .A(n47083), .B(n47082), .Y(n47113) );
  NAND2X1 U49193 ( .A(n2540), .B(n40273), .Y(n47085) );
  NAND2X1 U49194 ( .A(n2546), .B(n43048), .Y(n47084) );
  NAND2X1 U49195 ( .A(n47085), .B(n47084), .Y(n47089) );
  NAND2X1 U49196 ( .A(n2538), .B(n43050), .Y(n47087) );
  NAND2X1 U49197 ( .A(n2523), .B(n43052), .Y(n47086) );
  NAND2X1 U49198 ( .A(n47087), .B(n47086), .Y(n47088) );
  NOR2X1 U49199 ( .A(n47089), .B(n47088), .Y(n47095) );
  NOR2X1 U49200 ( .A(n43370), .B(n36875), .Y(n47093) );
  NAND2X1 U49201 ( .A(n2526), .B(n38577), .Y(n47091) );
  NAND2X1 U49202 ( .A(n2548), .B(n43057), .Y(n47090) );
  NAND2X1 U49203 ( .A(n47091), .B(n47090), .Y(n47092) );
  NOR2X1 U49204 ( .A(n47093), .B(n47092), .Y(n47094) );
  NAND2X1 U49205 ( .A(n47095), .B(n47094), .Y(n47111) );
  NAND2X1 U49206 ( .A(n2544), .B(n43061), .Y(n47097) );
  NAND2X1 U49207 ( .A(n2542), .B(n39132), .Y(n47096) );
  NAND2X1 U49208 ( .A(n47097), .B(n47096), .Y(n47101) );
  NAND2X1 U49209 ( .A(n2534), .B(n40158), .Y(n47099) );
  NAND2X1 U49210 ( .A(n2524), .B(n43067), .Y(n47098) );
  NAND2X1 U49211 ( .A(n47099), .B(n47098), .Y(n47100) );
  NOR2X1 U49212 ( .A(n47101), .B(n47100), .Y(n47109) );
  NAND2X1 U49213 ( .A(n2530), .B(n38528), .Y(n47103) );
  NAND2X1 U49214 ( .A(n2536), .B(n43349), .Y(n47102) );
  NAND2X1 U49215 ( .A(n47103), .B(n47102), .Y(n47107) );
  NAND2X1 U49216 ( .A(n2528), .B(n43069), .Y(n47105) );
  NAND2X1 U49217 ( .A(n2521), .B(n43072), .Y(n47104) );
  NAND2X1 U49218 ( .A(n47105), .B(n47104), .Y(n47106) );
  NOR2X1 U49219 ( .A(n47107), .B(n47106), .Y(n47108) );
  NAND2X1 U49220 ( .A(n47109), .B(n47108), .Y(n47110) );
  NOR2X1 U49221 ( .A(n47111), .B(n47110), .Y(n47112) );
  NAND2X1 U49222 ( .A(n47113), .B(n47112), .Y(n47114) );
  NAND2X1 U49223 ( .A(n42805), .B(n47114), .Y(n47115) );
  NAND2X1 U49224 ( .A(n47116), .B(n47115), .Y(n73216) );
  NOR2X1 U49225 ( .A(n49625), .B(n37119), .Y(n47118) );
  NOR2X1 U49226 ( .A(n38798), .B(n37120), .Y(n47117) );
  NOR2X1 U49227 ( .A(n47118), .B(n47117), .Y(n47120) );
  NAND2X1 U49228 ( .A(n2521), .B(n49647), .Y(n47119) );
  NAND2X1 U49229 ( .A(n47120), .B(n47119), .Y(n47165) );
  NOR2X1 U49230 ( .A(n42915), .B(n37192), .Y(n47161) );
  NAND2X1 U49231 ( .A(n2523), .B(n40520), .Y(n47122) );
  NAND2X1 U49232 ( .A(n2538), .B(n42626), .Y(n47121) );
  NAND2X1 U49233 ( .A(n47122), .B(n47121), .Y(n47128) );
  NOR2X1 U49234 ( .A(n42903), .B(n36865), .Y(n47124) );
  NOR2X1 U49235 ( .A(n49678), .B(n36872), .Y(n47123) );
  NOR2X1 U49236 ( .A(n47124), .B(n47123), .Y(n47126) );
  NAND2X1 U49237 ( .A(n2548), .B(n42618), .Y(n47125) );
  NAND2X1 U49238 ( .A(n47126), .B(n47125), .Y(n47127) );
  NOR2X1 U49239 ( .A(n47128), .B(n47127), .Y(n47138) );
  NAND2X1 U49240 ( .A(n2537), .B(n40424), .Y(n47130) );
  NAND2X1 U49241 ( .A(n2539), .B(n40535), .Y(n47129) );
  NAND2X1 U49242 ( .A(n47130), .B(n47129), .Y(n47136) );
  NOR2X1 U49243 ( .A(n45870), .B(n36867), .Y(n47132) );
  NOR2X1 U49244 ( .A(n42682), .B(n36876), .Y(n47131) );
  NOR2X1 U49245 ( .A(n47132), .B(n47131), .Y(n47134) );
  NAND2X1 U49246 ( .A(n2546), .B(n47895), .Y(n47133) );
  NAND2X1 U49247 ( .A(n47134), .B(n47133), .Y(n47135) );
  NOR2X1 U49248 ( .A(n47136), .B(n47135), .Y(n47137) );
  NAND2X1 U49249 ( .A(n47138), .B(n47137), .Y(n47158) );
  NAND2X1 U49250 ( .A(n2529), .B(n42779), .Y(n47140) );
  NAND2X1 U49251 ( .A(n2520), .B(n38709), .Y(n47139) );
  NAND2X1 U49252 ( .A(n47140), .B(n47139), .Y(n47146) );
  NOR2X1 U49253 ( .A(n42892), .B(n36871), .Y(n47142) );
  NOR2X1 U49254 ( .A(n42895), .B(n36875), .Y(n47141) );
  NOR2X1 U49255 ( .A(n47142), .B(n47141), .Y(n47144) );
  INVX1 U49256 ( .A(n49610), .Y(n73368) );
  NAND2X1 U49257 ( .A(n2527), .B(n42675), .Y(n47143) );
  NAND2X1 U49258 ( .A(n47144), .B(n47143), .Y(n47145) );
  NOR2X1 U49259 ( .A(n47146), .B(n47145), .Y(n47156) );
  INVX1 U49260 ( .A(n49605), .Y(n57615) );
  NAND2X1 U49261 ( .A(n2535), .B(n46177), .Y(n47148) );
  NAND2X1 U49262 ( .A(n2530), .B(n39319), .Y(n47147) );
  NAND2X1 U49263 ( .A(n47148), .B(n47147), .Y(n47154) );
  NOR2X1 U49264 ( .A(n49665), .B(n36879), .Y(n47150) );
  NOR2X1 U49265 ( .A(n42893), .B(n36874), .Y(n47149) );
  NOR2X1 U49266 ( .A(n47149), .B(n47150), .Y(n47152) );
  NAND2X1 U49267 ( .A(n2531), .B(n40515), .Y(n47151) );
  NAND2X1 U49268 ( .A(n47152), .B(n47151), .Y(n47153) );
  NOR2X1 U49269 ( .A(n47154), .B(n47153), .Y(n47155) );
  NAND2X1 U49270 ( .A(n47156), .B(n47155), .Y(n47157) );
  NOR2X1 U49271 ( .A(n47158), .B(n47157), .Y(n47159) );
  NOR2X1 U49272 ( .A(n47159), .B(n42887), .Y(n47160) );
  NOR2X1 U49273 ( .A(n47161), .B(n47160), .Y(n47164) );
  NOR2X1 U49274 ( .A(n40277), .B(n37154), .Y(n47163) );
  NOR2X1 U49275 ( .A(n42901), .B(n37160), .Y(n47162) );
  NOR2X1 U49276 ( .A(n42900), .B(n37164), .Y(n47167) );
  NOR2X1 U49277 ( .A(n43150), .B(n40360), .Y(n47166) );
  NOR2X1 U49278 ( .A(n47167), .B(n47166), .Y(n47169) );
  NAND2X1 U49279 ( .A(writeback_exec_value_w[16]), .B(n43020), .Y(n47168) );
  NAND2X1 U49280 ( .A(n47169), .B(n47168), .Y(n47177) );
  NOR2X1 U49281 ( .A(n42910), .B(n37168), .Y(n47171) );
  NOR2X1 U49282 ( .A(n46727), .B(n37171), .Y(n47170) );
  NOR2X1 U49283 ( .A(n47171), .B(n47170), .Y(n47175) );
  NOR2X1 U49284 ( .A(n49637), .B(n37170), .Y(n47173) );
  NOR2X1 U49285 ( .A(n42918), .B(n37172), .Y(n47172) );
  NOR2X1 U49286 ( .A(n47173), .B(n47172), .Y(n47174) );
  NAND2X1 U49287 ( .A(n47175), .B(n47174), .Y(n47176) );
  NAND2X1 U49288 ( .A(n43901), .B(n43724), .Y(n57838) );
  INVX1 U49289 ( .A(n57838), .Y(n57637) );
  INVX1 U49290 ( .A(n31921), .Y(n47178) );
  NOR2X1 U49291 ( .A(n47178), .B(n429), .Y(n47180) );
  NAND2X1 U49292 ( .A(n34489), .B(n34490), .Y(n47179) );
  NOR2X1 U49293 ( .A(n43092), .B(n43455), .Y(n47182) );
  NOR2X1 U49294 ( .A(n43021), .B(n43095), .Y(n47181) );
  NAND2X1 U49295 ( .A(n2250), .B(n43362), .Y(n47184) );
  NAND2X1 U49296 ( .A(n2225), .B(n38406), .Y(n47183) );
  NAND2X1 U49297 ( .A(n47184), .B(n47183), .Y(n47188) );
  NAND2X1 U49298 ( .A(n2232), .B(n43343), .Y(n47186) );
  NAND2X1 U49299 ( .A(n2240), .B(n38602), .Y(n47185) );
  NAND2X1 U49300 ( .A(n47186), .B(n47185), .Y(n47187) );
  NOR2X1 U49301 ( .A(n47188), .B(n47187), .Y(n47196) );
  NAND2X1 U49302 ( .A(n2222), .B(n43030), .Y(n47190) );
  NAND2X1 U49303 ( .A(n2228), .B(n43033), .Y(n47189) );
  NAND2X1 U49304 ( .A(n47190), .B(n47189), .Y(n47194) );
  NAND2X1 U49305 ( .A(n2242), .B(n38534), .Y(n47192) );
  NAND2X1 U49306 ( .A(n2234), .B(n43352), .Y(n47191) );
  NAND2X1 U49307 ( .A(n47192), .B(n47191), .Y(n47193) );
  NOR2X1 U49308 ( .A(n47194), .B(n47193), .Y(n47195) );
  NAND2X1 U49309 ( .A(n47196), .B(n47195), .Y(n47212) );
  NAND2X1 U49310 ( .A(n2238), .B(n43355), .Y(n47198) );
  NAND2X1 U49311 ( .A(n2236), .B(n43039), .Y(n47197) );
  NAND2X1 U49312 ( .A(n47198), .B(n47197), .Y(n47202) );
  NAND2X1 U49313 ( .A(n1793), .B(n39801), .Y(n47200) );
  NAND2X1 U49314 ( .A(n2244), .B(n43043), .Y(n47199) );
  NAND2X1 U49315 ( .A(n47200), .B(n47199), .Y(n47201) );
  NOR2X1 U49316 ( .A(n47202), .B(n47201), .Y(n47210) );
  NAND2X1 U49317 ( .A(n2248), .B(n43359), .Y(n47204) );
  NAND2X1 U49318 ( .A(n2223), .B(n43346), .Y(n47203) );
  NAND2X1 U49319 ( .A(n47204), .B(n47203), .Y(n47208) );
  NAND2X1 U49320 ( .A(n2230), .B(n43339), .Y(n47206) );
  NAND2X1 U49321 ( .A(n2246), .B(n43366), .Y(n47205) );
  NAND2X1 U49322 ( .A(n47206), .B(n47205), .Y(n47207) );
  NOR2X1 U49323 ( .A(n47208), .B(n47207), .Y(n47209) );
  NAND2X1 U49324 ( .A(n47210), .B(n47209), .Y(n47211) );
  NOR2X1 U49325 ( .A(n47212), .B(n47211), .Y(n47242) );
  NAND2X1 U49326 ( .A(n2243), .B(n40273), .Y(n47214) );
  NAND2X1 U49327 ( .A(n2249), .B(n43048), .Y(n47213) );
  NAND2X1 U49328 ( .A(n47214), .B(n47213), .Y(n47218) );
  NAND2X1 U49329 ( .A(n2241), .B(n43050), .Y(n47216) );
  NAND2X1 U49330 ( .A(n2227), .B(n43052), .Y(n47215) );
  NAND2X1 U49331 ( .A(n47216), .B(n47215), .Y(n47217) );
  NOR2X1 U49332 ( .A(n47218), .B(n47217), .Y(n47224) );
  NOR2X1 U49333 ( .A(n43371), .B(n36890), .Y(n47222) );
  NAND2X1 U49334 ( .A(n2229), .B(n38577), .Y(n47220) );
  NAND2X1 U49335 ( .A(n1794), .B(n43057), .Y(n47219) );
  NAND2X1 U49336 ( .A(n47220), .B(n47219), .Y(n47221) );
  NOR2X1 U49337 ( .A(n47222), .B(n47221), .Y(n47223) );
  NAND2X1 U49338 ( .A(n47224), .B(n47223), .Y(n47240) );
  NAND2X1 U49339 ( .A(n2247), .B(n43061), .Y(n47226) );
  NAND2X1 U49340 ( .A(n2245), .B(n39139), .Y(n47225) );
  NAND2X1 U49341 ( .A(n47226), .B(n47225), .Y(n47230) );
  NAND2X1 U49342 ( .A(n2237), .B(n40158), .Y(n47228) );
  NAND2X1 U49343 ( .A(n2226), .B(n43067), .Y(n47227) );
  NAND2X1 U49344 ( .A(n47228), .B(n47227), .Y(n47229) );
  NOR2X1 U49345 ( .A(n47230), .B(n47229), .Y(n47238) );
  NAND2X1 U49346 ( .A(n2233), .B(n38528), .Y(n47232) );
  NAND2X1 U49347 ( .A(n2239), .B(n43350), .Y(n47231) );
  NAND2X1 U49348 ( .A(n47232), .B(n47231), .Y(n47236) );
  NAND2X1 U49349 ( .A(n2231), .B(n43069), .Y(n47234) );
  NAND2X1 U49350 ( .A(n2224), .B(n43072), .Y(n47233) );
  NAND2X1 U49351 ( .A(n47234), .B(n47233), .Y(n47235) );
  NOR2X1 U49352 ( .A(n47236), .B(n47235), .Y(n47237) );
  NAND2X1 U49353 ( .A(n47238), .B(n47237), .Y(n47239) );
  NOR2X1 U49354 ( .A(n47240), .B(n47239), .Y(n47241) );
  NAND2X1 U49355 ( .A(n47242), .B(n47241), .Y(n47243) );
  NOR2X1 U49356 ( .A(n40862), .B(n37122), .Y(n47245) );
  NOR2X1 U49357 ( .A(n40517), .B(n37127), .Y(n47244) );
  NOR2X1 U49358 ( .A(n47245), .B(n47244), .Y(n47247) );
  NAND2X1 U49359 ( .A(n2224), .B(n42706), .Y(n47246) );
  NAND2X1 U49360 ( .A(n47247), .B(n47246), .Y(n47292) );
  NAND2X1 U49361 ( .A(n2227), .B(n40519), .Y(n47249) );
  NAND2X1 U49362 ( .A(n2241), .B(n42626), .Y(n47248) );
  NAND2X1 U49363 ( .A(n47249), .B(n47248), .Y(n47255) );
  NOR2X1 U49364 ( .A(n42903), .B(n36878), .Y(n47251) );
  NOR2X1 U49365 ( .A(n42904), .B(n36885), .Y(n47250) );
  NOR2X1 U49366 ( .A(n47251), .B(n47250), .Y(n47253) );
  NAND2X1 U49367 ( .A(n1794), .B(n42617), .Y(n47252) );
  NAND2X1 U49368 ( .A(n47253), .B(n47252), .Y(n47254) );
  NOR2X1 U49369 ( .A(n47255), .B(n47254), .Y(n47265) );
  NAND2X1 U49370 ( .A(n2240), .B(n40426), .Y(n47257) );
  NAND2X1 U49371 ( .A(n2242), .B(n40536), .Y(n47256) );
  NAND2X1 U49372 ( .A(n47257), .B(n47256), .Y(n47263) );
  NOR2X1 U49373 ( .A(n42646), .B(n36882), .Y(n47259) );
  NOR2X1 U49374 ( .A(n38213), .B(n36888), .Y(n47258) );
  NOR2X1 U49375 ( .A(n47259), .B(n47258), .Y(n47261) );
  NAND2X1 U49376 ( .A(n2243), .B(n42680), .Y(n47260) );
  NAND2X1 U49377 ( .A(n47261), .B(n47260), .Y(n47262) );
  NOR2X1 U49378 ( .A(n47263), .B(n47262), .Y(n47264) );
  NAND2X1 U49379 ( .A(n47265), .B(n47264), .Y(n47285) );
  NAND2X1 U49380 ( .A(n2232), .B(n42777), .Y(n47267) );
  NAND2X1 U49381 ( .A(n2223), .B(n38709), .Y(n47266) );
  NAND2X1 U49382 ( .A(n47267), .B(n47266), .Y(n47273) );
  NOR2X1 U49383 ( .A(n36609), .B(n36883), .Y(n47269) );
  NOR2X1 U49384 ( .A(n42896), .B(n36890), .Y(n47268) );
  NOR2X1 U49385 ( .A(n47269), .B(n47268), .Y(n47271) );
  NAND2X1 U49386 ( .A(n47271), .B(n47270), .Y(n47272) );
  NOR2X1 U49387 ( .A(n47273), .B(n47272), .Y(n47283) );
  NAND2X1 U49388 ( .A(n2238), .B(n46177), .Y(n47275) );
  NAND2X1 U49389 ( .A(n47275), .B(n47274), .Y(n47281) );
  NOR2X1 U49390 ( .A(n49665), .B(n36889), .Y(n47277) );
  NOR2X1 U49391 ( .A(n40851), .B(n36895), .Y(n47276) );
  NOR2X1 U49392 ( .A(n47277), .B(n47276), .Y(n47279) );
  NAND2X1 U49393 ( .A(n2234), .B(n40515), .Y(n47278) );
  NAND2X1 U49394 ( .A(n47279), .B(n47278), .Y(n47280) );
  NOR2X1 U49395 ( .A(n47281), .B(n47280), .Y(n47282) );
  NAND2X1 U49396 ( .A(n47283), .B(n47282), .Y(n47284) );
  NOR2X1 U49397 ( .A(n47285), .B(n47284), .Y(n47286) );
  NOR2X1 U49398 ( .A(n47286), .B(n42889), .Y(n47288) );
  NOR2X1 U49399 ( .A(n42914), .B(n37188), .Y(n47287) );
  NOR2X1 U49400 ( .A(n47288), .B(n47287), .Y(n47291) );
  NOR2X1 U49401 ( .A(n39335), .B(n37157), .Y(n47290) );
  NOR2X1 U49402 ( .A(n42901), .B(n37161), .Y(n47289) );
  NAND2X1 U49403 ( .A(writeback_exec_value_w[15]), .B(n43020), .Y(n47293) );
  NAND2X1 U49404 ( .A(n47294), .B(n47293), .Y(n47302) );
  NOR2X1 U49405 ( .A(n49710), .B(n37158), .Y(n47296) );
  NOR2X1 U49406 ( .A(n46727), .B(n37163), .Y(n47295) );
  NOR2X1 U49407 ( .A(n47296), .B(n47295), .Y(n47300) );
  NOR2X1 U49408 ( .A(n42911), .B(n37162), .Y(n47298) );
  NOR2X1 U49409 ( .A(n42919), .B(n37167), .Y(n47297) );
  NOR2X1 U49410 ( .A(n47298), .B(n47297), .Y(n47299) );
  NAND2X1 U49411 ( .A(n47300), .B(n47299), .Y(n47301) );
  NAND2X1 U49412 ( .A(n43895), .B(n43787), .Y(n57828) );
  NAND2X1 U49413 ( .A(n43789), .B(n43890), .Y(n57830) );
  NOR2X1 U49414 ( .A(n42908), .B(n37173), .Y(n47303) );
  NAND2X1 U49415 ( .A(n3015), .B(n49647), .Y(n47304) );
  NAND2X1 U49416 ( .A(n47305), .B(n47304), .Y(n47346) );
  NAND2X1 U49417 ( .A(n3018), .B(n49674), .Y(n47307) );
  NAND2X1 U49418 ( .A(n3032), .B(n42627), .Y(n47306) );
  NAND2X1 U49419 ( .A(n47307), .B(n47306), .Y(n47313) );
  NOR2X1 U49420 ( .A(n45640), .B(n36847), .Y(n47309) );
  NOR2X1 U49421 ( .A(n38753), .B(n36857), .Y(n47308) );
  NOR2X1 U49422 ( .A(n47309), .B(n47308), .Y(n47311) );
  NAND2X1 U49423 ( .A(n1798), .B(n42620), .Y(n47310) );
  NAND2X1 U49424 ( .A(n47311), .B(n47310), .Y(n47312) );
  NOR2X1 U49425 ( .A(n47313), .B(n47312), .Y(n47323) );
  NAND2X1 U49426 ( .A(n3031), .B(n40424), .Y(n47315) );
  NAND2X1 U49427 ( .A(n47315), .B(n47314), .Y(n47321) );
  NOR2X1 U49428 ( .A(n42646), .B(n36854), .Y(n47317) );
  NOR2X1 U49429 ( .A(n42858), .B(n36859), .Y(n47316) );
  NOR2X1 U49430 ( .A(n47317), .B(n47316), .Y(n47319) );
  NAND2X1 U49431 ( .A(n3034), .B(n42680), .Y(n47318) );
  NAND2X1 U49432 ( .A(n47319), .B(n47318), .Y(n47320) );
  NOR2X1 U49433 ( .A(n47321), .B(n47320), .Y(n47322) );
  NAND2X1 U49434 ( .A(n47323), .B(n47322), .Y(n47339) );
  NAND2X1 U49435 ( .A(n3023), .B(n42779), .Y(n47325) );
  NAND2X1 U49436 ( .A(n3014), .B(n38709), .Y(n47324) );
  NAND2X1 U49437 ( .A(n47325), .B(n47324), .Y(n47331) );
  NOR2X1 U49438 ( .A(n42891), .B(n36858), .Y(n47327) );
  NOR2X1 U49439 ( .A(n45651), .B(n36864), .Y(n47326) );
  NOR2X1 U49440 ( .A(n47327), .B(n47326), .Y(n47329) );
  NAND2X1 U49441 ( .A(n47329), .B(n47328), .Y(n47330) );
  NAND2X1 U49442 ( .A(n3029), .B(n57615), .Y(n47333) );
  NAND2X1 U49443 ( .A(n47333), .B(n47332), .Y(n47337) );
  NOR2X1 U49444 ( .A(n49400), .B(n36863), .Y(n47335) );
  NOR2X1 U49445 ( .A(n42894), .B(n36869), .Y(n47334) );
  NOR2X1 U49446 ( .A(n42916), .B(n37176), .Y(n47340) );
  NOR2X1 U49447 ( .A(n47340), .B(n47341), .Y(n47344) );
  NOR2X1 U49448 ( .A(n39335), .B(n37174), .Y(n47342) );
  NAND2X1 U49449 ( .A(n47343), .B(n47344), .Y(n47345) );
  NAND2X1 U49450 ( .A(mem_d_data_rd_i[14]), .B(n31921), .Y(n47347) );
  NAND2X1 U49451 ( .A(n34489), .B(n47347), .Y(n47348) );
  NAND2X1 U49452 ( .A(writeback_exec_value_w[14]), .B(n43020), .Y(n47349) );
  NAND2X1 U49453 ( .A(n47350), .B(n47349), .Y(n47358) );
  NOR2X1 U49454 ( .A(n42909), .B(n37175), .Y(n47352) );
  NOR2X1 U49455 ( .A(n46727), .B(n37179), .Y(n47351) );
  NOR2X1 U49456 ( .A(n47352), .B(n47351), .Y(n47356) );
  NOR2X1 U49457 ( .A(n49637), .B(n37177), .Y(n47354) );
  NOR2X1 U49458 ( .A(n42917), .B(n37181), .Y(n47353) );
  NOR2X1 U49459 ( .A(n47354), .B(n47353), .Y(n47355) );
  NAND2X1 U49460 ( .A(n47356), .B(n47355), .Y(n47357) );
  NOR2X1 U49461 ( .A(n43142), .B(n43455), .Y(n47360) );
  NOR2X1 U49462 ( .A(n43021), .B(n43145), .Y(n47359) );
  NAND2X1 U49463 ( .A(n3041), .B(n43361), .Y(n47362) );
  NAND2X1 U49464 ( .A(n3016), .B(n38413), .Y(n47361) );
  NAND2X1 U49465 ( .A(n47362), .B(n47361), .Y(n47366) );
  NAND2X1 U49466 ( .A(n3023), .B(n38401), .Y(n47364) );
  NAND2X1 U49467 ( .A(n3031), .B(n38602), .Y(n47363) );
  NAND2X1 U49468 ( .A(n47364), .B(n47363), .Y(n47365) );
  NOR2X1 U49469 ( .A(n47366), .B(n47365), .Y(n47374) );
  NAND2X1 U49470 ( .A(n3013), .B(n38599), .Y(n47368) );
  NAND2X1 U49471 ( .A(n3019), .B(n43033), .Y(n47367) );
  NAND2X1 U49472 ( .A(n47368), .B(n47367), .Y(n47372) );
  NAND2X1 U49473 ( .A(n3033), .B(n38534), .Y(n47370) );
  NAND2X1 U49474 ( .A(n3025), .B(n43352), .Y(n47369) );
  NAND2X1 U49475 ( .A(n47370), .B(n47369), .Y(n47371) );
  NOR2X1 U49476 ( .A(n47372), .B(n47371), .Y(n47373) );
  NAND2X1 U49477 ( .A(n47374), .B(n47373), .Y(n47390) );
  NAND2X1 U49478 ( .A(n3029), .B(n43355), .Y(n47376) );
  NAND2X1 U49479 ( .A(n3027), .B(n40169), .Y(n47375) );
  NAND2X1 U49480 ( .A(n47376), .B(n47375), .Y(n47380) );
  NAND2X1 U49481 ( .A(n1796), .B(n39808), .Y(n47378) );
  NAND2X1 U49482 ( .A(n3035), .B(n43043), .Y(n47377) );
  NAND2X1 U49483 ( .A(n47378), .B(n47377), .Y(n47379) );
  NOR2X1 U49484 ( .A(n47380), .B(n47379), .Y(n47388) );
  NAND2X1 U49485 ( .A(n3039), .B(n38389), .Y(n47382) );
  NAND2X1 U49486 ( .A(n3014), .B(n43346), .Y(n47381) );
  NAND2X1 U49487 ( .A(n47382), .B(n47381), .Y(n47386) );
  NAND2X1 U49488 ( .A(n3021), .B(n43339), .Y(n47384) );
  NAND2X1 U49489 ( .A(n3037), .B(n43366), .Y(n47383) );
  NAND2X1 U49490 ( .A(n47384), .B(n47383), .Y(n47385) );
  NOR2X1 U49491 ( .A(n47386), .B(n47385), .Y(n47387) );
  NAND2X1 U49492 ( .A(n47388), .B(n47387), .Y(n47389) );
  NOR2X1 U49493 ( .A(n47390), .B(n47389), .Y(n47420) );
  NAND2X1 U49494 ( .A(n3034), .B(n40273), .Y(n47392) );
  NAND2X1 U49495 ( .A(n3040), .B(n43048), .Y(n47391) );
  NAND2X1 U49496 ( .A(n47392), .B(n47391), .Y(n47396) );
  NAND2X1 U49497 ( .A(n3032), .B(n43050), .Y(n47394) );
  NAND2X1 U49498 ( .A(n3018), .B(n43052), .Y(n47393) );
  NAND2X1 U49499 ( .A(n47394), .B(n47393), .Y(n47395) );
  NOR2X1 U49500 ( .A(n47396), .B(n47395), .Y(n47402) );
  NOR2X1 U49501 ( .A(n43370), .B(n36864), .Y(n47400) );
  NAND2X1 U49502 ( .A(n3020), .B(n38577), .Y(n47398) );
  NAND2X1 U49503 ( .A(n1798), .B(n40026), .Y(n47397) );
  NAND2X1 U49504 ( .A(n47398), .B(n47397), .Y(n47399) );
  NOR2X1 U49505 ( .A(n47400), .B(n47399), .Y(n47401) );
  NAND2X1 U49506 ( .A(n47402), .B(n47401), .Y(n47418) );
  NAND2X1 U49507 ( .A(n3038), .B(n43061), .Y(n47404) );
  NAND2X1 U49508 ( .A(n3036), .B(n39139), .Y(n47403) );
  NAND2X1 U49509 ( .A(n47404), .B(n47403), .Y(n47408) );
  NAND2X1 U49510 ( .A(n3028), .B(n40158), .Y(n47406) );
  NAND2X1 U49511 ( .A(n3017), .B(n38573), .Y(n47405) );
  NAND2X1 U49512 ( .A(n47406), .B(n47405), .Y(n47407) );
  NOR2X1 U49513 ( .A(n47408), .B(n47407), .Y(n47416) );
  NAND2X1 U49514 ( .A(n3024), .B(n38528), .Y(n47410) );
  NAND2X1 U49515 ( .A(n3030), .B(n43349), .Y(n47409) );
  NAND2X1 U49516 ( .A(n47410), .B(n47409), .Y(n47414) );
  NAND2X1 U49517 ( .A(n3022), .B(n43069), .Y(n47412) );
  NAND2X1 U49518 ( .A(n3015), .B(n43072), .Y(n47411) );
  NAND2X1 U49519 ( .A(n47412), .B(n47411), .Y(n47413) );
  NOR2X1 U49520 ( .A(n47414), .B(n47413), .Y(n47415) );
  NAND2X1 U49521 ( .A(n47416), .B(n47415), .Y(n47417) );
  NOR2X1 U49522 ( .A(n47418), .B(n47417), .Y(n47419) );
  NAND2X1 U49523 ( .A(n47420), .B(n47419), .Y(n47421) );
  NAND2X1 U49524 ( .A(n43722), .B(n43879), .Y(n57811) );
  NAND2X1 U49525 ( .A(n57830), .B(n57811), .Y(n57814) );
  INVX1 U49526 ( .A(n57814), .Y(n73435) );
  NOR2X1 U49527 ( .A(n49625), .B(n37252), .Y(n47424) );
  NAND2X1 U49528 ( .A(n42149), .B(n47422), .Y(n49169) );
  NOR2X1 U49529 ( .A(n49169), .B(n37258), .Y(n47423) );
  NOR2X1 U49530 ( .A(n47424), .B(n47423), .Y(n47426) );
  NAND2X1 U49531 ( .A(n2422), .B(n42706), .Y(n47425) );
  NAND2X1 U49532 ( .A(n47426), .B(n47425), .Y(n47473) );
  NAND2X1 U49533 ( .A(n2425), .B(n40519), .Y(n47428) );
  NAND2X1 U49534 ( .A(n2439), .B(n42625), .Y(n47427) );
  NAND2X1 U49535 ( .A(n47428), .B(n47427), .Y(n47434) );
  NOR2X1 U49536 ( .A(n45640), .B(n37076), .Y(n47430) );
  NOR2X1 U49537 ( .A(n42904), .B(n37083), .Y(n47429) );
  NOR2X1 U49538 ( .A(n47430), .B(n47429), .Y(n47432) );
  NAND2X1 U49539 ( .A(n2449), .B(n42617), .Y(n47431) );
  NAND2X1 U49540 ( .A(n47432), .B(n47431), .Y(n47433) );
  NOR2X1 U49541 ( .A(n47434), .B(n47433), .Y(n47444) );
  NAND2X1 U49542 ( .A(n2438), .B(n40426), .Y(n47436) );
  NAND2X1 U49543 ( .A(n2440), .B(n40536), .Y(n47435) );
  NAND2X1 U49544 ( .A(n47436), .B(n47435), .Y(n47442) );
  NOR2X1 U49545 ( .A(n42864), .B(n37080), .Y(n47438) );
  NOR2X1 U49546 ( .A(n38213), .B(n37086), .Y(n47437) );
  NOR2X1 U49547 ( .A(n47438), .B(n47437), .Y(n47440) );
  NAND2X1 U49548 ( .A(n2441), .B(n42678), .Y(n47439) );
  NAND2X1 U49549 ( .A(n47440), .B(n47439), .Y(n47441) );
  NOR2X1 U49550 ( .A(n47442), .B(n47441), .Y(n47443) );
  NAND2X1 U49551 ( .A(n47444), .B(n47443), .Y(n47464) );
  NAND2X1 U49552 ( .A(n2430), .B(n42779), .Y(n47446) );
  NAND2X1 U49553 ( .A(n47446), .B(n47445), .Y(n47452) );
  NOR2X1 U49554 ( .A(n36609), .B(n37082), .Y(n47448) );
  NOR2X1 U49555 ( .A(n42896), .B(n37087), .Y(n47447) );
  NOR2X1 U49556 ( .A(n47448), .B(n47447), .Y(n47450) );
  NAND2X1 U49557 ( .A(n2428), .B(n73368), .Y(n47449) );
  NAND2X1 U49558 ( .A(n47450), .B(n47449), .Y(n47451) );
  NOR2X1 U49559 ( .A(n47452), .B(n47451), .Y(n47462) );
  NAND2X1 U49560 ( .A(n2436), .B(n57615), .Y(n47454) );
  NAND2X1 U49561 ( .A(n2431), .B(n40537), .Y(n47453) );
  NAND2X1 U49562 ( .A(n47454), .B(n47453), .Y(n47460) );
  NOR2X1 U49563 ( .A(n45507), .B(n37088), .Y(n47456) );
  NOR2X1 U49564 ( .A(n40497), .B(n37090), .Y(n47455) );
  NOR2X1 U49565 ( .A(n47456), .B(n47455), .Y(n47458) );
  NAND2X1 U49566 ( .A(n2432), .B(n40515), .Y(n47457) );
  NAND2X1 U49567 ( .A(n47458), .B(n47457), .Y(n47459) );
  NOR2X1 U49568 ( .A(n47460), .B(n47459), .Y(n47461) );
  NAND2X1 U49569 ( .A(n47462), .B(n47461), .Y(n47463) );
  NOR2X1 U49570 ( .A(n47464), .B(n47463), .Y(n47465) );
  NOR2X1 U49571 ( .A(n47465), .B(n42889), .Y(n47467) );
  NOR2X1 U49572 ( .A(n42916), .B(n37266), .Y(n47466) );
  NOR2X1 U49573 ( .A(n47467), .B(n47466), .Y(n47471) );
  NOR2X1 U49574 ( .A(n40277), .B(n37263), .Y(n47469) );
  NOR2X1 U49575 ( .A(n39572), .B(n37268), .Y(n47468) );
  NOR2X1 U49576 ( .A(n47469), .B(n47468), .Y(n47470) );
  NAND2X1 U49577 ( .A(n47471), .B(n47470), .Y(n47472) );
  NOR2X1 U49578 ( .A(n42900), .B(n37259), .Y(n47477) );
  INVX1 U49579 ( .A(n31923), .Y(n73578) );
  NAND2X1 U49580 ( .A(mem_d_data_rd_i[25]), .B(n73578), .Y(n47474) );
  NAND2X1 U49581 ( .A(n34489), .B(n47474), .Y(n47475) );
  NOR2X1 U49582 ( .A(n43120), .B(n40360), .Y(n47476) );
  NOR2X1 U49583 ( .A(n47477), .B(n47476), .Y(n47479) );
  NAND2X1 U49584 ( .A(writeback_exec_value_w[9]), .B(n37976), .Y(n47478) );
  NAND2X1 U49585 ( .A(n47479), .B(n47478), .Y(n47487) );
  NOR2X1 U49586 ( .A(n42910), .B(n37264), .Y(n47481) );
  NOR2X1 U49587 ( .A(n38932), .B(n37269), .Y(n47480) );
  NOR2X1 U49588 ( .A(n47481), .B(n47480), .Y(n47485) );
  NOR2X1 U49589 ( .A(n49637), .B(n37267), .Y(n47483) );
  NOR2X1 U49590 ( .A(n42918), .B(n37270), .Y(n47482) );
  NOR2X1 U49591 ( .A(n47483), .B(n47482), .Y(n47484) );
  NAND2X1 U49592 ( .A(n47485), .B(n47484), .Y(n47486) );
  NOR2X1 U49593 ( .A(n43120), .B(n43455), .Y(n47489) );
  NOR2X1 U49594 ( .A(n43021), .B(n43123), .Y(n47488) );
  NOR2X1 U49595 ( .A(n47489), .B(n47488), .Y(n47552) );
  NAND2X1 U49596 ( .A(n2448), .B(n43361), .Y(n47491) );
  NAND2X1 U49597 ( .A(n2424), .B(n38409), .Y(n47490) );
  NAND2X1 U49598 ( .A(n47491), .B(n47490), .Y(n47495) );
  NAND2X1 U49599 ( .A(n2430), .B(n38401), .Y(n47493) );
  NAND2X1 U49600 ( .A(n2438), .B(n43028), .Y(n47492) );
  NAND2X1 U49601 ( .A(n47493), .B(n47492), .Y(n47494) );
  NOR2X1 U49602 ( .A(n47495), .B(n47494), .Y(n47503) );
  NAND2X1 U49603 ( .A(n1826), .B(n38599), .Y(n47497) );
  NAND2X1 U49604 ( .A(n2426), .B(n43033), .Y(n47496) );
  NAND2X1 U49605 ( .A(n47497), .B(n47496), .Y(n47501) );
  NAND2X1 U49606 ( .A(n2440), .B(n43037), .Y(n47499) );
  NAND2X1 U49607 ( .A(n2432), .B(n43352), .Y(n47498) );
  NAND2X1 U49608 ( .A(n47499), .B(n47498), .Y(n47500) );
  NOR2X1 U49609 ( .A(n47501), .B(n47500), .Y(n47502) );
  NAND2X1 U49610 ( .A(n47503), .B(n47502), .Y(n47519) );
  NAND2X1 U49611 ( .A(n2436), .B(n43356), .Y(n47505) );
  NAND2X1 U49612 ( .A(n2434), .B(n40169), .Y(n47504) );
  NAND2X1 U49613 ( .A(n47505), .B(n47504), .Y(n47509) );
  NAND2X1 U49614 ( .A(n2450), .B(n39807), .Y(n47507) );
  NAND2X1 U49615 ( .A(n2442), .B(n43043), .Y(n47506) );
  NAND2X1 U49616 ( .A(n47507), .B(n47506), .Y(n47508) );
  NOR2X1 U49617 ( .A(n47509), .B(n47508), .Y(n47517) );
  NAND2X1 U49618 ( .A(n2446), .B(n38389), .Y(n47511) );
  NAND2X1 U49619 ( .A(n2421), .B(n43346), .Y(n47510) );
  NAND2X1 U49620 ( .A(n47511), .B(n47510), .Y(n47515) );
  NAND2X1 U49621 ( .A(n2428), .B(n43339), .Y(n47513) );
  NAND2X1 U49622 ( .A(n2444), .B(n43366), .Y(n47512) );
  NAND2X1 U49623 ( .A(n47513), .B(n47512), .Y(n47514) );
  NOR2X1 U49624 ( .A(n47515), .B(n47514), .Y(n47516) );
  NAND2X1 U49625 ( .A(n47517), .B(n47516), .Y(n47518) );
  NOR2X1 U49626 ( .A(n47519), .B(n47518), .Y(n47549) );
  NAND2X1 U49627 ( .A(n2441), .B(n40273), .Y(n47521) );
  NAND2X1 U49628 ( .A(n2447), .B(n43048), .Y(n47520) );
  NAND2X1 U49629 ( .A(n47521), .B(n47520), .Y(n47525) );
  NAND2X1 U49630 ( .A(n2439), .B(n49841), .Y(n47523) );
  NAND2X1 U49631 ( .A(n2425), .B(n43052), .Y(n47522) );
  NAND2X1 U49632 ( .A(n47523), .B(n47522), .Y(n47524) );
  NOR2X1 U49633 ( .A(n47525), .B(n47524), .Y(n47531) );
  NOR2X1 U49634 ( .A(n43371), .B(n37087), .Y(n47529) );
  NAND2X1 U49635 ( .A(n2427), .B(n43055), .Y(n47527) );
  NAND2X1 U49636 ( .A(n2449), .B(n40026), .Y(n47526) );
  NAND2X1 U49637 ( .A(n47527), .B(n47526), .Y(n47528) );
  NOR2X1 U49638 ( .A(n47529), .B(n47528), .Y(n47530) );
  NAND2X1 U49639 ( .A(n47531), .B(n47530), .Y(n47547) );
  NAND2X1 U49640 ( .A(n2445), .B(n43061), .Y(n47533) );
  NAND2X1 U49641 ( .A(n2443), .B(n39135), .Y(n47532) );
  NAND2X1 U49642 ( .A(n47533), .B(n47532), .Y(n47537) );
  NAND2X1 U49643 ( .A(n2435), .B(n40158), .Y(n47535) );
  NAND2X1 U49644 ( .A(n2423), .B(n38573), .Y(n47534) );
  NAND2X1 U49645 ( .A(n47535), .B(n47534), .Y(n47536) );
  NOR2X1 U49646 ( .A(n47537), .B(n47536), .Y(n47545) );
  NAND2X1 U49647 ( .A(n2431), .B(n43373), .Y(n47539) );
  NAND2X1 U49648 ( .A(n2437), .B(n43350), .Y(n47538) );
  NAND2X1 U49649 ( .A(n47539), .B(n47538), .Y(n47543) );
  NAND2X1 U49650 ( .A(n2429), .B(n43069), .Y(n47541) );
  NAND2X1 U49651 ( .A(n2422), .B(n43072), .Y(n47540) );
  NAND2X1 U49652 ( .A(n47541), .B(n47540), .Y(n47542) );
  NOR2X1 U49653 ( .A(n47543), .B(n47542), .Y(n47544) );
  NAND2X1 U49654 ( .A(n47545), .B(n47544), .Y(n47546) );
  NOR2X1 U49655 ( .A(n47547), .B(n47546), .Y(n47548) );
  NAND2X1 U49656 ( .A(n47549), .B(n47548), .Y(n47550) );
  NAND2X1 U49657 ( .A(n42804), .B(n47550), .Y(n47551) );
  NOR2X1 U49658 ( .A(n42907), .B(n36899), .Y(n47554) );
  NOR2X1 U49659 ( .A(n40042), .B(n36900), .Y(n47553) );
  NOR2X1 U49660 ( .A(n47554), .B(n47553), .Y(n47556) );
  NAND2X1 U49661 ( .A(n2039), .B(n49647), .Y(n47555) );
  NAND2X1 U49662 ( .A(n47556), .B(n47555), .Y(n47603) );
  NAND2X1 U49663 ( .A(n2041), .B(n40520), .Y(n47558) );
  NAND2X1 U49664 ( .A(n2055), .B(n42626), .Y(n47557) );
  NAND2X1 U49665 ( .A(n47558), .B(n47557), .Y(n47564) );
  NOR2X1 U49666 ( .A(n42902), .B(n36905), .Y(n47560) );
  NOR2X1 U49667 ( .A(n42904), .B(n36893), .Y(n47559) );
  NOR2X1 U49668 ( .A(n47560), .B(n47559), .Y(n47562) );
  NAND2X1 U49669 ( .A(n2065), .B(n42618), .Y(n47561) );
  NAND2X1 U49670 ( .A(n47562), .B(n47561), .Y(n47563) );
  NOR2X1 U49671 ( .A(n47564), .B(n47563), .Y(n47574) );
  NAND2X1 U49672 ( .A(n2054), .B(n40424), .Y(n47566) );
  NAND2X1 U49673 ( .A(n2056), .B(n49685), .Y(n47565) );
  NAND2X1 U49674 ( .A(n47566), .B(n47565), .Y(n47572) );
  NOR2X1 U49675 ( .A(n42864), .B(n37140), .Y(n47568) );
  NOR2X1 U49676 ( .A(n38213), .B(n36903), .Y(n47567) );
  NOR2X1 U49677 ( .A(n47568), .B(n47567), .Y(n47570) );
  NAND2X1 U49678 ( .A(n2057), .B(n42680), .Y(n47569) );
  NAND2X1 U49679 ( .A(n47570), .B(n47569), .Y(n47571) );
  NOR2X1 U49680 ( .A(n47572), .B(n47571), .Y(n47573) );
  NAND2X1 U49681 ( .A(n47574), .B(n47573), .Y(n47594) );
  NAND2X1 U49682 ( .A(n2046), .B(n42779), .Y(n47576) );
  NAND2X1 U49683 ( .A(n2037), .B(n38709), .Y(n47575) );
  NAND2X1 U49684 ( .A(n47576), .B(n47575), .Y(n47582) );
  NOR2X1 U49685 ( .A(n36609), .B(n37032), .Y(n47578) );
  NOR2X1 U49686 ( .A(n42895), .B(n37093), .Y(n47577) );
  NOR2X1 U49687 ( .A(n47578), .B(n47577), .Y(n47580) );
  NAND2X1 U49688 ( .A(n2044), .B(n42675), .Y(n47579) );
  NAND2X1 U49689 ( .A(n47580), .B(n47579), .Y(n47581) );
  NOR2X1 U49690 ( .A(n47582), .B(n47581), .Y(n47592) );
  NAND2X1 U49691 ( .A(n2052), .B(n42781), .Y(n47584) );
  NAND2X1 U49692 ( .A(n2047), .B(n39318), .Y(n47583) );
  NAND2X1 U49693 ( .A(n47584), .B(n47583), .Y(n47590) );
  NOR2X1 U49694 ( .A(n49665), .B(n36897), .Y(n47586) );
  NOR2X1 U49695 ( .A(n40497), .B(n37147), .Y(n47585) );
  NOR2X1 U49696 ( .A(n47586), .B(n47585), .Y(n47588) );
  NAND2X1 U49697 ( .A(n2048), .B(n40515), .Y(n47587) );
  NAND2X1 U49698 ( .A(n47588), .B(n47587), .Y(n47589) );
  NOR2X1 U49699 ( .A(n47590), .B(n47589), .Y(n47591) );
  NAND2X1 U49700 ( .A(n47592), .B(n47591), .Y(n47593) );
  NOR2X1 U49701 ( .A(n47594), .B(n47593), .Y(n47595) );
  NOR2X1 U49702 ( .A(n47595), .B(n42890), .Y(n47597) );
  NOR2X1 U49703 ( .A(n42915), .B(n36898), .Y(n47596) );
  NOR2X1 U49704 ( .A(n47597), .B(n47596), .Y(n47601) );
  NOR2X1 U49705 ( .A(n39335), .B(n37028), .Y(n47599) );
  NOR2X1 U49706 ( .A(n39572), .B(n36913), .Y(n47598) );
  NOR2X1 U49707 ( .A(n47599), .B(n47598), .Y(n47600) );
  NAND2X1 U49708 ( .A(n47601), .B(n47600), .Y(n47602) );
  NOR2X1 U49709 ( .A(n39353), .B(n37092), .Y(n47607) );
  NOR2X1 U49710 ( .A(n34083), .B(n34082), .Y(n47605) );
  NOR2X1 U49711 ( .A(n34081), .B(n34080), .Y(n47604) );
  NAND2X1 U49712 ( .A(n47605), .B(n47604), .Y(n47618) );
  NOR2X1 U49713 ( .A(n43074), .B(n42899), .Y(n47606) );
  NOR2X1 U49714 ( .A(n47607), .B(n47606), .Y(n47609) );
  NAND2X1 U49715 ( .A(writeback_exec_value_w[3]), .B(n43020), .Y(n47608) );
  NAND2X1 U49716 ( .A(n47609), .B(n47608), .Y(n47617) );
  NOR2X1 U49717 ( .A(n49710), .B(n37024), .Y(n47611) );
  NOR2X1 U49718 ( .A(n38932), .B(n37091), .Y(n47610) );
  NOR2X1 U49719 ( .A(n47611), .B(n47610), .Y(n47615) );
  NOR2X1 U49720 ( .A(n40855), .B(n37026), .Y(n47613) );
  NOR2X1 U49721 ( .A(n42919), .B(n36902), .Y(n47612) );
  NOR2X1 U49722 ( .A(n47613), .B(n47612), .Y(n47614) );
  NAND2X1 U49723 ( .A(n47615), .B(n47614), .Y(n47616) );
  NAND2X1 U49724 ( .A(writeback_exec_value_w[3]), .B(n43025), .Y(n47620) );
  NAND2X1 U49725 ( .A(n38271), .B(n47618), .Y(n47619) );
  NOR2X1 U49726 ( .A(n48360), .B(n37024), .Y(n47623) );
  NOR2X1 U49727 ( .A(n57625), .B(n37032), .Y(n47622) );
  NOR2X1 U49728 ( .A(n47623), .B(n47622), .Y(n47629) );
  NOR2X1 U49729 ( .A(n47624), .B(n37026), .Y(n47627) );
  NOR2X1 U49730 ( .A(n47625), .B(n37040), .Y(n47626) );
  NOR2X1 U49731 ( .A(n47627), .B(n47626), .Y(n47628) );
  NAND2X1 U49732 ( .A(n47629), .B(n47628), .Y(n47643) );
  NOR2X1 U49733 ( .A(n57609), .B(n37028), .Y(n47635) );
  NOR2X1 U49734 ( .A(n43015), .B(n38366), .Y(n47630) );
  NAND2X1 U49735 ( .A(n47630), .B(n2037), .Y(n47633) );
  NOR2X1 U49736 ( .A(n42670), .B(n42869), .Y(n47631) );
  NAND2X1 U49737 ( .A(n47631), .B(n2040), .Y(n47632) );
  NAND2X1 U49738 ( .A(n47633), .B(n47632), .Y(n47634) );
  NOR2X1 U49739 ( .A(n47635), .B(n47634), .Y(n47641) );
  NOR2X1 U49740 ( .A(n47636), .B(n37039), .Y(n47639) );
  NOR2X1 U49741 ( .A(n47637), .B(n37047), .Y(n47638) );
  NOR2X1 U49742 ( .A(n47639), .B(n47638), .Y(n47640) );
  NAND2X1 U49743 ( .A(n47641), .B(n47640), .Y(n47642) );
  NOR2X1 U49744 ( .A(n47643), .B(n47642), .Y(n47702) );
  NAND2X1 U49745 ( .A(n48199), .B(n39669), .Y(n47644) );
  NOR2X1 U49746 ( .A(n36893), .B(n47644), .Y(n47646) );
  NOR2X1 U49747 ( .A(n47646), .B(n47645), .Y(n47652) );
  NAND2X1 U49748 ( .A(n48205), .B(n39669), .Y(n47647) );
  NOR2X1 U49749 ( .A(n36897), .B(n47647), .Y(n47650) );
  NAND2X1 U49750 ( .A(n42743), .B(n43019), .Y(n47648) );
  NOR2X1 U49751 ( .A(n36904), .B(n47648), .Y(n47649) );
  NOR2X1 U49752 ( .A(n47650), .B(n47649), .Y(n47651) );
  NAND2X1 U49753 ( .A(n47652), .B(n47651), .Y(n47663) );
  NAND2X1 U49754 ( .A(n40448), .B(n42757), .Y(n47653) );
  NOR2X1 U49755 ( .A(n36900), .B(n47653), .Y(n47656) );
  NAND2X1 U49756 ( .A(n47674), .B(n48372), .Y(n47654) );
  NOR2X1 U49757 ( .A(n36905), .B(n47654), .Y(n47655) );
  NOR2X1 U49758 ( .A(n47656), .B(n47655), .Y(n47661) );
  NAND2X1 U49759 ( .A(n47674), .B(n58130), .Y(n47657) );
  NOR2X1 U49760 ( .A(n36909), .B(n47657), .Y(n47658) );
  NOR2X1 U49761 ( .A(n47659), .B(n47658), .Y(n47660) );
  NAND2X1 U49762 ( .A(n47661), .B(n47660), .Y(n47662) );
  NAND2X1 U49763 ( .A(n48370), .B(n42673), .Y(n47664) );
  NOR2X1 U49764 ( .A(n36898), .B(n47664), .Y(n47667) );
  NAND2X1 U49765 ( .A(n42756), .B(n48370), .Y(n47665) );
  NOR2X1 U49766 ( .A(n36902), .B(n47665), .Y(n47666) );
  NOR2X1 U49767 ( .A(n47667), .B(n47666), .Y(n47673) );
  NAND2X1 U49768 ( .A(n42742), .B(n43018), .Y(n47668) );
  NOR2X1 U49769 ( .A(n36901), .B(n47668), .Y(n47671) );
  NAND2X1 U49770 ( .A(n40448), .B(n43018), .Y(n47669) );
  NOR2X1 U49771 ( .A(n36907), .B(n47669), .Y(n47670) );
  NOR2X1 U49772 ( .A(n47671), .B(n47670), .Y(n47672) );
  NAND2X1 U49773 ( .A(n47673), .B(n47672), .Y(n47684) );
  NAND2X1 U49774 ( .A(n47674), .B(n42673), .Y(n47675) );
  NOR2X1 U49775 ( .A(n36910), .B(n47675), .Y(n47676) );
  NOR2X1 U49776 ( .A(n47677), .B(n47676), .Y(n47682) );
  NAND2X1 U49777 ( .A(n39584), .B(n40076), .Y(n47678) );
  NOR2X1 U49778 ( .A(n36913), .B(n47678), .Y(n47679) );
  NOR2X1 U49779 ( .A(n47680), .B(n47679), .Y(n47681) );
  NAND2X1 U49780 ( .A(n47682), .B(n47681), .Y(n47683) );
  NOR2X1 U49781 ( .A(n47685), .B(n37092), .Y(n47687) );
  NOR2X1 U49782 ( .A(n43369), .B(n37093), .Y(n47686) );
  NOR2X1 U49783 ( .A(n47687), .B(n47686), .Y(n47698) );
  NOR2X1 U49784 ( .A(n37091), .B(n39799), .Y(n47696) );
  NAND2X1 U49785 ( .A(n40448), .B(n39669), .Y(n47688) );
  NOR2X1 U49786 ( .A(n36899), .B(n47688), .Y(n47691) );
  NAND2X1 U49787 ( .A(n42744), .B(n48372), .Y(n47689) );
  NOR2X1 U49788 ( .A(n36903), .B(n47689), .Y(n47690) );
  NOR2X1 U49789 ( .A(n47691), .B(n47690), .Y(n47694) );
  NOR2X1 U49790 ( .A(n43015), .B(n42861), .Y(n47692) );
  NAND2X1 U49791 ( .A(n47692), .B(n2042), .Y(n47693) );
  NAND2X1 U49792 ( .A(n47694), .B(n47693), .Y(n47695) );
  NOR2X1 U49793 ( .A(n47696), .B(n47695), .Y(n47697) );
  NAND2X1 U49794 ( .A(n47698), .B(n47697), .Y(n47699) );
  NOR2X1 U49795 ( .A(n47699), .B(n47700), .Y(n47701) );
  NAND2X1 U49796 ( .A(n47702), .B(n47701), .Y(n47703) );
  NAND2X1 U49797 ( .A(n42804), .B(n47703), .Y(n63825) );
  NAND2X1 U49798 ( .A(n43807), .B(n40392), .Y(n57793) );
  OR2X1 U49799 ( .A(n35166), .B(n35165), .Y(n47705) );
  OR2X1 U49800 ( .A(n35168), .B(n35167), .Y(n47704) );
  NOR2X1 U49801 ( .A(n43329), .B(n47706), .Y(n47707) );
  NOR2X1 U49802 ( .A(n48109), .B(n36482), .Y(n47708) );
  NAND2X1 U49803 ( .A(n2015), .B(n47708), .Y(n47711) );
  NOR2X1 U49804 ( .A(n48109), .B(n42738), .Y(n47709) );
  NAND2X1 U49805 ( .A(n47709), .B(n2018), .Y(n47710) );
  NAND2X1 U49806 ( .A(n47711), .B(n47710), .Y(n47717) );
  NOR2X1 U49807 ( .A(n47965), .B(n36482), .Y(n47712) );
  NAND2X1 U49808 ( .A(n47712), .B(n2031), .Y(n47715) );
  NOR2X1 U49809 ( .A(n48126), .B(n42879), .Y(n47713) );
  NAND2X1 U49810 ( .A(n47713), .B(n2029), .Y(n47714) );
  NAND2X1 U49811 ( .A(n47715), .B(n47714), .Y(n47716) );
  NOR2X1 U49812 ( .A(n47717), .B(n47716), .Y(n47729) );
  NOR2X1 U49813 ( .A(n48116), .B(n42861), .Y(n47718) );
  NAND2X1 U49814 ( .A(n47718), .B(n2033), .Y(n47721) );
  NOR2X1 U49815 ( .A(n48109), .B(n48611), .Y(n47719) );
  NAND2X1 U49816 ( .A(n47719), .B(n2014), .Y(n47720) );
  NAND2X1 U49817 ( .A(n47721), .B(n47720), .Y(n47727) );
  NOR2X1 U49818 ( .A(n48109), .B(n42745), .Y(n47722) );
  NAND2X1 U49819 ( .A(n2016), .B(n47722), .Y(n47725) );
  NOR2X1 U49820 ( .A(n48109), .B(n42880), .Y(n47723) );
  NAND2X1 U49821 ( .A(n2013), .B(n47723), .Y(n47724) );
  NAND2X1 U49822 ( .A(n47725), .B(n47724), .Y(n47726) );
  NOR2X1 U49823 ( .A(n47727), .B(n47726), .Y(n47728) );
  NAND2X1 U49824 ( .A(n47729), .B(n47728), .Y(n47748) );
  NOR2X1 U49825 ( .A(n48585), .B(n42746), .Y(n47730) );
  NAND2X1 U49826 ( .A(n2010), .B(n47730), .Y(n47733) );
  NOR2X1 U49827 ( .A(n48585), .B(n42862), .Y(n47731) );
  NAND2X1 U49828 ( .A(n47731), .B(n2011), .Y(n47732) );
  NAND2X1 U49829 ( .A(n47733), .B(n47732), .Y(n47734) );
  NOR2X1 U49830 ( .A(n42495), .B(n47734), .Y(n47746) );
  NOR2X1 U49831 ( .A(n48116), .B(n48611), .Y(n47735) );
  NAND2X1 U49832 ( .A(n47735), .B(n2030), .Y(n47738) );
  NOR2X1 U49833 ( .A(n48595), .B(n42745), .Y(n47736) );
  NAND2X1 U49834 ( .A(n47736), .B(n2032), .Y(n47737) );
  NAND2X1 U49835 ( .A(n47738), .B(n47737), .Y(n47744) );
  NOR2X1 U49836 ( .A(n48126), .B(n42737), .Y(n47739) );
  NAND2X1 U49837 ( .A(n2034), .B(n47739), .Y(n47742) );
  NOR2X1 U49838 ( .A(n48585), .B(n42737), .Y(n47740) );
  NAND2X1 U49839 ( .A(n47740), .B(n2012), .Y(n47741) );
  NAND2X1 U49840 ( .A(n47742), .B(n47741), .Y(n47743) );
  NOR2X1 U49841 ( .A(n47744), .B(n47743), .Y(n47745) );
  NAND2X1 U49842 ( .A(n47746), .B(n47745), .Y(n47747) );
  NOR2X1 U49843 ( .A(n47748), .B(n47747), .Y(n62915) );
  NOR2X1 U49844 ( .A(n48585), .B(n48611), .Y(n47749) );
  NAND2X1 U49845 ( .A(n2008), .B(n47749), .Y(n47752) );
  NAND2X1 U49846 ( .A(n1832), .B(n40018), .Y(n47750) );
  OR2X1 U49847 ( .A(n48585), .B(n47750), .Y(n47751) );
  NAND2X1 U49848 ( .A(n47752), .B(n47751), .Y(n47758) );
  NOR2X1 U49849 ( .A(n48607), .B(n48611), .Y(n47753) );
  NAND2X1 U49850 ( .A(n47753), .B(n2022), .Y(n47756) );
  NOR2X1 U49851 ( .A(n48607), .B(n42738), .Y(n47754) );
  NAND2X1 U49852 ( .A(n2026), .B(n47754), .Y(n47755) );
  NAND2X1 U49853 ( .A(n47756), .B(n47755), .Y(n47757) );
  NOR2X1 U49854 ( .A(n47758), .B(n47757), .Y(n47770) );
  NOR2X1 U49855 ( .A(n48560), .B(n47965), .Y(n47759) );
  NAND2X1 U49856 ( .A(n47759), .B(n2027), .Y(n47762) );
  NOR2X1 U49857 ( .A(n48585), .B(n42855), .Y(n47760) );
  NAND2X1 U49858 ( .A(n47760), .B(n1831), .Y(n47761) );
  NAND2X1 U49859 ( .A(n47762), .B(n47761), .Y(n47768) );
  NOR2X1 U49860 ( .A(n48585), .B(n38366), .Y(n47763) );
  NAND2X1 U49861 ( .A(n2007), .B(n47763), .Y(n47766) );
  NOR2X1 U49862 ( .A(n48585), .B(n42870), .Y(n47764) );
  NAND2X1 U49863 ( .A(n47764), .B(n2009), .Y(n47765) );
  NAND2X1 U49864 ( .A(n47766), .B(n47765), .Y(n47767) );
  NOR2X1 U49865 ( .A(n47768), .B(n47767), .Y(n47769) );
  NAND2X1 U49866 ( .A(n47770), .B(n47769), .Y(n47794) );
  NAND2X1 U49867 ( .A(n2019), .B(n40018), .Y(n47771) );
  OR2X1 U49868 ( .A(n39883), .B(n47771), .Y(n47774) );
  NOR2X1 U49869 ( .A(n42853), .B(n48595), .Y(n47772) );
  NAND2X1 U49870 ( .A(n47772), .B(n2028), .Y(n47773) );
  NAND2X1 U49871 ( .A(n47774), .B(n47773), .Y(n47780) );
  NOR2X1 U49872 ( .A(n42853), .B(n48109), .Y(n47775) );
  NAND2X1 U49873 ( .A(n47775), .B(n2006), .Y(n47778) );
  NOR2X1 U49874 ( .A(n48109), .B(n42860), .Y(n47776) );
  NAND2X1 U49875 ( .A(n2017), .B(n47776), .Y(n47777) );
  NAND2X1 U49876 ( .A(n47778), .B(n47777), .Y(n47779) );
  NOR2X1 U49877 ( .A(n47780), .B(n47779), .Y(n47792) );
  NOR2X1 U49878 ( .A(n39882), .B(n42860), .Y(n47781) );
  NAND2X1 U49879 ( .A(n2025), .B(n47781), .Y(n47784) );
  NOR2X1 U49880 ( .A(n39883), .B(n42879), .Y(n47782) );
  NAND2X1 U49881 ( .A(n2021), .B(n47782), .Y(n47783) );
  NAND2X1 U49882 ( .A(n47784), .B(n47783), .Y(n47790) );
  NOR2X1 U49883 ( .A(n48607), .B(n42869), .Y(n47785) );
  NAND2X1 U49884 ( .A(n2023), .B(n47785), .Y(n47788) );
  NOR2X1 U49885 ( .A(n39883), .B(n42745), .Y(n47786) );
  NAND2X1 U49886 ( .A(n2024), .B(n47786), .Y(n47787) );
  NAND2X1 U49887 ( .A(n47788), .B(n47787), .Y(n47789) );
  NOR2X1 U49888 ( .A(n47790), .B(n47789), .Y(n47791) );
  NAND2X1 U49889 ( .A(n47792), .B(n47791), .Y(n47793) );
  NOR2X1 U49890 ( .A(n47794), .B(n47793), .Y(n62916) );
  NAND2X1 U49891 ( .A(n62915), .B(n62916), .Y(n63188) );
  NAND2X1 U49892 ( .A(n42802), .B(n63188), .Y(n62460) );
  NOR2X1 U49893 ( .A(n42908), .B(n37305), .Y(n47796) );
  NOR2X1 U49894 ( .A(n49169), .B(n37306), .Y(n47795) );
  NOR2X1 U49895 ( .A(n47796), .B(n47795), .Y(n47798) );
  NAND2X1 U49896 ( .A(n2008), .B(n49647), .Y(n47797) );
  NAND2X1 U49897 ( .A(n47798), .B(n47797), .Y(n47846) );
  NAND2X1 U49898 ( .A(n2010), .B(n40519), .Y(n47800) );
  NAND2X1 U49899 ( .A(n2024), .B(n42627), .Y(n47799) );
  NAND2X1 U49900 ( .A(n47800), .B(n47799), .Y(n47806) );
  NOR2X1 U49901 ( .A(n49677), .B(n37233), .Y(n47802) );
  NOR2X1 U49902 ( .A(n38753), .B(n37236), .Y(n47801) );
  NOR2X1 U49903 ( .A(n47802), .B(n47801), .Y(n47804) );
  NAND2X1 U49904 ( .A(n2034), .B(n42619), .Y(n47803) );
  NAND2X1 U49905 ( .A(n47804), .B(n47803), .Y(n47805) );
  NOR2X1 U49906 ( .A(n47806), .B(n47805), .Y(n47816) );
  NAND2X1 U49907 ( .A(n2023), .B(n40425), .Y(n47808) );
  NAND2X1 U49908 ( .A(n2025), .B(n40535), .Y(n47807) );
  NAND2X1 U49909 ( .A(n47808), .B(n47807), .Y(n47814) );
  NOR2X1 U49910 ( .A(n42647), .B(n37234), .Y(n47810) );
  NOR2X1 U49911 ( .A(n42858), .B(n37237), .Y(n47809) );
  NOR2X1 U49912 ( .A(n47810), .B(n47809), .Y(n47812) );
  NAND2X1 U49913 ( .A(n2026), .B(n42678), .Y(n47811) );
  NAND2X1 U49914 ( .A(n47812), .B(n47811), .Y(n47813) );
  NOR2X1 U49915 ( .A(n47814), .B(n47813), .Y(n47815) );
  NAND2X1 U49916 ( .A(n47816), .B(n47815), .Y(n47836) );
  NAND2X1 U49917 ( .A(n2015), .B(n42777), .Y(n47818) );
  NAND2X1 U49918 ( .A(n2007), .B(n38708), .Y(n47817) );
  NAND2X1 U49919 ( .A(n47818), .B(n47817), .Y(n47824) );
  NOR2X1 U49920 ( .A(n42891), .B(n37235), .Y(n47820) );
  NOR2X1 U49921 ( .A(n42896), .B(n37238), .Y(n47819) );
  NOR2X1 U49922 ( .A(n47820), .B(n47819), .Y(n47822) );
  NAND2X1 U49923 ( .A(n2013), .B(n42675), .Y(n47821) );
  NAND2X1 U49924 ( .A(n47822), .B(n47821), .Y(n47823) );
  NOR2X1 U49925 ( .A(n47824), .B(n47823), .Y(n47834) );
  NAND2X1 U49926 ( .A(n2021), .B(n39645), .Y(n47826) );
  NAND2X1 U49927 ( .A(n2016), .B(n40537), .Y(n47825) );
  NAND2X1 U49928 ( .A(n47826), .B(n47825), .Y(n47832) );
  NOR2X1 U49929 ( .A(n42912), .B(n37239), .Y(n47828) );
  NOR2X1 U49930 ( .A(n42893), .B(n37240), .Y(n47827) );
  NOR2X1 U49931 ( .A(n47828), .B(n47827), .Y(n47830) );
  NAND2X1 U49932 ( .A(n2017), .B(n40514), .Y(n47829) );
  NAND2X1 U49933 ( .A(n47830), .B(n47829), .Y(n47831) );
  NOR2X1 U49934 ( .A(n47832), .B(n47831), .Y(n47833) );
  NAND2X1 U49935 ( .A(n47834), .B(n47833), .Y(n47835) );
  NOR2X1 U49936 ( .A(n47836), .B(n47835), .Y(n47837) );
  NOR2X1 U49937 ( .A(n47837), .B(n42890), .Y(n47840) );
  INVX1 U49938 ( .A(n2020), .Y(n47838) );
  NOR2X1 U49939 ( .A(n42914), .B(n47838), .Y(n47839) );
  NOR2X1 U49940 ( .A(n47840), .B(n47839), .Y(n47844) );
  NOR2X1 U49941 ( .A(n40277), .B(n37309), .Y(n47842) );
  NOR2X1 U49942 ( .A(n49624), .B(n37311), .Y(n47841) );
  NOR2X1 U49943 ( .A(n47842), .B(n47841), .Y(n47843) );
  NAND2X1 U49944 ( .A(n47844), .B(n47843), .Y(n47845) );
  NOR2X1 U49945 ( .A(n47846), .B(n47845), .Y(n47860) );
  NOR2X1 U49946 ( .A(n40406), .B(n37307), .Y(n47848) );
  NOR2X1 U49947 ( .A(n43329), .B(n42898), .Y(n47847) );
  NOR2X1 U49948 ( .A(n47848), .B(n47847), .Y(n47850) );
  NAND2X1 U49949 ( .A(writeback_exec_value_w[2]), .B(n38805), .Y(n47849) );
  NAND2X1 U49950 ( .A(n47850), .B(n47849), .Y(n47858) );
  NOR2X1 U49951 ( .A(n42909), .B(n37308), .Y(n47852) );
  NOR2X1 U49952 ( .A(n38932), .B(n37312), .Y(n47851) );
  NOR2X1 U49953 ( .A(n47852), .B(n47851), .Y(n47856) );
  NOR2X1 U49954 ( .A(n49637), .B(n37310), .Y(n47854) );
  NOR2X1 U49955 ( .A(n42917), .B(n37313), .Y(n47853) );
  NOR2X1 U49956 ( .A(n47854), .B(n47853), .Y(n47855) );
  NAND2X1 U49957 ( .A(n47856), .B(n47855), .Y(n47857) );
  NOR2X1 U49958 ( .A(n47858), .B(n47857), .Y(n47859) );
  NAND2X1 U49959 ( .A(n47860), .B(n47859), .Y(n72823) );
  NOR2X1 U49960 ( .A(n49625), .B(n48180), .Y(n47862) );
  NOR2X1 U49961 ( .A(n40041), .B(n48211), .Y(n47861) );
  NOR2X1 U49962 ( .A(n47862), .B(n47861), .Y(n47864) );
  NAND2X1 U49963 ( .A(n1977), .B(n49647), .Y(n47863) );
  NAND2X1 U49964 ( .A(n47864), .B(n47863), .Y(n47912) );
  NAND2X1 U49965 ( .A(n1992), .B(n40424), .Y(n47866) );
  NAND2X1 U49966 ( .A(n1990), .B(n57615), .Y(n47865) );
  NAND2X1 U49967 ( .A(n47866), .B(n47865), .Y(n47872) );
  NOR2X1 U49968 ( .A(n42628), .B(n36814), .Y(n47868) );
  NOR2X1 U49969 ( .A(n42684), .B(n37198), .Y(n47867) );
  NOR2X1 U49970 ( .A(n47868), .B(n47867), .Y(n47870) );
  NAND2X1 U49971 ( .A(n1994), .B(n40536), .Y(n47869) );
  NAND2X1 U49972 ( .A(n47870), .B(n47869), .Y(n47871) );
  NOR2X1 U49973 ( .A(n47872), .B(n47871), .Y(n47882) );
  NAND2X1 U49974 ( .A(n1984), .B(n42778), .Y(n47874) );
  NAND2X1 U49975 ( .A(n1982), .B(n73368), .Y(n47873) );
  NAND2X1 U49976 ( .A(n47874), .B(n47873), .Y(n47880) );
  NOR2X1 U49977 ( .A(n42896), .B(n36862), .Y(n47876) );
  NOR2X1 U49978 ( .A(n49599), .B(n36810), .Y(n47875) );
  NOR2X1 U49979 ( .A(n47876), .B(n47875), .Y(n47878) );
  NAND2X1 U49980 ( .A(n1985), .B(n39319), .Y(n47877) );
  NAND2X1 U49981 ( .A(n47878), .B(n47877), .Y(n47879) );
  NOR2X1 U49982 ( .A(n47880), .B(n47879), .Y(n47881) );
  NAND2X1 U49983 ( .A(n47882), .B(n47881), .Y(n47903) );
  NAND2X1 U49984 ( .A(n1978), .B(n38844), .Y(n47884) );
  NAND2X1 U49985 ( .A(n1976), .B(n42819), .Y(n47883) );
  NAND2X1 U49986 ( .A(n47884), .B(n47883), .Y(n47890) );
  NOR2X1 U49987 ( .A(n36609), .B(n37196), .Y(n47886) );
  NOR2X1 U49988 ( .A(n39654), .B(n36815), .Y(n47885) );
  NOR2X1 U49989 ( .A(n47886), .B(n47885), .Y(n47888) );
  NAND2X1 U49990 ( .A(n1980), .B(n40249), .Y(n47887) );
  NAND2X1 U49991 ( .A(n47888), .B(n47887), .Y(n47889) );
  NOR2X1 U49992 ( .A(n47890), .B(n47889), .Y(n47901) );
  NAND2X1 U49993 ( .A(n2000), .B(n57617), .Y(n47892) );
  NAND2X1 U49994 ( .A(n1998), .B(n38085), .Y(n47891) );
  NAND2X1 U49995 ( .A(n47892), .B(n47891), .Y(n47899) );
  NOR2X1 U49996 ( .A(n42903), .B(n37201), .Y(n47894) );
  NOR2X1 U49997 ( .A(n42623), .B(n37211), .Y(n47893) );
  NOR2X1 U49998 ( .A(n47894), .B(n47893), .Y(n47897) );
  NAND2X1 U49999 ( .A(n2001), .B(n47895), .Y(n47896) );
  NAND2X1 U50000 ( .A(n47897), .B(n47896), .Y(n47898) );
  NOR2X1 U50001 ( .A(n47899), .B(n47898), .Y(n47900) );
  NAND2X1 U50002 ( .A(n47901), .B(n47900), .Y(n47902) );
  NOR2X1 U50003 ( .A(n47903), .B(n47902), .Y(n47904) );
  NOR2X1 U50004 ( .A(n47904), .B(n42888), .Y(n47906) );
  NOR2X1 U50005 ( .A(n42914), .B(n37296), .Y(n47905) );
  NOR2X1 U50006 ( .A(n47906), .B(n47905), .Y(n47910) );
  NOR2X1 U50007 ( .A(n39335), .B(n37295), .Y(n47908) );
  NOR2X1 U50008 ( .A(n39572), .B(n37297), .Y(n47907) );
  NOR2X1 U50009 ( .A(n47908), .B(n47907), .Y(n47909) );
  NAND2X1 U50010 ( .A(n47910), .B(n47909), .Y(n47911) );
  NOR2X1 U50011 ( .A(n42900), .B(n37294), .Y(n47916) );
  NOR2X1 U50012 ( .A(n32011), .B(n32010), .Y(n47914) );
  NOR2X1 U50013 ( .A(n32008), .B(n32007), .Y(n47913) );
  NAND2X1 U50014 ( .A(n47914), .B(n47913), .Y(n62903) );
  NOR2X1 U50015 ( .A(n43080), .B(n42898), .Y(n47915) );
  NOR2X1 U50016 ( .A(n47916), .B(n47915), .Y(n47918) );
  NAND2X1 U50017 ( .A(writeback_exec_value_w[1]), .B(n38805), .Y(n47917) );
  NAND2X1 U50018 ( .A(n47918), .B(n47917), .Y(n47926) );
  NOR2X1 U50019 ( .A(n42910), .B(n48161), .Y(n47920) );
  NOR2X1 U50020 ( .A(n42913), .B(n36860), .Y(n47919) );
  NOR2X1 U50021 ( .A(n47920), .B(n47919), .Y(n47924) );
  NOR2X1 U50022 ( .A(n42911), .B(n36802), .Y(n47922) );
  NOR2X1 U50023 ( .A(n42918), .B(n36820), .Y(n47921) );
  NOR2X1 U50024 ( .A(n47922), .B(n47921), .Y(n47923) );
  NAND2X1 U50025 ( .A(n47924), .B(n47923), .Y(n47925) );
  NOR2X1 U50026 ( .A(n48105), .B(n48104), .Y(n47927) );
  NAND2X1 U50027 ( .A(n47927), .B(writeback_exec_value_w[0]), .Y(n62902) );
  NAND2X1 U50028 ( .A(n38793), .B(n62907), .Y(n61182) );
  INVX1 U50029 ( .A(n61182), .Y(n48107) );
  NOR2X1 U50030 ( .A(n35309), .B(n35308), .Y(n47929) );
  NOR2X1 U50031 ( .A(n35304), .B(n35303), .Y(n47928) );
  NAND2X1 U50032 ( .A(n47929), .B(n47928), .Y(n62904) );
  NAND2X1 U50033 ( .A(n48107), .B(n62904), .Y(n47930) );
  NOR2X1 U50034 ( .A(n42793), .B(n42663), .Y(n47931) );
  NAND2X1 U50035 ( .A(n47931), .B(n1960), .Y(n47932) );
  NOR2X1 U50036 ( .A(n42871), .B(n47932), .Y(n47936) );
  NOR2X1 U50037 ( .A(n42792), .B(n42662), .Y(n47933) );
  NAND2X1 U50038 ( .A(n47933), .B(n1958), .Y(n47934) );
  NOR2X1 U50039 ( .A(n42880), .B(n47934), .Y(n47935) );
  NOR2X1 U50040 ( .A(n47936), .B(n47935), .Y(n47944) );
  NAND2X1 U50041 ( .A(n38115), .B(n42667), .Y(n47938) );
  NAND2X1 U50042 ( .A(n42724), .B(n42689), .Y(n47937) );
  NOR2X1 U50043 ( .A(n47938), .B(n47937), .Y(n47942) );
  NOR2X1 U50044 ( .A(n1959), .B(n42794), .Y(n47940) );
  NOR2X1 U50045 ( .A(n1945), .B(n42789), .Y(n47939) );
  NOR2X1 U50046 ( .A(n47940), .B(n47939), .Y(n47941) );
  NAND2X1 U50047 ( .A(n47942), .B(n47941), .Y(n47943) );
  NAND2X1 U50048 ( .A(n47944), .B(n47943), .Y(n47960) );
  NOR2X1 U50049 ( .A(n42795), .B(n42664), .Y(n47945) );
  NAND2X1 U50050 ( .A(n47945), .B(n1961), .Y(n47946) );
  NOR2X1 U50051 ( .A(n42745), .B(n47946), .Y(n47950) );
  NOR2X1 U50052 ( .A(n42794), .B(n42663), .Y(n47947) );
  NAND2X1 U50053 ( .A(n47947), .B(n1957), .Y(n47948) );
  NOR2X1 U50054 ( .A(n42853), .B(n47948), .Y(n47949) );
  NOR2X1 U50055 ( .A(n47950), .B(n47949), .Y(n47958) );
  NAND2X1 U50056 ( .A(n42685), .B(n42669), .Y(n47952) );
  NAND2X1 U50057 ( .A(n42723), .B(n42731), .Y(n47951) );
  NOR2X1 U50058 ( .A(n47952), .B(n47951), .Y(n47956) );
  NOR2X1 U50059 ( .A(n1948), .B(n42790), .Y(n47954) );
  NOR2X1 U50060 ( .A(n1962), .B(n42795), .Y(n47953) );
  NOR2X1 U50061 ( .A(n47954), .B(n47953), .Y(n47955) );
  NAND2X1 U50062 ( .A(n47956), .B(n47955), .Y(n47957) );
  NAND2X1 U50063 ( .A(n47958), .B(n47957), .Y(n47959) );
  NAND2X1 U50064 ( .A(n42790), .B(n42664), .Y(n48109) );
  INVX1 U50065 ( .A(n48109), .Y(n48015) );
  NAND2X1 U50066 ( .A(n1950), .B(n42751), .Y(n47961) );
  NOR2X1 U50067 ( .A(n38366), .B(n47961), .Y(n47964) );
  NAND2X1 U50068 ( .A(n1951), .B(n42751), .Y(n47962) );
  NOR2X1 U50069 ( .A(n39647), .B(n47962), .Y(n47963) );
  NOR2X1 U50070 ( .A(n47964), .B(n47963), .Y(n47968) );
  NAND2X1 U50071 ( .A(n42792), .B(n42665), .Y(n47965) );
  NOR2X1 U50072 ( .A(n36799), .B(n47965), .Y(n47966) );
  NAND2X1 U50073 ( .A(n47966), .B(n48205), .Y(n47967) );
  NAND2X1 U50074 ( .A(n47968), .B(n47967), .Y(n47984) );
  NOR2X1 U50075 ( .A(n42668), .B(n42790), .Y(n47969) );
  NAND2X1 U50076 ( .A(n47969), .B(n1968), .Y(n47970) );
  NOR2X1 U50077 ( .A(n42870), .B(n47970), .Y(n47976) );
  NOR2X1 U50078 ( .A(n48186), .B(n48171), .Y(n47971) );
  NAND2X1 U50079 ( .A(n47971), .B(n1954), .Y(n47974) );
  NAND2X1 U50080 ( .A(n47974), .B(n47973), .Y(n47975) );
  NOR2X1 U50081 ( .A(n47976), .B(n47975), .Y(n47982) );
  NAND2X1 U50082 ( .A(opcode_opcode_w[18]), .B(n42795), .Y(n48114) );
  INVX1 U50083 ( .A(n48114), .Y(n48176) );
  NAND2X1 U50084 ( .A(n48176), .B(n42744), .Y(n47977) );
  NOR2X1 U50085 ( .A(n36812), .B(n47977), .Y(n47980) );
  NAND2X1 U50086 ( .A(n1944), .B(n48176), .Y(n47978) );
  NOR2X1 U50087 ( .A(n42879), .B(n47978), .Y(n47979) );
  NOR2X1 U50088 ( .A(n47980), .B(n47979), .Y(n47981) );
  NAND2X1 U50089 ( .A(n47982), .B(n47981), .Y(n47983) );
  NOR2X1 U50090 ( .A(n42667), .B(n42787), .Y(n47985) );
  NAND2X1 U50091 ( .A(n47985), .B(n1969), .Y(n47986) );
  NOR2X1 U50092 ( .A(n42746), .B(n47986), .Y(n47990) );
  NOR2X1 U50093 ( .A(n42667), .B(n42787), .Y(n47987) );
  NAND2X1 U50094 ( .A(n47987), .B(n1970), .Y(n47988) );
  NOR2X1 U50095 ( .A(n48186), .B(n47988), .Y(n47989) );
  NOR2X1 U50096 ( .A(n47990), .B(n47989), .Y(n47996) );
  NAND2X1 U50097 ( .A(n1952), .B(n42856), .Y(n47991) );
  NOR2X1 U50098 ( .A(n42869), .B(n47991), .Y(n47994) );
  NAND2X1 U50099 ( .A(n1943), .B(n42751), .Y(n47992) );
  NOR2X1 U50100 ( .A(n42853), .B(n47992), .Y(n47993) );
  NOR2X1 U50101 ( .A(n47994), .B(n47993), .Y(n47995) );
  NAND2X1 U50102 ( .A(n47996), .B(n47995), .Y(n48002) );
  NOR2X1 U50103 ( .A(n48585), .B(n36482), .Y(n47997) );
  NAND2X1 U50104 ( .A(n47997), .B(n1946), .Y(n48000) );
  NOR2X1 U50105 ( .A(n48585), .B(n42854), .Y(n47998) );
  NAND2X1 U50106 ( .A(n47998), .B(n1791), .Y(n47999) );
  NAND2X1 U50107 ( .A(n48000), .B(n47999), .Y(n48001) );
  NOR2X1 U50108 ( .A(n48002), .B(n48001), .Y(n48035) );
  NOR2X1 U50109 ( .A(n42669), .B(n42786), .Y(n48003) );
  NAND2X1 U50110 ( .A(n48003), .B(n1965), .Y(n48004) );
  NOR2X1 U50111 ( .A(n42854), .B(n48004), .Y(n48007) );
  NAND2X1 U50112 ( .A(opcode_opcode_w[18]), .B(n42788), .Y(n48138) );
  INVX1 U50113 ( .A(n48138), .Y(n48208) );
  NAND2X1 U50114 ( .A(n1963), .B(n48208), .Y(n48005) );
  NOR2X1 U50115 ( .A(n42736), .B(n48005), .Y(n48006) );
  NOR2X1 U50116 ( .A(n48007), .B(n48006), .Y(n48014) );
  NOR2X1 U50117 ( .A(opcode_opcode_w[18]), .B(n42789), .Y(n48008) );
  NOR2X1 U50118 ( .A(n42788), .B(n42664), .Y(n48009) );
  NAND2X1 U50119 ( .A(n48009), .B(n1949), .Y(n48010) );
  NOR2X1 U50120 ( .A(n42736), .B(n48010), .Y(n48011) );
  NOR2X1 U50121 ( .A(n48012), .B(n48011), .Y(n48013) );
  NAND2X1 U50122 ( .A(n48014), .B(n48013), .Y(n48033) );
  NAND2X1 U50123 ( .A(n1955), .B(n42751), .Y(n48016) );
  NOR2X1 U50124 ( .A(n42733), .B(n48016), .Y(n48024) );
  NAND2X1 U50125 ( .A(n42795), .B(n48094), .Y(n48018) );
  NAND2X1 U50126 ( .A(n42788), .B(n48089), .Y(n48017) );
  NAND2X1 U50127 ( .A(n48018), .B(n48017), .Y(n48022) );
  NOR2X1 U50128 ( .A(n42729), .B(n42723), .Y(n48020) );
  NOR2X1 U50129 ( .A(n42687), .B(n42665), .Y(n48019) );
  NAND2X1 U50130 ( .A(n48020), .B(n48019), .Y(n48021) );
  NOR2X1 U50131 ( .A(n48022), .B(n48021), .Y(n48023) );
  NOR2X1 U50132 ( .A(n48024), .B(n48023), .Y(n48031) );
  NOR2X1 U50133 ( .A(n42668), .B(n42790), .Y(n48025) );
  NAND2X1 U50134 ( .A(n48025), .B(n1967), .Y(n48026) );
  NOR2X1 U50135 ( .A(n39647), .B(n48026), .Y(n48029) );
  NAND2X1 U50136 ( .A(n42792), .B(n42663), .Y(n48184) );
  NOR2X1 U50137 ( .A(n48560), .B(n48027), .Y(n48028) );
  NOR2X1 U50138 ( .A(n48029), .B(n48028), .Y(n48030) );
  NAND2X1 U50139 ( .A(n48031), .B(n48030), .Y(n48032) );
  NOR2X1 U50140 ( .A(n48033), .B(n48032), .Y(n48034) );
  NAND2X1 U50141 ( .A(n48035), .B(n48034), .Y(n61177) );
  NOR2X1 U50142 ( .A(n42907), .B(n37298), .Y(n48037) );
  NOR2X1 U50143 ( .A(n40042), .B(n37299), .Y(n48036) );
  NOR2X1 U50144 ( .A(n48037), .B(n48036), .Y(n48039) );
  NAND2X1 U50145 ( .A(n1945), .B(n42707), .Y(n48038) );
  NAND2X1 U50146 ( .A(n48039), .B(n48038), .Y(n48088) );
  NAND2X1 U50147 ( .A(n1947), .B(n40520), .Y(n48041) );
  NAND2X1 U50148 ( .A(n1961), .B(n42627), .Y(n48040) );
  NAND2X1 U50149 ( .A(n48041), .B(n48040), .Y(n48047) );
  NOR2X1 U50150 ( .A(n42902), .B(n37217), .Y(n48043) );
  NOR2X1 U50151 ( .A(n42906), .B(n37220), .Y(n48042) );
  NOR2X1 U50152 ( .A(n48043), .B(n48042), .Y(n48045) );
  NAND2X1 U50153 ( .A(n1971), .B(n42620), .Y(n48044) );
  NAND2X1 U50154 ( .A(n48045), .B(n48044), .Y(n48046) );
  NOR2X1 U50155 ( .A(n48047), .B(n48046), .Y(n48058) );
  NAND2X1 U50156 ( .A(n1960), .B(n40426), .Y(n48049) );
  NAND2X1 U50157 ( .A(n1962), .B(n49685), .Y(n48048) );
  NAND2X1 U50158 ( .A(n48049), .B(n48048), .Y(n48056) );
  NOR2X1 U50159 ( .A(n42864), .B(n37218), .Y(n48052) );
  INVX1 U50160 ( .A(n1969), .Y(n48050) );
  NOR2X1 U50161 ( .A(n38213), .B(n48050), .Y(n48051) );
  NOR2X1 U50162 ( .A(n48052), .B(n48051), .Y(n48054) );
  NAND2X1 U50163 ( .A(n1963), .B(n42679), .Y(n48053) );
  NAND2X1 U50164 ( .A(n48054), .B(n48053), .Y(n48055) );
  NOR2X1 U50165 ( .A(n48056), .B(n48055), .Y(n48057) );
  NAND2X1 U50166 ( .A(n48058), .B(n48057), .Y(n48078) );
  NAND2X1 U50167 ( .A(n1952), .B(n42777), .Y(n48060) );
  NAND2X1 U50168 ( .A(n1944), .B(n38709), .Y(n48059) );
  NAND2X1 U50169 ( .A(n48060), .B(n48059), .Y(n48066) );
  NOR2X1 U50170 ( .A(n36609), .B(n37219), .Y(n48062) );
  NOR2X1 U50171 ( .A(n42896), .B(n37222), .Y(n48061) );
  NOR2X1 U50172 ( .A(n48062), .B(n48061), .Y(n48064) );
  NAND2X1 U50173 ( .A(n1950), .B(n73368), .Y(n48063) );
  NAND2X1 U50174 ( .A(n48064), .B(n48063), .Y(n48065) );
  NOR2X1 U50175 ( .A(n48066), .B(n48065), .Y(n48076) );
  NAND2X1 U50176 ( .A(n1958), .B(n46177), .Y(n48068) );
  NAND2X1 U50177 ( .A(n1953), .B(n39319), .Y(n48067) );
  NAND2X1 U50178 ( .A(n48068), .B(n48067), .Y(n48074) );
  NOR2X1 U50179 ( .A(n40857), .B(n36799), .Y(n48070) );
  NOR2X1 U50180 ( .A(n42893), .B(n37226), .Y(n48069) );
  NOR2X1 U50181 ( .A(n48070), .B(n48069), .Y(n48072) );
  NAND2X1 U50182 ( .A(n1954), .B(n40515), .Y(n48071) );
  NAND2X1 U50183 ( .A(n48072), .B(n48071), .Y(n48073) );
  NOR2X1 U50184 ( .A(n48074), .B(n48073), .Y(n48075) );
  NAND2X1 U50185 ( .A(n48076), .B(n48075), .Y(n48077) );
  NOR2X1 U50186 ( .A(n48078), .B(n48077), .Y(n48079) );
  NOR2X1 U50187 ( .A(n48079), .B(n42889), .Y(n48081) );
  NOR2X1 U50188 ( .A(n42916), .B(n37301), .Y(n48080) );
  NOR2X1 U50189 ( .A(n48081), .B(n48080), .Y(n48086) );
  INVX1 U50190 ( .A(n1964), .Y(n48082) );
  NOR2X1 U50191 ( .A(n39335), .B(n48082), .Y(n48084) );
  NOR2X1 U50192 ( .A(n39572), .B(n37302), .Y(n48083) );
  NOR2X1 U50193 ( .A(n48084), .B(n48083), .Y(n48085) );
  NAND2X1 U50194 ( .A(n48086), .B(n48085), .Y(n48087) );
  NOR2X1 U50195 ( .A(n39353), .B(n48089), .Y(n48091) );
  NOR2X1 U50196 ( .A(n43451), .B(n42899), .Y(n48090) );
  NOR2X1 U50197 ( .A(n48091), .B(n48090), .Y(n48093) );
  NAND2X1 U50198 ( .A(writeback_exec_value_w[0]), .B(n37976), .Y(n48092) );
  NAND2X1 U50199 ( .A(n48093), .B(n48092), .Y(n48102) );
  NOR2X1 U50200 ( .A(n49710), .B(n37300), .Y(n48096) );
  NOR2X1 U50201 ( .A(n42913), .B(n48094), .Y(n48095) );
  NOR2X1 U50202 ( .A(n48096), .B(n48095), .Y(n48100) );
  NOR2X1 U50203 ( .A(n40855), .B(n37303), .Y(n48098) );
  NOR2X1 U50204 ( .A(n42919), .B(n37304), .Y(n48097) );
  NOR2X1 U50205 ( .A(n48098), .B(n48097), .Y(n48099) );
  NAND2X1 U50206 ( .A(n48100), .B(n48099), .Y(n48101) );
  NAND2X1 U50207 ( .A(n36719), .B(n43732), .Y(n48103) );
  NAND2X1 U50208 ( .A(n43755), .B(n48103), .Y(n48226) );
  INVX1 U50209 ( .A(n48103), .Y(n57670) );
  NAND2X1 U50210 ( .A(n57670), .B(n43752), .Y(n48224) );
  NOR2X1 U50211 ( .A(n48105), .B(n48104), .Y(n48106) );
  NAND2X1 U50212 ( .A(n48106), .B(writeback_exec_value_w[1]), .Y(n62909) );
  NAND2X1 U50213 ( .A(n48107), .B(n62903), .Y(n48108) );
  NAND2X1 U50214 ( .A(n62909), .B(n48108), .Y(n62455) );
  NOR2X1 U50215 ( .A(n48109), .B(n36801), .Y(n48110) );
  NAND2X1 U50216 ( .A(n48110), .B(n42743), .Y(n48113) );
  NOR2X1 U50217 ( .A(n42855), .B(n48116), .Y(n48111) );
  NAND2X1 U50218 ( .A(n48111), .B(n1997), .Y(n48112) );
  NAND2X1 U50219 ( .A(n48113), .B(n48112), .Y(n48120) );
  NOR2X1 U50220 ( .A(n48114), .B(n36802), .Y(n48115) );
  INVX1 U50221 ( .A(n1998), .Y(n48117) );
  NOR2X1 U50222 ( .A(n48117), .B(n47965), .Y(n48118) );
  NOR2X1 U50223 ( .A(n48120), .B(n48119), .Y(n48145) );
  NOR2X1 U50224 ( .A(n42668), .B(n42786), .Y(n48121) );
  NAND2X1 U50225 ( .A(n48121), .B(n2000), .Y(n48122) );
  NOR2X1 U50226 ( .A(n48122), .B(n42871), .Y(n48125) );
  NAND2X1 U50227 ( .A(n1981), .B(n48176), .Y(n48123) );
  NOR2X1 U50228 ( .A(n42736), .B(n48123), .Y(n48124) );
  NOR2X1 U50229 ( .A(n48125), .B(n48124), .Y(n48130) );
  INVX1 U50230 ( .A(n2001), .Y(n48127) );
  NAND2X1 U50231 ( .A(n42793), .B(n42664), .Y(n48126) );
  NOR2X1 U50232 ( .A(n48127), .B(n48595), .Y(n48128) );
  NAND2X1 U50233 ( .A(n48128), .B(n42742), .Y(n48129) );
  NAND2X1 U50234 ( .A(n48130), .B(n48129), .Y(n48143) );
  NOR2X1 U50235 ( .A(n42668), .B(n42788), .Y(n48131) );
  NAND2X1 U50236 ( .A(n48131), .B(n2003), .Y(n48132) );
  NOR2X1 U50237 ( .A(n42736), .B(n48132), .Y(n48135) );
  NAND2X1 U50238 ( .A(n1995), .B(n48208), .Y(n48133) );
  NOR2X1 U50239 ( .A(n42738), .B(n48133), .Y(n48134) );
  NOR2X1 U50240 ( .A(n48135), .B(n48134), .Y(n48141) );
  NOR2X1 U50241 ( .A(n42686), .B(n42728), .Y(n48136) );
  NAND2X1 U50242 ( .A(n48136), .B(n42725), .Y(n48137) );
  NOR2X1 U50243 ( .A(n39883), .B(n48137), .Y(n48139) );
  NAND2X1 U50244 ( .A(n48139), .B(n1988), .Y(n48140) );
  NAND2X1 U50245 ( .A(n48141), .B(n48140), .Y(n48142) );
  NOR2X1 U50246 ( .A(n48143), .B(n48142), .Y(n48144) );
  NAND2X1 U50247 ( .A(n48145), .B(n48144), .Y(n62897) );
  NAND2X1 U50248 ( .A(n40449), .B(n40018), .Y(n48146) );
  NOR2X1 U50249 ( .A(n36860), .B(n48146), .Y(n48152) );
  NOR2X1 U50250 ( .A(n39882), .B(n42855), .Y(n48147) );
  NAND2X1 U50251 ( .A(n48147), .B(n1989), .Y(n48150) );
  NOR2X1 U50252 ( .A(n48560), .B(n48116), .Y(n48148) );
  NAND2X1 U50253 ( .A(n48148), .B(n1996), .Y(n48149) );
  NAND2X1 U50254 ( .A(n48150), .B(n48149), .Y(n48151) );
  NOR2X1 U50255 ( .A(n48152), .B(n48151), .Y(n48157) );
  NAND2X1 U50256 ( .A(n42734), .B(n48015), .Y(n48153) );
  NOR2X1 U50257 ( .A(n36862), .B(n48153), .Y(n48155) );
  NOR2X1 U50258 ( .A(n42854), .B(n38572), .Y(n48154) );
  NOR2X1 U50259 ( .A(n48155), .B(n48154), .Y(n48156) );
  NAND2X1 U50260 ( .A(n48157), .B(n48156), .Y(n62896) );
  NOR2X1 U50261 ( .A(n42786), .B(n42663), .Y(n48158) );
  NAND2X1 U50262 ( .A(n48158), .B(n1980), .Y(n48159) );
  NOR2X1 U50263 ( .A(n48186), .B(n48159), .Y(n48170) );
  NAND2X1 U50264 ( .A(n38115), .B(n42689), .Y(n48160) );
  NOR2X1 U50265 ( .A(n48161), .B(n48160), .Y(n48165) );
  NAND2X1 U50266 ( .A(n42687), .B(n42730), .Y(n48162) );
  NOR2X1 U50267 ( .A(n48163), .B(n48162), .Y(n48164) );
  NOR2X1 U50268 ( .A(n48165), .B(n48164), .Y(n48168) );
  NOR2X1 U50269 ( .A(n42663), .B(n42727), .Y(n48166) );
  NAND2X1 U50270 ( .A(n48166), .B(n42786), .Y(n48167) );
  NOR2X1 U50271 ( .A(n48168), .B(n48167), .Y(n48169) );
  NOR2X1 U50272 ( .A(n48170), .B(n48169), .Y(n48173) );
  NAND2X1 U50273 ( .A(n42786), .B(n42662), .Y(n48171) );
  NAND2X1 U50274 ( .A(n48173), .B(n48172), .Y(n48193) );
  NOR2X1 U50275 ( .A(n42722), .B(n42731), .Y(n48174) );
  NAND2X1 U50276 ( .A(n48208), .B(n42378), .Y(n48175) );
  NOR2X1 U50277 ( .A(n36814), .B(n48175), .Y(n48179) );
  NAND2X1 U50278 ( .A(n48176), .B(n42378), .Y(n48177) );
  NOR2X1 U50279 ( .A(n36815), .B(n48177), .Y(n48178) );
  NOR2X1 U50280 ( .A(n48179), .B(n48178), .Y(n48191) );
  NOR2X1 U50281 ( .A(n42727), .B(n48180), .Y(n48182) );
  NOR2X1 U50282 ( .A(opcode_opcode_w[17]), .B(n42730), .Y(n48181) );
  NAND2X1 U50283 ( .A(n48182), .B(n48181), .Y(n48183) );
  NOR2X1 U50284 ( .A(n48126), .B(n48183), .Y(n48189) );
  NOR2X1 U50285 ( .A(n42668), .B(n42790), .Y(n48185) );
  NAND2X1 U50286 ( .A(n48185), .B(n2002), .Y(n48187) );
  NOR2X1 U50287 ( .A(n48187), .B(n48186), .Y(n48188) );
  NOR2X1 U50288 ( .A(n48189), .B(n48188), .Y(n48190) );
  NAND2X1 U50289 ( .A(n48191), .B(n48190), .Y(n48192) );
  NOR2X1 U50290 ( .A(n42667), .B(n42794), .Y(n48194) );
  NAND2X1 U50291 ( .A(n48194), .B(n1984), .Y(n48197) );
  NOR2X1 U50292 ( .A(n42787), .B(n42663), .Y(n48195) );
  NAND2X1 U50293 ( .A(n48195), .B(n1978), .Y(n48196) );
  NAND2X1 U50294 ( .A(n48197), .B(n48196), .Y(n48198) );
  NAND2X1 U50295 ( .A(n48199), .B(n48198), .Y(n48207) );
  NOR2X1 U50296 ( .A(n42667), .B(n42795), .Y(n48200) );
  NAND2X1 U50297 ( .A(n48200), .B(n1982), .Y(n48203) );
  NOR2X1 U50298 ( .A(n42789), .B(n42663), .Y(n48201) );
  NAND2X1 U50299 ( .A(n48201), .B(n1976), .Y(n48202) );
  NAND2X1 U50300 ( .A(n48203), .B(n48202), .Y(n48204) );
  NAND2X1 U50301 ( .A(n48205), .B(n48204), .Y(n48206) );
  NAND2X1 U50302 ( .A(n48207), .B(n48206), .Y(n48223) );
  NAND2X1 U50303 ( .A(n1990), .B(n48208), .Y(n48209) );
  NOR2X1 U50304 ( .A(n42880), .B(n48209), .Y(n48218) );
  NAND2X1 U50305 ( .A(n42789), .B(n42665), .Y(n48210) );
  NOR2X1 U50306 ( .A(n48211), .B(n48210), .Y(n48215) );
  NAND2X1 U50307 ( .A(n42668), .B(n42793), .Y(n48212) );
  NOR2X1 U50308 ( .A(n48213), .B(n48212), .Y(n48214) );
  NOR2X1 U50309 ( .A(n48215), .B(n48214), .Y(n48216) );
  NOR2X1 U50310 ( .A(n48216), .B(n39647), .Y(n48217) );
  NOR2X1 U50311 ( .A(n48218), .B(n48217), .Y(n48221) );
  NOR2X1 U50312 ( .A(n39882), .B(n42869), .Y(n48219) );
  NAND2X1 U50313 ( .A(n48219), .B(n1992), .Y(n48220) );
  NAND2X1 U50314 ( .A(n48221), .B(n48220), .Y(n48222) );
  NAND2X1 U50315 ( .A(n48224), .B(n42719), .Y(n48225) );
  NAND2X1 U50316 ( .A(n43818), .B(n43457), .Y(n57632) );
  NOR2X1 U50317 ( .A(n42192), .B(n42046), .Y(n48227) );
  NAND2X1 U50318 ( .A(n43474), .B(n43804), .Y(n57790) );
  NAND2X1 U50319 ( .A(n48227), .B(n57790), .Y(n48228) );
  NAND2X1 U50320 ( .A(n57793), .B(n48228), .Y(n48690) );
  INVX1 U50321 ( .A(n48690), .Y(n48531) );
  NAND2X1 U50322 ( .A(writeback_exec_value_w[5]), .B(n43025), .Y(n48232) );
  NAND2X1 U50323 ( .A(n33679), .B(n33680), .Y(n48230) );
  NAND2X1 U50324 ( .A(n33676), .B(n33677), .Y(n48229) );
  OR2X1 U50325 ( .A(n48230), .B(n48229), .Y(n48516) );
  NAND2X1 U50326 ( .A(n38271), .B(n48516), .Y(n48231) );
  NAND2X1 U50327 ( .A(n48232), .B(n48231), .Y(n63834) );
  INVX1 U50328 ( .A(n63834), .Y(n63835) );
  NOR2X1 U50329 ( .A(n48184), .B(n42862), .Y(n48233) );
  NAND2X1 U50330 ( .A(n48233), .B(n2128), .Y(n48236) );
  NOR2X1 U50331 ( .A(n42670), .B(n42870), .Y(n48234) );
  NAND2X1 U50332 ( .A(n48234), .B(n2104), .Y(n48235) );
  NAND2X1 U50333 ( .A(n48236), .B(n48235), .Y(n48242) );
  NOR2X1 U50334 ( .A(n42753), .B(n42869), .Y(n48237) );
  NAND2X1 U50335 ( .A(n48237), .B(n2110), .Y(n48240) );
  NOR2X1 U50336 ( .A(n42674), .B(n42870), .Y(n48238) );
  NAND2X1 U50337 ( .A(n48238), .B(n2118), .Y(n48239) );
  NAND2X1 U50338 ( .A(n48240), .B(n48239), .Y(n48241) );
  NOR2X1 U50339 ( .A(n48242), .B(n48241), .Y(n48254) );
  NOR2X1 U50340 ( .A(n42670), .B(n42854), .Y(n48243) );
  NAND2X1 U50341 ( .A(n48243), .B(n1806), .Y(n48246) );
  NOR2X1 U50342 ( .A(n43016), .B(n42862), .Y(n48244) );
  NAND2X1 U50343 ( .A(n48244), .B(n2106), .Y(n48245) );
  NAND2X1 U50344 ( .A(n48246), .B(n48245), .Y(n48252) );
  NOR2X1 U50345 ( .A(n42672), .B(n42861), .Y(n48247) );
  NAND2X1 U50346 ( .A(n48247), .B(n2120), .Y(n48250) );
  NOR2X1 U50347 ( .A(n42753), .B(n42861), .Y(n48248) );
  NAND2X1 U50348 ( .A(n48248), .B(n2112), .Y(n48249) );
  NAND2X1 U50349 ( .A(n48250), .B(n48249), .Y(n48251) );
  NOR2X1 U50350 ( .A(n48252), .B(n48251), .Y(n48253) );
  NAND2X1 U50351 ( .A(n48254), .B(n48253), .Y(n48275) );
  NOR2X1 U50352 ( .A(n42674), .B(n42880), .Y(n48255) );
  NAND2X1 U50353 ( .A(n48255), .B(n2116), .Y(n48257) );
  NAND2X1 U50354 ( .A(n2114), .B(n43038), .Y(n48256) );
  NAND2X1 U50355 ( .A(n48257), .B(n48256), .Y(n48261) );
  NAND2X1 U50356 ( .A(n1807), .B(n39803), .Y(n48259) );
  NAND2X1 U50357 ( .A(n2122), .B(n43043), .Y(n48258) );
  NAND2X1 U50358 ( .A(n48259), .B(n48258), .Y(n48260) );
  NOR2X1 U50359 ( .A(n48261), .B(n48260), .Y(n48273) );
  NOR2X1 U50360 ( .A(n48184), .B(n36482), .Y(n48262) );
  NAND2X1 U50361 ( .A(n48262), .B(n2126), .Y(n48265) );
  NOR2X1 U50362 ( .A(n43016), .B(n38366), .Y(n48263) );
  NAND2X1 U50363 ( .A(n48263), .B(n2101), .Y(n48264) );
  NAND2X1 U50364 ( .A(n48265), .B(n48264), .Y(n48271) );
  NOR2X1 U50365 ( .A(n42752), .B(n42879), .Y(n48266) );
  NAND2X1 U50366 ( .A(n48266), .B(n2108), .Y(n48269) );
  NOR2X1 U50367 ( .A(n48184), .B(n42880), .Y(n48267) );
  NAND2X1 U50368 ( .A(n48267), .B(n2124), .Y(n48268) );
  NAND2X1 U50369 ( .A(n48269), .B(n48268), .Y(n48270) );
  NOR2X1 U50370 ( .A(n48271), .B(n48270), .Y(n48272) );
  NAND2X1 U50371 ( .A(n48273), .B(n48272), .Y(n48274) );
  NOR2X1 U50372 ( .A(n48275), .B(n48274), .Y(n48309) );
  NAND2X1 U50373 ( .A(n2121), .B(n43045), .Y(n48277) );
  NAND2X1 U50374 ( .A(n2127), .B(n43048), .Y(n48276) );
  NAND2X1 U50375 ( .A(n48277), .B(n48276), .Y(n48282) );
  NAND2X1 U50376 ( .A(n2119), .B(n49841), .Y(n48280) );
  NOR2X1 U50377 ( .A(n42670), .B(n42745), .Y(n48278) );
  NAND2X1 U50378 ( .A(n48278), .B(n2105), .Y(n48279) );
  NAND2X1 U50379 ( .A(n48280), .B(n48279), .Y(n48281) );
  NOR2X1 U50380 ( .A(n48282), .B(n48281), .Y(n48288) );
  NOR2X1 U50381 ( .A(n57625), .B(n37112), .Y(n48286) );
  NAND2X1 U50382 ( .A(n2113), .B(n38764), .Y(n48284) );
  NAND2X1 U50383 ( .A(n2129), .B(n43056), .Y(n48283) );
  NAND2X1 U50384 ( .A(n48284), .B(n48283), .Y(n48285) );
  NOR2X1 U50385 ( .A(n48286), .B(n48285), .Y(n48287) );
  NAND2X1 U50386 ( .A(n48288), .B(n48287), .Y(n48307) );
  NAND2X1 U50387 ( .A(n2125), .B(n43061), .Y(n48290) );
  NAND2X1 U50388 ( .A(n2123), .B(n39132), .Y(n48289) );
  NAND2X1 U50389 ( .A(n48290), .B(n48289), .Y(n48294) );
  NAND2X1 U50390 ( .A(n2115), .B(n43064), .Y(n48292) );
  NAND2X1 U50391 ( .A(n2102), .B(n43066), .Y(n48291) );
  NAND2X1 U50392 ( .A(n48292), .B(n48291), .Y(n48293) );
  NOR2X1 U50393 ( .A(n48294), .B(n48293), .Y(n48305) );
  NOR2X1 U50394 ( .A(n42753), .B(n39647), .Y(n48295) );
  NAND2X1 U50395 ( .A(n48295), .B(n2109), .Y(n48298) );
  NOR2X1 U50396 ( .A(n43016), .B(n39647), .Y(n48296) );
  NAND2X1 U50397 ( .A(n48296), .B(n2103), .Y(n48297) );
  NAND2X1 U50398 ( .A(n48298), .B(n48297), .Y(n48303) );
  NAND2X1 U50399 ( .A(n2117), .B(n40154), .Y(n48301) );
  NOR2X1 U50400 ( .A(n42752), .B(n42746), .Y(n48299) );
  NAND2X1 U50401 ( .A(n48299), .B(n2111), .Y(n48300) );
  NAND2X1 U50402 ( .A(n48301), .B(n48300), .Y(n48302) );
  NOR2X1 U50403 ( .A(n48303), .B(n48302), .Y(n48304) );
  NAND2X1 U50404 ( .A(n48305), .B(n48304), .Y(n48306) );
  NOR2X1 U50405 ( .A(n48307), .B(n48306), .Y(n48308) );
  NAND2X1 U50406 ( .A(n48309), .B(n48308), .Y(n63833) );
  NAND2X1 U50407 ( .A(n42806), .B(n63833), .Y(n63550) );
  NOR2X1 U50408 ( .A(n33542), .B(n33541), .Y(n48311) );
  NOR2X1 U50409 ( .A(n33540), .B(n33539), .Y(n48310) );
  NAND2X1 U50410 ( .A(n48311), .B(n48310), .Y(n48452) );
  NOR2X1 U50411 ( .A(n48184), .B(n42861), .Y(n48312) );
  NAND2X1 U50412 ( .A(n48312), .B(n2096), .Y(n48315) );
  NOR2X1 U50413 ( .A(n42670), .B(n42870), .Y(n48313) );
  NAND2X1 U50414 ( .A(n48313), .B(n2072), .Y(n48314) );
  NAND2X1 U50415 ( .A(n48315), .B(n48314), .Y(n48321) );
  NOR2X1 U50416 ( .A(n42857), .B(n36482), .Y(n48316) );
  NAND2X1 U50417 ( .A(n2078), .B(n48316), .Y(n48319) );
  NOR2X1 U50418 ( .A(n48607), .B(n42869), .Y(n48317) );
  NAND2X1 U50419 ( .A(n2086), .B(n48317), .Y(n48318) );
  NAND2X1 U50420 ( .A(n48319), .B(n48318), .Y(n48320) );
  NOR2X1 U50421 ( .A(n48321), .B(n48320), .Y(n48333) );
  NOR2X1 U50422 ( .A(n43015), .B(n42855), .Y(n48322) );
  NAND2X1 U50423 ( .A(n48322), .B(n1815), .Y(n48325) );
  NOR2X1 U50424 ( .A(n42670), .B(n42862), .Y(n48323) );
  NAND2X1 U50425 ( .A(n48323), .B(n2074), .Y(n48324) );
  NAND2X1 U50426 ( .A(n48325), .B(n48324), .Y(n48331) );
  NOR2X1 U50427 ( .A(n39883), .B(n42861), .Y(n48326) );
  NAND2X1 U50428 ( .A(n2088), .B(n48326), .Y(n48329) );
  NOR2X1 U50429 ( .A(n42755), .B(n42862), .Y(n48327) );
  NAND2X1 U50430 ( .A(n2080), .B(n48327), .Y(n48328) );
  NAND2X1 U50431 ( .A(n48329), .B(n48328), .Y(n48330) );
  NOR2X1 U50432 ( .A(n48331), .B(n48330), .Y(n48332) );
  NAND2X1 U50433 ( .A(n48333), .B(n48332), .Y(n48356) );
  NOR2X1 U50434 ( .A(n48607), .B(n38366), .Y(n48334) );
  NAND2X1 U50435 ( .A(n2084), .B(n48334), .Y(n48337) );
  NOR2X1 U50436 ( .A(n48560), .B(n48607), .Y(n48335) );
  NAND2X1 U50437 ( .A(n48335), .B(n2082), .Y(n48336) );
  NAND2X1 U50438 ( .A(n48337), .B(n48336), .Y(n48342) );
  NOR2X1 U50439 ( .A(n48560), .B(n43015), .Y(n48338) );
  NAND2X1 U50440 ( .A(n48338), .B(n1816), .Y(n48340) );
  NAND2X1 U50441 ( .A(n48340), .B(n48339), .Y(n48341) );
  NOR2X1 U50442 ( .A(n48342), .B(n48341), .Y(n48354) );
  NOR2X1 U50443 ( .A(n48126), .B(n42870), .Y(n48343) );
  NAND2X1 U50444 ( .A(n48343), .B(n2094), .Y(n48346) );
  NOR2X1 U50445 ( .A(n42670), .B(n42879), .Y(n48344) );
  NAND2X1 U50446 ( .A(n2069), .B(n48344), .Y(n48345) );
  NAND2X1 U50447 ( .A(n48346), .B(n48345), .Y(n48352) );
  NOR2X1 U50448 ( .A(n42754), .B(n42880), .Y(n48347) );
  NAND2X1 U50449 ( .A(n2076), .B(n48347), .Y(n48350) );
  NOR2X1 U50450 ( .A(n48184), .B(n38366), .Y(n48348) );
  NAND2X1 U50451 ( .A(n48348), .B(n2092), .Y(n48349) );
  NAND2X1 U50452 ( .A(n48350), .B(n48349), .Y(n48351) );
  NOR2X1 U50453 ( .A(n48352), .B(n48351), .Y(n48353) );
  NAND2X1 U50454 ( .A(n48354), .B(n48353), .Y(n48355) );
  NOR2X1 U50455 ( .A(n48356), .B(n48355), .Y(n63200) );
  NAND2X1 U50456 ( .A(n40448), .B(n42756), .Y(n48357) );
  NOR2X1 U50457 ( .A(n36949), .B(n48357), .Y(n48358) );
  NOR2X1 U50458 ( .A(n48359), .B(n48358), .Y(n48365) );
  NAND2X1 U50459 ( .A(n40448), .B(n42673), .Y(n48360) );
  NOR2X1 U50460 ( .A(n36945), .B(n48360), .Y(n48363) );
  NAND2X1 U50461 ( .A(n42743), .B(n42758), .Y(n48361) );
  NOR2X1 U50462 ( .A(n36965), .B(n48361), .Y(n48362) );
  NOR2X1 U50463 ( .A(n48363), .B(n48362), .Y(n48364) );
  NAND2X1 U50464 ( .A(n48365), .B(n48364), .Y(n48379) );
  NAND2X1 U50465 ( .A(n42756), .B(n40076), .Y(n48366) );
  NOR2X1 U50466 ( .A(n36947), .B(n48366), .Y(n48369) );
  NAND2X1 U50467 ( .A(n40076), .B(n42673), .Y(n48367) );
  NOR2X1 U50468 ( .A(n36969), .B(n48367), .Y(n48368) );
  NOR2X1 U50469 ( .A(n48369), .B(n48368), .Y(n48377) );
  NAND2X1 U50470 ( .A(n48372), .B(n40076), .Y(n48371) );
  NOR2X1 U50471 ( .A(n36961), .B(n48371), .Y(n48375) );
  NAND2X1 U50472 ( .A(n39669), .B(n40448), .Y(n48373) );
  NOR2X1 U50473 ( .A(n36982), .B(n48373), .Y(n48374) );
  NOR2X1 U50474 ( .A(n48375), .B(n48374), .Y(n48376) );
  NAND2X1 U50475 ( .A(n48377), .B(n48376), .Y(n48378) );
  NOR2X1 U50476 ( .A(n48379), .B(n48378), .Y(n48398) );
  NAND2X1 U50477 ( .A(n42735), .B(n39669), .Y(n48380) );
  NOR2X1 U50478 ( .A(n36936), .B(n48380), .Y(n48383) );
  NAND2X1 U50479 ( .A(n42734), .B(n43018), .Y(n48381) );
  NOR2X1 U50480 ( .A(n36942), .B(n48381), .Y(n48382) );
  NOR2X1 U50481 ( .A(n48383), .B(n48382), .Y(n48385) );
  NAND2X1 U50482 ( .A(n2081), .B(n38764), .Y(n48384) );
  NAND2X1 U50483 ( .A(n48385), .B(n48384), .Y(n48396) );
  NAND2X1 U50484 ( .A(n42742), .B(n43017), .Y(n48386) );
  NOR2X1 U50485 ( .A(n36941), .B(n48386), .Y(n48388) );
  NOR2X1 U50486 ( .A(n48388), .B(n48387), .Y(n48394) );
  NAND2X1 U50487 ( .A(n42744), .B(n39584), .Y(n48389) );
  NOR2X1 U50488 ( .A(n36944), .B(n48389), .Y(n48392) );
  NAND2X1 U50489 ( .A(n42735), .B(n42673), .Y(n48390) );
  NOR2X1 U50490 ( .A(n36966), .B(n48390), .Y(n48391) );
  NOR2X1 U50491 ( .A(n48392), .B(n48391), .Y(n48393) );
  NAND2X1 U50492 ( .A(n48394), .B(n48393), .Y(n48395) );
  NOR2X1 U50493 ( .A(n48396), .B(n48395), .Y(n48397) );
  NAND2X1 U50494 ( .A(n42515), .B(n48399), .Y(n62923) );
  NAND2X1 U50495 ( .A(n39946), .B(n43469), .Y(n48530) );
  NOR2X1 U50496 ( .A(n42908), .B(n36982), .Y(n48401) );
  NOR2X1 U50497 ( .A(n40041), .B(n36949), .Y(n48400) );
  NOR2X1 U50498 ( .A(n48401), .B(n48400), .Y(n48403) );
  NAND2X1 U50499 ( .A(n2071), .B(n42707), .Y(n48402) );
  NAND2X1 U50500 ( .A(n48403), .B(n48402), .Y(n48451) );
  NAND2X1 U50501 ( .A(n2073), .B(n40519), .Y(n48405) );
  NAND2X1 U50502 ( .A(n2087), .B(n42625), .Y(n48404) );
  NAND2X1 U50503 ( .A(n48405), .B(n48404), .Y(n48411) );
  NOR2X1 U50504 ( .A(n42903), .B(n37138), .Y(n48407) );
  NOR2X1 U50505 ( .A(n42906), .B(n37143), .Y(n48406) );
  NOR2X1 U50506 ( .A(n48407), .B(n48406), .Y(n48409) );
  NAND2X1 U50507 ( .A(n2097), .B(n42617), .Y(n48408) );
  NAND2X1 U50508 ( .A(n48409), .B(n48408), .Y(n48410) );
  NOR2X1 U50509 ( .A(n48411), .B(n48410), .Y(n48421) );
  NAND2X1 U50510 ( .A(n2086), .B(n40426), .Y(n48413) );
  NAND2X1 U50511 ( .A(n2088), .B(n40536), .Y(n48412) );
  NAND2X1 U50512 ( .A(n48413), .B(n48412), .Y(n48419) );
  NOR2X1 U50513 ( .A(n42865), .B(n37141), .Y(n48415) );
  NOR2X1 U50514 ( .A(n42858), .B(n36944), .Y(n48414) );
  NOR2X1 U50515 ( .A(n48415), .B(n48414), .Y(n48417) );
  NAND2X1 U50516 ( .A(n2089), .B(n42681), .Y(n48416) );
  NAND2X1 U50517 ( .A(n48417), .B(n48416), .Y(n48418) );
  NOR2X1 U50518 ( .A(n48419), .B(n48418), .Y(n48420) );
  NAND2X1 U50519 ( .A(n48421), .B(n48420), .Y(n48441) );
  NAND2X1 U50520 ( .A(n2078), .B(n42778), .Y(n48423) );
  NAND2X1 U50521 ( .A(n2069), .B(n38710), .Y(n48422) );
  NAND2X1 U50522 ( .A(n48423), .B(n48422), .Y(n48429) );
  NOR2X1 U50523 ( .A(n42891), .B(n36942), .Y(n48425) );
  NOR2X1 U50524 ( .A(n42896), .B(n37145), .Y(n48424) );
  NOR2X1 U50525 ( .A(n48425), .B(n48424), .Y(n48427) );
  NAND2X1 U50526 ( .A(n2076), .B(n42675), .Y(n48426) );
  NAND2X1 U50527 ( .A(n48427), .B(n48426), .Y(n48428) );
  NOR2X1 U50528 ( .A(n48429), .B(n48428), .Y(n48439) );
  NAND2X1 U50529 ( .A(n2084), .B(n46177), .Y(n48431) );
  NAND2X1 U50530 ( .A(n2079), .B(n39318), .Y(n48430) );
  NAND2X1 U50531 ( .A(n48431), .B(n48430), .Y(n48437) );
  NOR2X1 U50532 ( .A(n40857), .B(n37146), .Y(n48433) );
  NOR2X1 U50533 ( .A(n40851), .B(n37149), .Y(n48432) );
  NOR2X1 U50534 ( .A(n48433), .B(n48432), .Y(n48435) );
  NAND2X1 U50535 ( .A(n2080), .B(n40514), .Y(n48434) );
  NAND2X1 U50536 ( .A(n48435), .B(n48434), .Y(n48436) );
  NOR2X1 U50537 ( .A(n48437), .B(n48436), .Y(n48438) );
  NAND2X1 U50538 ( .A(n48439), .B(n48438), .Y(n48440) );
  NOR2X1 U50539 ( .A(n48441), .B(n48440), .Y(n48442) );
  NOR2X1 U50540 ( .A(n48442), .B(n42890), .Y(n48444) );
  NOR2X1 U50541 ( .A(n42915), .B(n36969), .Y(n48443) );
  NOR2X1 U50542 ( .A(n48444), .B(n48443), .Y(n48449) );
  INVX1 U50543 ( .A(n2090), .Y(n48445) );
  NOR2X1 U50544 ( .A(n39335), .B(n48445), .Y(n48447) );
  NOR2X1 U50545 ( .A(n49624), .B(n36961), .Y(n48446) );
  NOR2X1 U50546 ( .A(n48447), .B(n48446), .Y(n48448) );
  NAND2X1 U50547 ( .A(n48449), .B(n48448), .Y(n48450) );
  NOR2X1 U50548 ( .A(n40407), .B(n37291), .Y(n48454) );
  NOR2X1 U50549 ( .A(n43261), .B(n42899), .Y(n48453) );
  NOR2X1 U50550 ( .A(n48454), .B(n48453), .Y(n48456) );
  NAND2X1 U50551 ( .A(writeback_exec_value_w[4]), .B(n37976), .Y(n48455) );
  NAND2X1 U50552 ( .A(n48456), .B(n48455), .Y(n48464) );
  NOR2X1 U50553 ( .A(n42909), .B(n36945), .Y(n48458) );
  NOR2X1 U50554 ( .A(n38932), .B(n37293), .Y(n48457) );
  NOR2X1 U50555 ( .A(n48458), .B(n48457), .Y(n48462) );
  NOR2X1 U50556 ( .A(n40855), .B(n37292), .Y(n48460) );
  NOR2X1 U50557 ( .A(n42917), .B(n36947), .Y(n48459) );
  NOR2X1 U50558 ( .A(n48460), .B(n48459), .Y(n48461) );
  NAND2X1 U50559 ( .A(n48462), .B(n48461), .Y(n48463) );
  NOR2X1 U50560 ( .A(n49625), .B(n37279), .Y(n48466) );
  NOR2X1 U50561 ( .A(n40042), .B(n37283), .Y(n48465) );
  NOR2X1 U50562 ( .A(n48466), .B(n48465), .Y(n48468) );
  NAND2X1 U50563 ( .A(n2103), .B(n42706), .Y(n48467) );
  NAND2X1 U50564 ( .A(n48468), .B(n48467), .Y(n48515) );
  NAND2X1 U50565 ( .A(n2105), .B(n40520), .Y(n48470) );
  NAND2X1 U50566 ( .A(n2119), .B(n42627), .Y(n48469) );
  NAND2X1 U50567 ( .A(n48470), .B(n48469), .Y(n48476) );
  NOR2X1 U50568 ( .A(n42902), .B(n37109), .Y(n48472) );
  NOR2X1 U50569 ( .A(n42905), .B(n37113), .Y(n48471) );
  NOR2X1 U50570 ( .A(n48472), .B(n48471), .Y(n48474) );
  NAND2X1 U50571 ( .A(n2129), .B(n42620), .Y(n48473) );
  NAND2X1 U50572 ( .A(n48474), .B(n48473), .Y(n48475) );
  NOR2X1 U50573 ( .A(n48476), .B(n48475), .Y(n48486) );
  NAND2X1 U50574 ( .A(n2118), .B(n40425), .Y(n48478) );
  NAND2X1 U50575 ( .A(n2120), .B(n40536), .Y(n48477) );
  NAND2X1 U50576 ( .A(n48478), .B(n48477), .Y(n48484) );
  NOR2X1 U50577 ( .A(n42647), .B(n37110), .Y(n48480) );
  NOR2X1 U50578 ( .A(n42858), .B(n37115), .Y(n48479) );
  NOR2X1 U50579 ( .A(n48480), .B(n48479), .Y(n48482) );
  NAND2X1 U50580 ( .A(n2121), .B(n42678), .Y(n48481) );
  NAND2X1 U50581 ( .A(n48482), .B(n48481), .Y(n48483) );
  NOR2X1 U50582 ( .A(n48484), .B(n48483), .Y(n48485) );
  NAND2X1 U50583 ( .A(n48486), .B(n48485), .Y(n48506) );
  NAND2X1 U50584 ( .A(n2110), .B(n42777), .Y(n48488) );
  NAND2X1 U50585 ( .A(n2101), .B(n38710), .Y(n48487) );
  NAND2X1 U50586 ( .A(n48488), .B(n48487), .Y(n48494) );
  NOR2X1 U50587 ( .A(n42892), .B(n37112), .Y(n48490) );
  NOR2X1 U50588 ( .A(n42896), .B(n37116), .Y(n48489) );
  NOR2X1 U50589 ( .A(n48490), .B(n48489), .Y(n48492) );
  NAND2X1 U50590 ( .A(n2108), .B(n46174), .Y(n48491) );
  NAND2X1 U50591 ( .A(n48492), .B(n48491), .Y(n48493) );
  NOR2X1 U50592 ( .A(n48494), .B(n48493), .Y(n48504) );
  NAND2X1 U50593 ( .A(n2116), .B(n57615), .Y(n48496) );
  NAND2X1 U50594 ( .A(n2111), .B(n40537), .Y(n48495) );
  NAND2X1 U50595 ( .A(n48496), .B(n48495), .Y(n48502) );
  NOR2X1 U50596 ( .A(n38627), .B(n42875), .Y(n48498) );
  NOR2X1 U50597 ( .A(n40497), .B(n37117), .Y(n48497) );
  NOR2X1 U50598 ( .A(n48498), .B(n48497), .Y(n48500) );
  NAND2X1 U50599 ( .A(n2112), .B(n40515), .Y(n48499) );
  NAND2X1 U50600 ( .A(n48500), .B(n48499), .Y(n48501) );
  NOR2X1 U50601 ( .A(n48502), .B(n48501), .Y(n48503) );
  NAND2X1 U50602 ( .A(n48504), .B(n48503), .Y(n48505) );
  NOR2X1 U50603 ( .A(n48506), .B(n48505), .Y(n48507) );
  NOR2X1 U50604 ( .A(n48507), .B(n42890), .Y(n48509) );
  NOR2X1 U50605 ( .A(n42915), .B(n37286), .Y(n48508) );
  NOR2X1 U50606 ( .A(n48509), .B(n48508), .Y(n48513) );
  NOR2X1 U50607 ( .A(n40277), .B(n37284), .Y(n48511) );
  NOR2X1 U50608 ( .A(n42901), .B(n37287), .Y(n48510) );
  NOR2X1 U50609 ( .A(n48511), .B(n48510), .Y(n48512) );
  NAND2X1 U50610 ( .A(n48513), .B(n48512), .Y(n48514) );
  NOR2X1 U50611 ( .A(n42900), .B(n37282), .Y(n48518) );
  NOR2X1 U50612 ( .A(n43114), .B(n42899), .Y(n48517) );
  NOR2X1 U50613 ( .A(n48518), .B(n48517), .Y(n48520) );
  NAND2X1 U50614 ( .A(writeback_exec_value_w[5]), .B(n37976), .Y(n48519) );
  NAND2X1 U50615 ( .A(n48520), .B(n48519), .Y(n48528) );
  NOR2X1 U50616 ( .A(n42910), .B(n37285), .Y(n48522) );
  NOR2X1 U50617 ( .A(n42913), .B(n37289), .Y(n48521) );
  NOR2X1 U50618 ( .A(n48522), .B(n48521), .Y(n48526) );
  NOR2X1 U50619 ( .A(n49637), .B(n37288), .Y(n48524) );
  NOR2X1 U50620 ( .A(n42918), .B(n37290), .Y(n48523) );
  NOR2X1 U50621 ( .A(n48524), .B(n48523), .Y(n48525) );
  NAND2X1 U50622 ( .A(n48526), .B(n48525), .Y(n48527) );
  NAND2X1 U50623 ( .A(n43763), .B(n38611), .Y(n48529) );
  NAND2X1 U50624 ( .A(n48530), .B(n48529), .Y(n57771) );
  NAND2X1 U50625 ( .A(n48531), .B(n57771), .Y(n48535) );
  NOR2X1 U50626 ( .A(n43769), .B(n39943), .Y(n48533) );
  NAND2X1 U50627 ( .A(n48690), .B(n43466), .Y(n48532) );
  NAND2X1 U50628 ( .A(n48533), .B(n48532), .Y(n48534) );
  NAND2X1 U50629 ( .A(n48535), .B(n48534), .Y(n48695) );
  NAND2X1 U50630 ( .A(writeback_exec_value_w[6]), .B(n43026), .Y(n48539) );
  NAND2X1 U50631 ( .A(n34760), .B(n34761), .Y(n48537) );
  NAND2X1 U50632 ( .A(n34758), .B(n34759), .Y(n48536) );
  OR2X1 U50633 ( .A(n48537), .B(n48536), .Y(n48676) );
  NAND2X1 U50634 ( .A(n38271), .B(n48676), .Y(n48538) );
  NAND2X1 U50635 ( .A(n48539), .B(n48538), .Y(n64081) );
  INVX1 U50636 ( .A(n64081), .Y(n64083) );
  NOR2X1 U50637 ( .A(n48184), .B(n42862), .Y(n48540) );
  NAND2X1 U50638 ( .A(n48540), .B(n2345), .Y(n48542) );
  NAND2X1 U50639 ( .A(n2321), .B(n38407), .Y(n48541) );
  NAND2X1 U50640 ( .A(n48542), .B(n48541), .Y(n48546) );
  NAND2X1 U50641 ( .A(n2327), .B(n43344), .Y(n48544) );
  NAND2X1 U50642 ( .A(n2335), .B(n43028), .Y(n48543) );
  NAND2X1 U50643 ( .A(n48544), .B(n48543), .Y(n48545) );
  NOR2X1 U50644 ( .A(n48546), .B(n48545), .Y(n48556) );
  NAND2X1 U50645 ( .A(n1833), .B(n43029), .Y(n48548) );
  NAND2X1 U50646 ( .A(n2323), .B(n43033), .Y(n48547) );
  NAND2X1 U50647 ( .A(n48548), .B(n48547), .Y(n48554) );
  NOR2X1 U50648 ( .A(n42674), .B(n42861), .Y(n48549) );
  NAND2X1 U50649 ( .A(n48549), .B(n2337), .Y(n48552) );
  NOR2X1 U50650 ( .A(n42752), .B(n42862), .Y(n48550) );
  NAND2X1 U50651 ( .A(n48550), .B(n2329), .Y(n48551) );
  NAND2X1 U50652 ( .A(n48552), .B(n48551), .Y(n48553) );
  NOR2X1 U50653 ( .A(n48554), .B(n48553), .Y(n48555) );
  NAND2X1 U50654 ( .A(n48556), .B(n48555), .Y(n48575) );
  NAND2X1 U50655 ( .A(n2333), .B(n41786), .Y(n48559) );
  NOR2X1 U50656 ( .A(n48560), .B(n42672), .Y(n48557) );
  NAND2X1 U50657 ( .A(n48557), .B(n2331), .Y(n48558) );
  NAND2X1 U50658 ( .A(n48559), .B(n48558), .Y(n48565) );
  NAND2X1 U50659 ( .A(n2347), .B(n39804), .Y(n48563) );
  NOR2X1 U50660 ( .A(n48560), .B(n48184), .Y(n48561) );
  NAND2X1 U50661 ( .A(n48561), .B(n2339), .Y(n48562) );
  NAND2X1 U50662 ( .A(n48563), .B(n48562), .Y(n48564) );
  NOR2X1 U50663 ( .A(n48565), .B(n48564), .Y(n48573) );
  NAND2X1 U50664 ( .A(n2343), .B(n43360), .Y(n48567) );
  NAND2X1 U50665 ( .A(n2318), .B(n43346), .Y(n48566) );
  NAND2X1 U50666 ( .A(n48567), .B(n48566), .Y(n48571) );
  NAND2X1 U50667 ( .A(n2325), .B(n43339), .Y(n48569) );
  NAND2X1 U50668 ( .A(n2341), .B(n43366), .Y(n48568) );
  NAND2X1 U50669 ( .A(n48569), .B(n48568), .Y(n48570) );
  NOR2X1 U50670 ( .A(n48571), .B(n48570), .Y(n48572) );
  NAND2X1 U50671 ( .A(n48573), .B(n48572), .Y(n48574) );
  NOR2X1 U50672 ( .A(n48575), .B(n48574), .Y(n48623) );
  NOR2X1 U50673 ( .A(n42674), .B(n42738), .Y(n48576) );
  NAND2X1 U50674 ( .A(n48576), .B(n2338), .Y(n48579) );
  NOR2X1 U50675 ( .A(n48184), .B(n42745), .Y(n48577) );
  NAND2X1 U50676 ( .A(n48577), .B(n2344), .Y(n48578) );
  NAND2X1 U50677 ( .A(n48579), .B(n48578), .Y(n48584) );
  NOR2X1 U50678 ( .A(n42672), .B(n42746), .Y(n48580) );
  NAND2X1 U50679 ( .A(n48580), .B(n2336), .Y(n48582) );
  NAND2X1 U50680 ( .A(n2322), .B(n43052), .Y(n48581) );
  NAND2X1 U50681 ( .A(n48582), .B(n48581), .Y(n48583) );
  NOR2X1 U50682 ( .A(n48584), .B(n48583), .Y(n48593) );
  NOR2X1 U50683 ( .A(n43370), .B(n37104), .Y(n48591) );
  NOR2X1 U50684 ( .A(n43016), .B(n42737), .Y(n48586) );
  NAND2X1 U50685 ( .A(n48586), .B(n2324), .Y(n48589) );
  NOR2X1 U50686 ( .A(n48184), .B(n42737), .Y(n48587) );
  NAND2X1 U50687 ( .A(n48587), .B(n2346), .Y(n48588) );
  NAND2X1 U50688 ( .A(n48589), .B(n48588), .Y(n48590) );
  NOR2X1 U50689 ( .A(n48591), .B(n48590), .Y(n48592) );
  NAND2X1 U50690 ( .A(n48593), .B(n48592), .Y(n48621) );
  NOR2X1 U50691 ( .A(n39647), .B(n48184), .Y(n48594) );
  NAND2X1 U50692 ( .A(n48594), .B(n2342), .Y(n48598) );
  NOR2X1 U50693 ( .A(n42854), .B(n48184), .Y(n48596) );
  NAND2X1 U50694 ( .A(n48596), .B(n2340), .Y(n48597) );
  NAND2X1 U50695 ( .A(n48598), .B(n48597), .Y(n48604) );
  NOR2X1 U50696 ( .A(n42672), .B(n42854), .Y(n48599) );
  NAND2X1 U50697 ( .A(n48599), .B(n2332), .Y(n48602) );
  NOR2X1 U50698 ( .A(n42855), .B(n42752), .Y(n48600) );
  NAND2X1 U50699 ( .A(n48600), .B(n2319), .Y(n48601) );
  NAND2X1 U50700 ( .A(n48602), .B(n48601), .Y(n48603) );
  NOR2X1 U50701 ( .A(n48604), .B(n48603), .Y(n48619) );
  NOR2X1 U50702 ( .A(n42753), .B(n42746), .Y(n48606) );
  NAND2X1 U50703 ( .A(n48606), .B(n2328), .Y(n48610) );
  NOR2X1 U50704 ( .A(n42672), .B(n39647), .Y(n48608) );
  NAND2X1 U50705 ( .A(n48608), .B(n2334), .Y(n48609) );
  NAND2X1 U50706 ( .A(n48610), .B(n48609), .Y(n48617) );
  NOR2X1 U50707 ( .A(n42752), .B(n39647), .Y(n48613) );
  NAND2X1 U50708 ( .A(n48613), .B(n2326), .Y(n48615) );
  NAND2X1 U50709 ( .A(n2320), .B(n43072), .Y(n48614) );
  NAND2X1 U50710 ( .A(n48615), .B(n48614), .Y(n48616) );
  NOR2X1 U50711 ( .A(n48617), .B(n48616), .Y(n48618) );
  NAND2X1 U50712 ( .A(n48619), .B(n48618), .Y(n48620) );
  NOR2X1 U50713 ( .A(n48621), .B(n48620), .Y(n48622) );
  NAND2X1 U50714 ( .A(n48623), .B(n48622), .Y(n64080) );
  NAND2X1 U50715 ( .A(n42801), .B(n64080), .Y(n48624) );
  NOR2X1 U50716 ( .A(n42907), .B(n37271), .Y(n48626) );
  NOR2X1 U50717 ( .A(n49169), .B(n37272), .Y(n48625) );
  NOR2X1 U50718 ( .A(n48626), .B(n48625), .Y(n48628) );
  NAND2X1 U50719 ( .A(n2320), .B(n42706), .Y(n48627) );
  NAND2X1 U50720 ( .A(n48628), .B(n48627), .Y(n48675) );
  NAND2X1 U50721 ( .A(n2322), .B(n40519), .Y(n48630) );
  NAND2X1 U50722 ( .A(n2336), .B(n42626), .Y(n48629) );
  NAND2X1 U50723 ( .A(n48630), .B(n48629), .Y(n48636) );
  NOR2X1 U50724 ( .A(n42903), .B(n37099), .Y(n48632) );
  NOR2X1 U50725 ( .A(n49678), .B(n37102), .Y(n48631) );
  NOR2X1 U50726 ( .A(n48632), .B(n48631), .Y(n48634) );
  NAND2X1 U50727 ( .A(n2346), .B(n42621), .Y(n48633) );
  NAND2X1 U50728 ( .A(n48634), .B(n48633), .Y(n48635) );
  NOR2X1 U50729 ( .A(n48636), .B(n48635), .Y(n48646) );
  NAND2X1 U50730 ( .A(n2335), .B(n40426), .Y(n48638) );
  NAND2X1 U50731 ( .A(n2337), .B(n49685), .Y(n48637) );
  NAND2X1 U50732 ( .A(n48638), .B(n48637), .Y(n48644) );
  NOR2X1 U50733 ( .A(n42864), .B(n37101), .Y(n48640) );
  NOR2X1 U50734 ( .A(n38213), .B(n37103), .Y(n48639) );
  NOR2X1 U50735 ( .A(n48640), .B(n48639), .Y(n48642) );
  NAND2X1 U50736 ( .A(n2338), .B(n42681), .Y(n48641) );
  NAND2X1 U50737 ( .A(n48642), .B(n48641), .Y(n48643) );
  NOR2X1 U50738 ( .A(n48644), .B(n48643), .Y(n48645) );
  NAND2X1 U50739 ( .A(n48646), .B(n48645), .Y(n48666) );
  NAND2X1 U50740 ( .A(n2327), .B(n42777), .Y(n48648) );
  NAND2X1 U50741 ( .A(n2318), .B(n42819), .Y(n48647) );
  NAND2X1 U50742 ( .A(n48648), .B(n48647), .Y(n48654) );
  NOR2X1 U50743 ( .A(n36609), .B(n37100), .Y(n48650) );
  NOR2X1 U50744 ( .A(n42896), .B(n37104), .Y(n48649) );
  NOR2X1 U50745 ( .A(n48650), .B(n48649), .Y(n48652) );
  NAND2X1 U50746 ( .A(n2325), .B(n73368), .Y(n48651) );
  NAND2X1 U50747 ( .A(n48652), .B(n48651), .Y(n48653) );
  NOR2X1 U50748 ( .A(n48654), .B(n48653), .Y(n48664) );
  NAND2X1 U50749 ( .A(n2333), .B(n42781), .Y(n48656) );
  NAND2X1 U50750 ( .A(n2328), .B(n39319), .Y(n48655) );
  NAND2X1 U50751 ( .A(n48656), .B(n48655), .Y(n48662) );
  NOR2X1 U50752 ( .A(n42912), .B(n37105), .Y(n48658) );
  NOR2X1 U50753 ( .A(n42893), .B(n37106), .Y(n48657) );
  NOR2X1 U50754 ( .A(n48658), .B(n48657), .Y(n48660) );
  NAND2X1 U50755 ( .A(n2329), .B(n40514), .Y(n48659) );
  NAND2X1 U50756 ( .A(n48660), .B(n48659), .Y(n48661) );
  NOR2X1 U50757 ( .A(n48662), .B(n48661), .Y(n48663) );
  NAND2X1 U50758 ( .A(n48664), .B(n48663), .Y(n48665) );
  NOR2X1 U50759 ( .A(n48666), .B(n48665), .Y(n48667) );
  NOR2X1 U50760 ( .A(n48667), .B(n42885), .Y(n48669) );
  NOR2X1 U50761 ( .A(n42915), .B(n37275), .Y(n48668) );
  NOR2X1 U50762 ( .A(n48669), .B(n48668), .Y(n48673) );
  NOR2X1 U50763 ( .A(n39335), .B(n37274), .Y(n48671) );
  NOR2X1 U50764 ( .A(n39572), .B(n37277), .Y(n48670) );
  NOR2X1 U50765 ( .A(n48671), .B(n48670), .Y(n48672) );
  NAND2X1 U50766 ( .A(n48673), .B(n48672), .Y(n48674) );
  NOR2X1 U50767 ( .A(n39354), .B(n37273), .Y(n48678) );
  NOR2X1 U50768 ( .A(n43108), .B(n42899), .Y(n48677) );
  NOR2X1 U50769 ( .A(n48678), .B(n48677), .Y(n48680) );
  NAND2X1 U50770 ( .A(writeback_exec_value_w[6]), .B(n43020), .Y(n48679) );
  NAND2X1 U50771 ( .A(n48680), .B(n48679), .Y(n48688) );
  NOR2X1 U50772 ( .A(n49710), .B(n37276), .Y(n48682) );
  NOR2X1 U50773 ( .A(n42913), .B(n37280), .Y(n48681) );
  NOR2X1 U50774 ( .A(n48682), .B(n48681), .Y(n48686) );
  NOR2X1 U50775 ( .A(n40855), .B(n37278), .Y(n48684) );
  NOR2X1 U50776 ( .A(n42919), .B(n37281), .Y(n48683) );
  NOR2X1 U50777 ( .A(n48684), .B(n48683), .Y(n48685) );
  NAND2X1 U50778 ( .A(n48686), .B(n48685), .Y(n48687) );
  NAND2X1 U50779 ( .A(n43845), .B(n43791), .Y(n57640) );
  NAND2X1 U50780 ( .A(n39944), .B(n38611), .Y(n48689) );
  NOR2X1 U50781 ( .A(n43746), .B(n43467), .Y(n48692) );
  NAND2X1 U50782 ( .A(n43768), .B(n48690), .Y(n48691) );
  NAND2X1 U50783 ( .A(n48692), .B(n48691), .Y(n48693) );
  NAND2X1 U50784 ( .A(n42068), .B(n48693), .Y(n48694) );
  NOR2X1 U50785 ( .A(n48695), .B(n48694), .Y(n48832) );
  OR2X1 U50786 ( .A(n35027), .B(n35026), .Y(n48697) );
  OR2X1 U50787 ( .A(n35029), .B(n35028), .Y(n48696) );
  NOR2X1 U50788 ( .A(n43103), .B(n43455), .Y(n48699) );
  NOR2X1 U50789 ( .A(n43021), .B(n43106), .Y(n48698) );
  NOR2X1 U50790 ( .A(n48699), .B(n48698), .Y(n48762) );
  NAND2X1 U50791 ( .A(n2610), .B(n43361), .Y(n48701) );
  NAND2X1 U50792 ( .A(n2586), .B(n38406), .Y(n48700) );
  NAND2X1 U50793 ( .A(n48701), .B(n48700), .Y(n48705) );
  NAND2X1 U50794 ( .A(n2592), .B(n43343), .Y(n48703) );
  NAND2X1 U50795 ( .A(n2600), .B(n43028), .Y(n48702) );
  NAND2X1 U50796 ( .A(n48703), .B(n48702), .Y(n48704) );
  NOR2X1 U50797 ( .A(n48705), .B(n48704), .Y(n48713) );
  NAND2X1 U50798 ( .A(n1821), .B(n43029), .Y(n48707) );
  NAND2X1 U50799 ( .A(n2588), .B(n43033), .Y(n48706) );
  NAND2X1 U50800 ( .A(n48707), .B(n48706), .Y(n48711) );
  NAND2X1 U50801 ( .A(n2602), .B(n43037), .Y(n48709) );
  NAND2X1 U50802 ( .A(n2594), .B(n43352), .Y(n48708) );
  NAND2X1 U50803 ( .A(n48709), .B(n48708), .Y(n48710) );
  NOR2X1 U50804 ( .A(n48711), .B(n48710), .Y(n48712) );
  NAND2X1 U50805 ( .A(n48713), .B(n48712), .Y(n48729) );
  NAND2X1 U50806 ( .A(n2598), .B(n41786), .Y(n48715) );
  NAND2X1 U50807 ( .A(n2596), .B(n43038), .Y(n48714) );
  NAND2X1 U50808 ( .A(n48715), .B(n48714), .Y(n48719) );
  NAND2X1 U50809 ( .A(n2612), .B(n39805), .Y(n48717) );
  NAND2X1 U50810 ( .A(n2604), .B(n43043), .Y(n48716) );
  NAND2X1 U50811 ( .A(n48717), .B(n48716), .Y(n48718) );
  NOR2X1 U50812 ( .A(n48719), .B(n48718), .Y(n48727) );
  NAND2X1 U50813 ( .A(n2608), .B(n43359), .Y(n48721) );
  NAND2X1 U50814 ( .A(n2583), .B(n43346), .Y(n48720) );
  NAND2X1 U50815 ( .A(n48721), .B(n48720), .Y(n48725) );
  NAND2X1 U50816 ( .A(n2590), .B(n43339), .Y(n48723) );
  NAND2X1 U50817 ( .A(n2606), .B(n43366), .Y(n48722) );
  NAND2X1 U50818 ( .A(n48723), .B(n48722), .Y(n48724) );
  NOR2X1 U50819 ( .A(n48725), .B(n48724), .Y(n48726) );
  NAND2X1 U50820 ( .A(n48727), .B(n48726), .Y(n48728) );
  NOR2X1 U50821 ( .A(n48729), .B(n48728), .Y(n48759) );
  NAND2X1 U50822 ( .A(n2603), .B(n43045), .Y(n48731) );
  NAND2X1 U50823 ( .A(n2609), .B(n43048), .Y(n48730) );
  NAND2X1 U50824 ( .A(n48731), .B(n48730), .Y(n48735) );
  NAND2X1 U50825 ( .A(n2601), .B(n49841), .Y(n48733) );
  NAND2X1 U50826 ( .A(n2587), .B(n43052), .Y(n48732) );
  NAND2X1 U50827 ( .A(n48733), .B(n48732), .Y(n48734) );
  NOR2X1 U50828 ( .A(n48735), .B(n48734), .Y(n48741) );
  NOR2X1 U50829 ( .A(n43371), .B(n36932), .Y(n48739) );
  NAND2X1 U50830 ( .A(n2589), .B(n43055), .Y(n48737) );
  NAND2X1 U50831 ( .A(n2611), .B(n43056), .Y(n48736) );
  NAND2X1 U50832 ( .A(n48737), .B(n48736), .Y(n48738) );
  NOR2X1 U50833 ( .A(n48739), .B(n48738), .Y(n48740) );
  NAND2X1 U50834 ( .A(n48741), .B(n48740), .Y(n48757) );
  NAND2X1 U50835 ( .A(n2607), .B(n43061), .Y(n48743) );
  NAND2X1 U50836 ( .A(n2605), .B(n39133), .Y(n48742) );
  NAND2X1 U50837 ( .A(n48743), .B(n48742), .Y(n48747) );
  NAND2X1 U50838 ( .A(n2597), .B(n43064), .Y(n48745) );
  NAND2X1 U50839 ( .A(n2585), .B(n43066), .Y(n48744) );
  NAND2X1 U50840 ( .A(n48745), .B(n48744), .Y(n48746) );
  NOR2X1 U50841 ( .A(n48747), .B(n48746), .Y(n48755) );
  NAND2X1 U50842 ( .A(n2593), .B(n43373), .Y(n48749) );
  NAND2X1 U50843 ( .A(n2599), .B(n40154), .Y(n48748) );
  NAND2X1 U50844 ( .A(n48749), .B(n48748), .Y(n48753) );
  NAND2X1 U50845 ( .A(n2591), .B(n43069), .Y(n48751) );
  NAND2X1 U50846 ( .A(n2584), .B(n43072), .Y(n48750) );
  NAND2X1 U50847 ( .A(n48751), .B(n48750), .Y(n48752) );
  NOR2X1 U50848 ( .A(n48753), .B(n48752), .Y(n48754) );
  NAND2X1 U50849 ( .A(n48755), .B(n48754), .Y(n48756) );
  NOR2X1 U50850 ( .A(n48757), .B(n48756), .Y(n48758) );
  NAND2X1 U50851 ( .A(n48759), .B(n48758), .Y(n48760) );
  NAND2X1 U50852 ( .A(n42802), .B(n48760), .Y(n48761) );
  NOR2X1 U50853 ( .A(n43794), .B(n38384), .Y(n48830) );
  NOR2X1 U50854 ( .A(n42908), .B(n37195), .Y(n48764) );
  NOR2X1 U50855 ( .A(n40041), .B(n37200), .Y(n48763) );
  NOR2X1 U50856 ( .A(n48764), .B(n48763), .Y(n48766) );
  NAND2X1 U50857 ( .A(n2584), .B(n42707), .Y(n48765) );
  NAND2X1 U50858 ( .A(n48766), .B(n48765), .Y(n48813) );
  NAND2X1 U50859 ( .A(n2587), .B(n40520), .Y(n48768) );
  NAND2X1 U50860 ( .A(n2601), .B(n42627), .Y(n48767) );
  NAND2X1 U50861 ( .A(n48768), .B(n48767), .Y(n48774) );
  NOR2X1 U50862 ( .A(n45640), .B(n36916), .Y(n48770) );
  NOR2X1 U50863 ( .A(n49678), .B(n36925), .Y(n48769) );
  NOR2X1 U50864 ( .A(n48770), .B(n48769), .Y(n48772) );
  NAND2X1 U50865 ( .A(n48772), .B(n48771), .Y(n48773) );
  NOR2X1 U50866 ( .A(n48774), .B(n48773), .Y(n48784) );
  NAND2X1 U50867 ( .A(n2600), .B(n40424), .Y(n48776) );
  NAND2X1 U50868 ( .A(n2602), .B(n49685), .Y(n48775) );
  NAND2X1 U50869 ( .A(n48776), .B(n48775), .Y(n48782) );
  NOR2X1 U50870 ( .A(n42864), .B(n36923), .Y(n48778) );
  NOR2X1 U50871 ( .A(n42859), .B(n36933), .Y(n48777) );
  NOR2X1 U50872 ( .A(n48778), .B(n48777), .Y(n48780) );
  NAND2X1 U50873 ( .A(n2603), .B(n42681), .Y(n48779) );
  NAND2X1 U50874 ( .A(n48780), .B(n48779), .Y(n48781) );
  NOR2X1 U50875 ( .A(n48782), .B(n48781), .Y(n48783) );
  NAND2X1 U50876 ( .A(n48784), .B(n48783), .Y(n48804) );
  NAND2X1 U50877 ( .A(n2592), .B(n38740), .Y(n48786) );
  NAND2X1 U50878 ( .A(n2583), .B(n38708), .Y(n48785) );
  NAND2X1 U50879 ( .A(n48786), .B(n48785), .Y(n48792) );
  NOR2X1 U50880 ( .A(n42891), .B(n36922), .Y(n48788) );
  NOR2X1 U50881 ( .A(n45651), .B(n36932), .Y(n48787) );
  NOR2X1 U50882 ( .A(n48788), .B(n48787), .Y(n48790) );
  NAND2X1 U50883 ( .A(n2590), .B(n46174), .Y(n48789) );
  NAND2X1 U50884 ( .A(n48790), .B(n48789), .Y(n48791) );
  NOR2X1 U50885 ( .A(n48792), .B(n48791), .Y(n48802) );
  NAND2X1 U50886 ( .A(n2598), .B(n39645), .Y(n48794) );
  NAND2X1 U50887 ( .A(n2593), .B(n39319), .Y(n48793) );
  NAND2X1 U50888 ( .A(n48794), .B(n48793), .Y(n48800) );
  NOR2X1 U50889 ( .A(n45507), .B(n36934), .Y(n48796) );
  NOR2X1 U50890 ( .A(n38166), .B(n42784), .Y(n48795) );
  NOR2X1 U50891 ( .A(n48796), .B(n48795), .Y(n48798) );
  NAND2X1 U50892 ( .A(n2594), .B(n40514), .Y(n48797) );
  NAND2X1 U50893 ( .A(n48798), .B(n48797), .Y(n48799) );
  NOR2X1 U50894 ( .A(n48800), .B(n48799), .Y(n48801) );
  NAND2X1 U50895 ( .A(n48802), .B(n48801), .Y(n48803) );
  NOR2X1 U50896 ( .A(n48804), .B(n48803), .Y(n48805) );
  NOR2X1 U50897 ( .A(n48805), .B(n42886), .Y(n48807) );
  NOR2X1 U50898 ( .A(n42916), .B(n37209), .Y(n48806) );
  NOR2X1 U50899 ( .A(n48807), .B(n48806), .Y(n48811) );
  NOR2X1 U50900 ( .A(n40277), .B(n37207), .Y(n48809) );
  NOR2X1 U50901 ( .A(n49624), .B(n37214), .Y(n48808) );
  NOR2X1 U50902 ( .A(n48809), .B(n48808), .Y(n48810) );
  NAND2X1 U50903 ( .A(n48811), .B(n48810), .Y(n48812) );
  NOR2X1 U50904 ( .A(n40407), .B(n37202), .Y(n48815) );
  NOR2X1 U50905 ( .A(n43103), .B(n42899), .Y(n48814) );
  NOR2X1 U50906 ( .A(n48815), .B(n48814), .Y(n48817) );
  NAND2X1 U50907 ( .A(writeback_exec_value_w[7]), .B(n38805), .Y(n48816) );
  NAND2X1 U50908 ( .A(n48817), .B(n48816), .Y(n48825) );
  NOR2X1 U50909 ( .A(n42909), .B(n37208), .Y(n48819) );
  NOR2X1 U50910 ( .A(n48819), .B(n48818), .Y(n48823) );
  NOR2X1 U50911 ( .A(n49637), .B(n37212), .Y(n48821) );
  NOR2X1 U50912 ( .A(n42917), .B(n37216), .Y(n48820) );
  NOR2X1 U50913 ( .A(n48821), .B(n48820), .Y(n48822) );
  NAND2X1 U50914 ( .A(n48823), .B(n48822), .Y(n48824) );
  NAND2X1 U50915 ( .A(n43792), .B(n43781), .Y(n48827) );
  NAND2X1 U50916 ( .A(n43847), .B(n38387), .Y(n48826) );
  NAND2X1 U50917 ( .A(n43847), .B(n39164), .Y(n48828) );
  NAND2X1 U50918 ( .A(n42069), .B(n48828), .Y(n48829) );
  NOR2X1 U50919 ( .A(n48830), .B(n48829), .Y(n48831) );
  NOR2X1 U50920 ( .A(n48832), .B(n48831), .Y(n48965) );
  NAND2X1 U50921 ( .A(mem_d_data_rd_i[24]), .B(n73578), .Y(n48833) );
  NAND2X1 U50922 ( .A(n34489), .B(n48833), .Y(n48834) );
  NOR2X1 U50923 ( .A(n43098), .B(n43455), .Y(n48836) );
  NOR2X1 U50924 ( .A(n43021), .B(n43101), .Y(n48835) );
  NOR2X1 U50925 ( .A(n48836), .B(n48835), .Y(n48899) );
  NAND2X1 U50926 ( .A(n2745), .B(n43361), .Y(n48838) );
  NAND2X1 U50927 ( .A(n2721), .B(n38408), .Y(n48837) );
  NAND2X1 U50928 ( .A(n48838), .B(n48837), .Y(n48842) );
  NAND2X1 U50929 ( .A(n2727), .B(n43342), .Y(n48840) );
  NAND2X1 U50930 ( .A(n2735), .B(n43028), .Y(n48839) );
  NAND2X1 U50931 ( .A(n48840), .B(n48839), .Y(n48841) );
  NOR2X1 U50932 ( .A(n48842), .B(n48841), .Y(n48850) );
  NAND2X1 U50933 ( .A(n1817), .B(n43029), .Y(n48844) );
  NAND2X1 U50934 ( .A(n2723), .B(n43033), .Y(n48843) );
  NAND2X1 U50935 ( .A(n48844), .B(n48843), .Y(n48848) );
  NAND2X1 U50936 ( .A(n2737), .B(n43037), .Y(n48846) );
  NAND2X1 U50937 ( .A(n2729), .B(n43352), .Y(n48845) );
  NAND2X1 U50938 ( .A(n48846), .B(n48845), .Y(n48847) );
  NOR2X1 U50939 ( .A(n48848), .B(n48847), .Y(n48849) );
  NAND2X1 U50940 ( .A(n48850), .B(n48849), .Y(n48866) );
  NAND2X1 U50941 ( .A(n2733), .B(n41786), .Y(n48852) );
  NAND2X1 U50942 ( .A(n2731), .B(n40169), .Y(n48851) );
  NAND2X1 U50943 ( .A(n48852), .B(n48851), .Y(n48856) );
  NAND2X1 U50944 ( .A(n2747), .B(n39806), .Y(n48854) );
  NAND2X1 U50945 ( .A(n2739), .B(n43043), .Y(n48853) );
  NAND2X1 U50946 ( .A(n48854), .B(n48853), .Y(n48855) );
  NOR2X1 U50947 ( .A(n48856), .B(n48855), .Y(n48864) );
  NAND2X1 U50948 ( .A(n2743), .B(n43358), .Y(n48858) );
  NAND2X1 U50949 ( .A(n2718), .B(n43346), .Y(n48857) );
  NAND2X1 U50950 ( .A(n48858), .B(n48857), .Y(n48862) );
  NAND2X1 U50951 ( .A(n2725), .B(n43339), .Y(n48860) );
  NAND2X1 U50952 ( .A(n2741), .B(n43366), .Y(n48859) );
  NAND2X1 U50953 ( .A(n48860), .B(n48859), .Y(n48861) );
  NOR2X1 U50954 ( .A(n48862), .B(n48861), .Y(n48863) );
  NAND2X1 U50955 ( .A(n48864), .B(n48863), .Y(n48865) );
  NOR2X1 U50956 ( .A(n48866), .B(n48865), .Y(n48896) );
  NAND2X1 U50957 ( .A(n2738), .B(n43045), .Y(n48868) );
  NAND2X1 U50958 ( .A(n2744), .B(n43048), .Y(n48867) );
  NAND2X1 U50959 ( .A(n48868), .B(n48867), .Y(n48872) );
  NAND2X1 U50960 ( .A(n2736), .B(n49841), .Y(n48870) );
  NAND2X1 U50961 ( .A(n2722), .B(n43052), .Y(n48869) );
  NAND2X1 U50962 ( .A(n48870), .B(n48869), .Y(n48871) );
  NOR2X1 U50963 ( .A(n48872), .B(n48871), .Y(n48878) );
  NOR2X1 U50964 ( .A(n43370), .B(n37066), .Y(n48876) );
  NAND2X1 U50965 ( .A(n2724), .B(n43055), .Y(n48874) );
  NAND2X1 U50966 ( .A(n2746), .B(n43056), .Y(n48873) );
  NAND2X1 U50967 ( .A(n48874), .B(n48873), .Y(n48875) );
  NOR2X1 U50968 ( .A(n48876), .B(n48875), .Y(n48877) );
  NAND2X1 U50969 ( .A(n48878), .B(n48877), .Y(n48894) );
  NAND2X1 U50970 ( .A(n2742), .B(n43061), .Y(n48880) );
  NAND2X1 U50971 ( .A(n2740), .B(n39134), .Y(n48879) );
  NAND2X1 U50972 ( .A(n48880), .B(n48879), .Y(n48884) );
  NAND2X1 U50973 ( .A(n2732), .B(n43064), .Y(n48882) );
  NAND2X1 U50974 ( .A(n2720), .B(n43066), .Y(n48881) );
  NAND2X1 U50975 ( .A(n48882), .B(n48881), .Y(n48883) );
  NOR2X1 U50976 ( .A(n48884), .B(n48883), .Y(n48892) );
  NAND2X1 U50977 ( .A(n2728), .B(n43373), .Y(n48886) );
  NAND2X1 U50978 ( .A(n2734), .B(n40154), .Y(n48885) );
  NAND2X1 U50979 ( .A(n48886), .B(n48885), .Y(n48890) );
  NAND2X1 U50980 ( .A(n2726), .B(n43069), .Y(n48888) );
  NAND2X1 U50981 ( .A(n2719), .B(n43072), .Y(n48887) );
  NAND2X1 U50982 ( .A(n48888), .B(n48887), .Y(n48889) );
  NOR2X1 U50983 ( .A(n48890), .B(n48889), .Y(n48891) );
  NAND2X1 U50984 ( .A(n48892), .B(n48891), .Y(n48893) );
  NOR2X1 U50985 ( .A(n48894), .B(n48893), .Y(n48895) );
  NAND2X1 U50986 ( .A(n48896), .B(n48895), .Y(n48897) );
  NAND2X1 U50987 ( .A(n42803), .B(n48897), .Y(n48898) );
  NOR2X1 U50988 ( .A(n49625), .B(n37241), .Y(n48901) );
  NOR2X1 U50989 ( .A(n40042), .B(n37243), .Y(n48900) );
  NOR2X1 U50990 ( .A(n48901), .B(n48900), .Y(n48903) );
  NAND2X1 U50991 ( .A(n2719), .B(n42707), .Y(n48902) );
  NAND2X1 U50992 ( .A(n48903), .B(n48902), .Y(n48950) );
  NAND2X1 U50993 ( .A(n2722), .B(n40520), .Y(n48905) );
  NAND2X1 U50994 ( .A(n2736), .B(n42626), .Y(n48904) );
  NAND2X1 U50995 ( .A(n48905), .B(n48904), .Y(n48911) );
  NOR2X1 U50996 ( .A(n42902), .B(n37049), .Y(n48907) );
  NOR2X1 U50997 ( .A(n42905), .B(n37059), .Y(n48906) );
  NOR2X1 U50998 ( .A(n48907), .B(n48906), .Y(n48909) );
  NAND2X1 U50999 ( .A(n2746), .B(n42618), .Y(n48908) );
  NAND2X1 U51000 ( .A(n48909), .B(n48908), .Y(n48910) );
  NOR2X1 U51001 ( .A(n48911), .B(n48910), .Y(n48921) );
  NAND2X1 U51002 ( .A(n2735), .B(n40425), .Y(n48913) );
  NAND2X1 U51003 ( .A(n2737), .B(n40535), .Y(n48912) );
  NAND2X1 U51004 ( .A(n48913), .B(n48912), .Y(n48919) );
  NOR2X1 U51005 ( .A(n42647), .B(n37056), .Y(n48915) );
  NOR2X1 U51006 ( .A(n42858), .B(n37063), .Y(n48914) );
  NOR2X1 U51007 ( .A(n48915), .B(n48914), .Y(n48917) );
  NAND2X1 U51008 ( .A(n2738), .B(n42679), .Y(n48916) );
  NAND2X1 U51009 ( .A(n48917), .B(n48916), .Y(n48918) );
  NOR2X1 U51010 ( .A(n48919), .B(n48918), .Y(n48920) );
  NAND2X1 U51011 ( .A(n48921), .B(n48920), .Y(n48941) );
  NAND2X1 U51012 ( .A(n2727), .B(n42778), .Y(n48923) );
  NAND2X1 U51013 ( .A(n48923), .B(n48922), .Y(n48929) );
  NOR2X1 U51014 ( .A(n36609), .B(n37058), .Y(n48925) );
  NOR2X1 U51015 ( .A(n42895), .B(n37066), .Y(n48924) );
  NOR2X1 U51016 ( .A(n48925), .B(n48924), .Y(n48927) );
  NAND2X1 U51017 ( .A(n2725), .B(n73368), .Y(n48926) );
  NAND2X1 U51018 ( .A(n48927), .B(n48926), .Y(n48928) );
  NOR2X1 U51019 ( .A(n48929), .B(n48928), .Y(n48939) );
  NAND2X1 U51020 ( .A(n2733), .B(n39645), .Y(n48931) );
  NAND2X1 U51021 ( .A(n2728), .B(n39318), .Y(n48930) );
  NAND2X1 U51022 ( .A(n48931), .B(n48930), .Y(n48937) );
  NOR2X1 U51023 ( .A(n45507), .B(n37065), .Y(n48933) );
  NOR2X1 U51024 ( .A(n40497), .B(n37072), .Y(n48932) );
  NOR2X1 U51025 ( .A(n48933), .B(n48932), .Y(n48935) );
  NAND2X1 U51026 ( .A(n2729), .B(n57613), .Y(n48934) );
  NAND2X1 U51027 ( .A(n48935), .B(n48934), .Y(n48936) );
  NOR2X1 U51028 ( .A(n48937), .B(n48936), .Y(n48938) );
  NAND2X1 U51029 ( .A(n48939), .B(n48938), .Y(n48940) );
  NOR2X1 U51030 ( .A(n48941), .B(n48940), .Y(n48942) );
  NOR2X1 U51031 ( .A(n48942), .B(n42887), .Y(n48944) );
  NOR2X1 U51032 ( .A(n42914), .B(n37246), .Y(n48943) );
  NOR2X1 U51033 ( .A(n48944), .B(n48943), .Y(n48948) );
  NOR2X1 U51034 ( .A(n39335), .B(n37245), .Y(n48946) );
  NOR2X1 U51035 ( .A(n42901), .B(n37248), .Y(n48945) );
  NOR2X1 U51036 ( .A(n48946), .B(n48945), .Y(n48947) );
  NAND2X1 U51037 ( .A(n48948), .B(n48947), .Y(n48949) );
  NOR2X1 U51038 ( .A(n48950), .B(n48949), .Y(n48964) );
  NOR2X1 U51039 ( .A(n42900), .B(n37242), .Y(n48952) );
  NOR2X1 U51040 ( .A(n43098), .B(n42899), .Y(n48951) );
  NOR2X1 U51041 ( .A(n48952), .B(n48951), .Y(n48954) );
  NAND2X1 U51042 ( .A(writeback_exec_value_w[8]), .B(n43020), .Y(n48953) );
  NAND2X1 U51043 ( .A(n48954), .B(n48953), .Y(n48962) );
  NOR2X1 U51044 ( .A(n42910), .B(n37244), .Y(n48956) );
  NOR2X1 U51045 ( .A(n38932), .B(n37249), .Y(n48955) );
  NOR2X1 U51046 ( .A(n48956), .B(n48955), .Y(n48960) );
  NOR2X1 U51047 ( .A(n42911), .B(n37247), .Y(n48958) );
  NOR2X1 U51048 ( .A(n42918), .B(n37250), .Y(n48957) );
  NOR2X1 U51049 ( .A(n48958), .B(n48957), .Y(n48959) );
  NAND2X1 U51050 ( .A(n48960), .B(n48959), .Y(n48961) );
  NOR2X1 U51051 ( .A(n48962), .B(n48961), .Y(n48963) );
  NAND2X1 U51052 ( .A(n48964), .B(n48963), .Y(n72760) );
  NAND2X1 U51053 ( .A(n44040), .B(n43737), .Y(n57639) );
  NAND2X1 U51054 ( .A(n38386), .B(n39163), .Y(n57636) );
  NAND2X1 U51055 ( .A(n57639), .B(n57636), .Y(n57757) );
  NOR2X1 U51056 ( .A(n48965), .B(n57757), .Y(n48966) );
  NAND2X1 U51057 ( .A(n43855), .B(n43758), .Y(n57672) );
  NOR2X1 U51058 ( .A(n42195), .B(n48967), .Y(n49101) );
  NAND2X1 U51059 ( .A(mem_d_data_rd_i[10]), .B(n31921), .Y(n48968) );
  NAND2X1 U51060 ( .A(n34489), .B(n48968), .Y(n48969) );
  NOR2X1 U51061 ( .A(n43125), .B(n43455), .Y(n48971) );
  NOR2X1 U51062 ( .A(n43021), .B(n43128), .Y(n48970) );
  NOR2X1 U51063 ( .A(n48971), .B(n48970), .Y(n49034) );
  NAND2X1 U51064 ( .A(n2379), .B(n43361), .Y(n48973) );
  NAND2X1 U51065 ( .A(n2355), .B(n38412), .Y(n48972) );
  NAND2X1 U51066 ( .A(n48973), .B(n48972), .Y(n48977) );
  NAND2X1 U51067 ( .A(n2361), .B(n38402), .Y(n48975) );
  NAND2X1 U51068 ( .A(n2369), .B(n38602), .Y(n48974) );
  NAND2X1 U51069 ( .A(n48975), .B(n48974), .Y(n48976) );
  NOR2X1 U51070 ( .A(n48977), .B(n48976), .Y(n48985) );
  NAND2X1 U51071 ( .A(n1830), .B(n38599), .Y(n48979) );
  NAND2X1 U51072 ( .A(n2357), .B(n43033), .Y(n48978) );
  NAND2X1 U51073 ( .A(n48979), .B(n48978), .Y(n48983) );
  NAND2X1 U51074 ( .A(n2371), .B(n43037), .Y(n48981) );
  NAND2X1 U51075 ( .A(n2363), .B(n43352), .Y(n48980) );
  NAND2X1 U51076 ( .A(n48981), .B(n48980), .Y(n48982) );
  NOR2X1 U51077 ( .A(n48983), .B(n48982), .Y(n48984) );
  NAND2X1 U51078 ( .A(n48985), .B(n48984), .Y(n49001) );
  NAND2X1 U51079 ( .A(n2367), .B(n43354), .Y(n48987) );
  NAND2X1 U51080 ( .A(n2365), .B(n40169), .Y(n48986) );
  NAND2X1 U51081 ( .A(n48987), .B(n48986), .Y(n48991) );
  NAND2X1 U51082 ( .A(n2381), .B(n39807), .Y(n48989) );
  NAND2X1 U51083 ( .A(n2373), .B(n43043), .Y(n48988) );
  NAND2X1 U51084 ( .A(n48989), .B(n48988), .Y(n48990) );
  NOR2X1 U51085 ( .A(n48991), .B(n48990), .Y(n48999) );
  NAND2X1 U51086 ( .A(n2377), .B(n38390), .Y(n48993) );
  NAND2X1 U51087 ( .A(n2352), .B(n43346), .Y(n48992) );
  NAND2X1 U51088 ( .A(n48993), .B(n48992), .Y(n48997) );
  NAND2X1 U51089 ( .A(n2359), .B(n43339), .Y(n48995) );
  NAND2X1 U51090 ( .A(n2375), .B(n43366), .Y(n48994) );
  NAND2X1 U51091 ( .A(n48995), .B(n48994), .Y(n48996) );
  NOR2X1 U51092 ( .A(n48997), .B(n48996), .Y(n48998) );
  NAND2X1 U51093 ( .A(n48999), .B(n48998), .Y(n49000) );
  NOR2X1 U51094 ( .A(n49001), .B(n49000), .Y(n49031) );
  NAND2X1 U51095 ( .A(n2372), .B(n40273), .Y(n49003) );
  NAND2X1 U51096 ( .A(n2378), .B(n43048), .Y(n49002) );
  NAND2X1 U51097 ( .A(n49003), .B(n49002), .Y(n49007) );
  NAND2X1 U51098 ( .A(n2370), .B(n49841), .Y(n49005) );
  NAND2X1 U51099 ( .A(n2356), .B(n43052), .Y(n49004) );
  NAND2X1 U51100 ( .A(n49005), .B(n49004), .Y(n49006) );
  NOR2X1 U51101 ( .A(n49007), .B(n49006), .Y(n49013) );
  NOR2X1 U51102 ( .A(n43370), .B(n37085), .Y(n49011) );
  NAND2X1 U51103 ( .A(n2358), .B(n38577), .Y(n49009) );
  NAND2X1 U51104 ( .A(n2380), .B(n40026), .Y(n49008) );
  NAND2X1 U51105 ( .A(n49009), .B(n49008), .Y(n49010) );
  NOR2X1 U51106 ( .A(n49011), .B(n49010), .Y(n49012) );
  NAND2X1 U51107 ( .A(n49013), .B(n49012), .Y(n49029) );
  NAND2X1 U51108 ( .A(n2376), .B(n43061), .Y(n49015) );
  NAND2X1 U51109 ( .A(n2374), .B(n39138), .Y(n49014) );
  NAND2X1 U51110 ( .A(n49015), .B(n49014), .Y(n49019) );
  NAND2X1 U51111 ( .A(n2366), .B(n40158), .Y(n49017) );
  NAND2X1 U51112 ( .A(n2354), .B(n38573), .Y(n49016) );
  NAND2X1 U51113 ( .A(n49017), .B(n49016), .Y(n49018) );
  NOR2X1 U51114 ( .A(n49019), .B(n49018), .Y(n49027) );
  NAND2X1 U51115 ( .A(n2362), .B(n43373), .Y(n49021) );
  NAND2X1 U51116 ( .A(n2368), .B(n43349), .Y(n49020) );
  NAND2X1 U51117 ( .A(n49021), .B(n49020), .Y(n49025) );
  NAND2X1 U51118 ( .A(n2360), .B(n43069), .Y(n49023) );
  NAND2X1 U51119 ( .A(n2353), .B(n43072), .Y(n49022) );
  NAND2X1 U51120 ( .A(n49023), .B(n49022), .Y(n49024) );
  NOR2X1 U51121 ( .A(n49025), .B(n49024), .Y(n49026) );
  NAND2X1 U51122 ( .A(n49027), .B(n49026), .Y(n49028) );
  NOR2X1 U51123 ( .A(n49029), .B(n49028), .Y(n49030) );
  NAND2X1 U51124 ( .A(n49031), .B(n49030), .Y(n49032) );
  NAND2X1 U51125 ( .A(n42806), .B(n49032), .Y(n49033) );
  NOR2X1 U51126 ( .A(n42907), .B(n37251), .Y(n49036) );
  NOR2X1 U51127 ( .A(n40041), .B(n37253), .Y(n49035) );
  NOR2X1 U51128 ( .A(n49036), .B(n49035), .Y(n49038) );
  NAND2X1 U51129 ( .A(n2353), .B(n42707), .Y(n49037) );
  NAND2X1 U51130 ( .A(n49038), .B(n49037), .Y(n49085) );
  NAND2X1 U51131 ( .A(n2356), .B(n40519), .Y(n49040) );
  NAND2X1 U51132 ( .A(n2370), .B(n42626), .Y(n49039) );
  NAND2X1 U51133 ( .A(n49040), .B(n49039), .Y(n49046) );
  NOR2X1 U51134 ( .A(n49677), .B(n37075), .Y(n49042) );
  NOR2X1 U51135 ( .A(n42906), .B(n37079), .Y(n49041) );
  NOR2X1 U51136 ( .A(n49042), .B(n49041), .Y(n49044) );
  NAND2X1 U51137 ( .A(n2380), .B(n42621), .Y(n49043) );
  NAND2X1 U51138 ( .A(n49044), .B(n49043), .Y(n49045) );
  NOR2X1 U51139 ( .A(n49046), .B(n49045), .Y(n49056) );
  NAND2X1 U51140 ( .A(n2369), .B(n40425), .Y(n49048) );
  NAND2X1 U51141 ( .A(n2371), .B(n49685), .Y(n49047) );
  NAND2X1 U51142 ( .A(n49048), .B(n49047), .Y(n49054) );
  NOR2X1 U51143 ( .A(n42647), .B(n37077), .Y(n49050) );
  NOR2X1 U51144 ( .A(n38213), .B(n37081), .Y(n49049) );
  NOR2X1 U51145 ( .A(n49050), .B(n49049), .Y(n49052) );
  NAND2X1 U51146 ( .A(n2372), .B(n42680), .Y(n49051) );
  NAND2X1 U51147 ( .A(n49052), .B(n49051), .Y(n49053) );
  NOR2X1 U51148 ( .A(n49054), .B(n49053), .Y(n49055) );
  NAND2X1 U51149 ( .A(n49056), .B(n49055), .Y(n49076) );
  NAND2X1 U51150 ( .A(n2361), .B(n42778), .Y(n49058) );
  NAND2X1 U51151 ( .A(n49058), .B(n49057), .Y(n49064) );
  NOR2X1 U51152 ( .A(n36609), .B(n37078), .Y(n49060) );
  NOR2X1 U51153 ( .A(n42896), .B(n37085), .Y(n49059) );
  NOR2X1 U51154 ( .A(n49060), .B(n49059), .Y(n49062) );
  NAND2X1 U51155 ( .A(n2359), .B(n42675), .Y(n49061) );
  NAND2X1 U51156 ( .A(n49062), .B(n49061), .Y(n49063) );
  NOR2X1 U51157 ( .A(n49064), .B(n49063), .Y(n49074) );
  NAND2X1 U51158 ( .A(n2367), .B(n42781), .Y(n49066) );
  NAND2X1 U51159 ( .A(n2362), .B(n39319), .Y(n49065) );
  NAND2X1 U51160 ( .A(n49066), .B(n49065), .Y(n49072) );
  NOR2X1 U51161 ( .A(n40857), .B(n37084), .Y(n49068) );
  NOR2X1 U51162 ( .A(n40851), .B(n37089), .Y(n49067) );
  NOR2X1 U51163 ( .A(n49068), .B(n49067), .Y(n49070) );
  NAND2X1 U51164 ( .A(n2363), .B(n57613), .Y(n49069) );
  NAND2X1 U51165 ( .A(n49070), .B(n49069), .Y(n49071) );
  NOR2X1 U51166 ( .A(n49072), .B(n49071), .Y(n49073) );
  NAND2X1 U51167 ( .A(n49074), .B(n49073), .Y(n49075) );
  NOR2X1 U51168 ( .A(n49076), .B(n49075), .Y(n49077) );
  NOR2X1 U51169 ( .A(n49077), .B(n42890), .Y(n49079) );
  NOR2X1 U51170 ( .A(n40847), .B(n37256), .Y(n49078) );
  NOR2X1 U51171 ( .A(n49079), .B(n49078), .Y(n49083) );
  NOR2X1 U51172 ( .A(n39335), .B(n37257), .Y(n49081) );
  NOR2X1 U51173 ( .A(n42901), .B(n37261), .Y(n49080) );
  NOR2X1 U51174 ( .A(n49081), .B(n49080), .Y(n49082) );
  NAND2X1 U51175 ( .A(n49083), .B(n49082), .Y(n49084) );
  NOR2X1 U51176 ( .A(n49085), .B(n49084), .Y(n49099) );
  NOR2X1 U51177 ( .A(n39353), .B(n37254), .Y(n49087) );
  NOR2X1 U51178 ( .A(n43125), .B(n40360), .Y(n49086) );
  NOR2X1 U51179 ( .A(n49087), .B(n49086), .Y(n49089) );
  NAND2X1 U51180 ( .A(writeback_exec_value_w[10]), .B(n43020), .Y(n49088) );
  NAND2X1 U51181 ( .A(n49089), .B(n49088), .Y(n49097) );
  NOR2X1 U51182 ( .A(n49710), .B(n37255), .Y(n49091) );
  NOR2X1 U51183 ( .A(n42913), .B(n37262), .Y(n49090) );
  NOR2X1 U51184 ( .A(n49091), .B(n49090), .Y(n49095) );
  NOR2X1 U51185 ( .A(n49637), .B(n37260), .Y(n49093) );
  NOR2X1 U51186 ( .A(n42919), .B(n37265), .Y(n49092) );
  NOR2X1 U51187 ( .A(n49093), .B(n49092), .Y(n49094) );
  NAND2X1 U51188 ( .A(n49095), .B(n49094), .Y(n49096) );
  NOR2X1 U51189 ( .A(n49097), .B(n49096), .Y(n49098) );
  NAND2X1 U51190 ( .A(n49099), .B(n49098), .Y(n72825) );
  NAND2X1 U51191 ( .A(n43864), .B(n43821), .Y(n57673) );
  INVX1 U51192 ( .A(n57673), .Y(n49100) );
  NOR2X1 U51193 ( .A(n49101), .B(n49100), .Y(n49239) );
  NAND2X1 U51194 ( .A(mem_d_data_rd_i[11]), .B(n31921), .Y(n49102) );
  NAND2X1 U51195 ( .A(n34489), .B(n49102), .Y(n49103) );
  NOR2X1 U51196 ( .A(n43130), .B(n43455), .Y(n49105) );
  NOR2X1 U51197 ( .A(n43021), .B(n43133), .Y(n49104) );
  NOR2X1 U51198 ( .A(n49105), .B(n49104), .Y(n49168) );
  NAND2X1 U51199 ( .A(n2280), .B(n43361), .Y(n49107) );
  NAND2X1 U51200 ( .A(n2256), .B(n38411), .Y(n49106) );
  NAND2X1 U51201 ( .A(n49107), .B(n49106), .Y(n49111) );
  NAND2X1 U51202 ( .A(n2262), .B(n43344), .Y(n49109) );
  NAND2X1 U51203 ( .A(n2270), .B(n38602), .Y(n49108) );
  NAND2X1 U51204 ( .A(n49109), .B(n49108), .Y(n49110) );
  NOR2X1 U51205 ( .A(n49111), .B(n49110), .Y(n49119) );
  NAND2X1 U51206 ( .A(n1835), .B(n38599), .Y(n49113) );
  NAND2X1 U51207 ( .A(n2258), .B(n43033), .Y(n49112) );
  NAND2X1 U51208 ( .A(n49113), .B(n49112), .Y(n49117) );
  NAND2X1 U51209 ( .A(n2272), .B(n38534), .Y(n49115) );
  NAND2X1 U51210 ( .A(n2264), .B(n43352), .Y(n49114) );
  NAND2X1 U51211 ( .A(n49115), .B(n49114), .Y(n49116) );
  NOR2X1 U51212 ( .A(n49117), .B(n49116), .Y(n49118) );
  NAND2X1 U51213 ( .A(n49119), .B(n49118), .Y(n49135) );
  NAND2X1 U51214 ( .A(n2268), .B(n43355), .Y(n49121) );
  NAND2X1 U51215 ( .A(n2266), .B(n40169), .Y(n49120) );
  NAND2X1 U51216 ( .A(n49121), .B(n49120), .Y(n49125) );
  NAND2X1 U51217 ( .A(n2282), .B(n39808), .Y(n49123) );
  NAND2X1 U51218 ( .A(n2274), .B(n43043), .Y(n49122) );
  NAND2X1 U51219 ( .A(n49123), .B(n49122), .Y(n49124) );
  NOR2X1 U51220 ( .A(n49125), .B(n49124), .Y(n49133) );
  NAND2X1 U51221 ( .A(n2278), .B(n43360), .Y(n49127) );
  NAND2X1 U51222 ( .A(n2253), .B(n43346), .Y(n49126) );
  NAND2X1 U51223 ( .A(n49127), .B(n49126), .Y(n49131) );
  NAND2X1 U51224 ( .A(n2260), .B(n43339), .Y(n49129) );
  NAND2X1 U51225 ( .A(n2276), .B(n43366), .Y(n49128) );
  NAND2X1 U51226 ( .A(n49129), .B(n49128), .Y(n49130) );
  NOR2X1 U51227 ( .A(n49131), .B(n49130), .Y(n49132) );
  NAND2X1 U51228 ( .A(n49133), .B(n49132), .Y(n49134) );
  NOR2X1 U51229 ( .A(n49135), .B(n49134), .Y(n49165) );
  NAND2X1 U51230 ( .A(n2273), .B(n40273), .Y(n49137) );
  NAND2X1 U51231 ( .A(n2279), .B(n43048), .Y(n49136) );
  NAND2X1 U51232 ( .A(n49137), .B(n49136), .Y(n49141) );
  NAND2X1 U51233 ( .A(n2271), .B(n43050), .Y(n49139) );
  NAND2X1 U51234 ( .A(n2257), .B(n43052), .Y(n49138) );
  NAND2X1 U51235 ( .A(n49139), .B(n49138), .Y(n49140) );
  NOR2X1 U51236 ( .A(n49141), .B(n49140), .Y(n49147) );
  NOR2X1 U51237 ( .A(n43370), .B(n36977), .Y(n49145) );
  NAND2X1 U51238 ( .A(n2259), .B(n38577), .Y(n49143) );
  NAND2X1 U51239 ( .A(n2281), .B(n40026), .Y(n49142) );
  NAND2X1 U51240 ( .A(n49143), .B(n49142), .Y(n49144) );
  NOR2X1 U51241 ( .A(n49145), .B(n49144), .Y(n49146) );
  NAND2X1 U51242 ( .A(n49147), .B(n49146), .Y(n49163) );
  NAND2X1 U51243 ( .A(n2277), .B(n43061), .Y(n49149) );
  NAND2X1 U51244 ( .A(n2275), .B(n39137), .Y(n49148) );
  NAND2X1 U51245 ( .A(n49149), .B(n49148), .Y(n49153) );
  NAND2X1 U51246 ( .A(n2267), .B(n40158), .Y(n49151) );
  NAND2X1 U51247 ( .A(n2255), .B(n38573), .Y(n49150) );
  NAND2X1 U51248 ( .A(n49151), .B(n49150), .Y(n49152) );
  NOR2X1 U51249 ( .A(n49153), .B(n49152), .Y(n49161) );
  NAND2X1 U51250 ( .A(n2263), .B(n38528), .Y(n49155) );
  NAND2X1 U51251 ( .A(n2269), .B(n43349), .Y(n49154) );
  NAND2X1 U51252 ( .A(n49155), .B(n49154), .Y(n49159) );
  NAND2X1 U51253 ( .A(n2261), .B(n43069), .Y(n49157) );
  NAND2X1 U51254 ( .A(n2254), .B(n43072), .Y(n49156) );
  NAND2X1 U51255 ( .A(n49157), .B(n49156), .Y(n49158) );
  NOR2X1 U51256 ( .A(n49159), .B(n49158), .Y(n49160) );
  NAND2X1 U51257 ( .A(n49161), .B(n49160), .Y(n49162) );
  NOR2X1 U51258 ( .A(n49163), .B(n49162), .Y(n49164) );
  NAND2X1 U51259 ( .A(n49165), .B(n49164), .Y(n49166) );
  NAND2X1 U51260 ( .A(n42801), .B(n49166), .Y(n49167) );
  NOR2X1 U51261 ( .A(n43822), .B(n43965), .Y(n49237) );
  NOR2X1 U51262 ( .A(n42908), .B(n37224), .Y(n49171) );
  NOR2X1 U51263 ( .A(n37221), .B(n49169), .Y(n49170) );
  NOR2X1 U51264 ( .A(n49171), .B(n49170), .Y(n49173) );
  NAND2X1 U51265 ( .A(n2254), .B(n42706), .Y(n49172) );
  NAND2X1 U51266 ( .A(n49173), .B(n49172), .Y(n49220) );
  NAND2X1 U51267 ( .A(n2257), .B(n40519), .Y(n49175) );
  NAND2X1 U51268 ( .A(n2271), .B(n42626), .Y(n49174) );
  NAND2X1 U51269 ( .A(n49175), .B(n49174), .Y(n49181) );
  NOR2X1 U51270 ( .A(n45640), .B(n36943), .Y(n49177) );
  NOR2X1 U51271 ( .A(n38753), .B(n36967), .Y(n49176) );
  NOR2X1 U51272 ( .A(n49177), .B(n49176), .Y(n49179) );
  NAND2X1 U51273 ( .A(n2281), .B(n42620), .Y(n49178) );
  NAND2X1 U51274 ( .A(n49179), .B(n49178), .Y(n49180) );
  NOR2X1 U51275 ( .A(n49181), .B(n49180), .Y(n49191) );
  NAND2X1 U51276 ( .A(n2270), .B(n40426), .Y(n49183) );
  NAND2X1 U51277 ( .A(n2272), .B(n40535), .Y(n49182) );
  NAND2X1 U51278 ( .A(n49183), .B(n49182), .Y(n49189) );
  NOR2X1 U51279 ( .A(n42865), .B(n36963), .Y(n49185) );
  NOR2X1 U51280 ( .A(n42858), .B(n36974), .Y(n49184) );
  NOR2X1 U51281 ( .A(n49185), .B(n49184), .Y(n49187) );
  NAND2X1 U51282 ( .A(n2273), .B(n42679), .Y(n49186) );
  NAND2X1 U51283 ( .A(n49187), .B(n49186), .Y(n49188) );
  NOR2X1 U51284 ( .A(n49189), .B(n49188), .Y(n49190) );
  NAND2X1 U51285 ( .A(n49191), .B(n49190), .Y(n49211) );
  NAND2X1 U51286 ( .A(n2262), .B(n42777), .Y(n49193) );
  NAND2X1 U51287 ( .A(n2253), .B(n38708), .Y(n49192) );
  NAND2X1 U51288 ( .A(n49193), .B(n49192), .Y(n49199) );
  NOR2X1 U51289 ( .A(n42891), .B(n36956), .Y(n49195) );
  NOR2X1 U51290 ( .A(n42895), .B(n36977), .Y(n49194) );
  NOR2X1 U51291 ( .A(n49195), .B(n49194), .Y(n49197) );
  NAND2X1 U51292 ( .A(n2260), .B(n46174), .Y(n49196) );
  NAND2X1 U51293 ( .A(n49197), .B(n49196), .Y(n49198) );
  NOR2X1 U51294 ( .A(n49199), .B(n49198), .Y(n49209) );
  NAND2X1 U51295 ( .A(n2268), .B(n39645), .Y(n49201) );
  NAND2X1 U51296 ( .A(n2263), .B(n39318), .Y(n49200) );
  NAND2X1 U51297 ( .A(n49201), .B(n49200), .Y(n49207) );
  NOR2X1 U51298 ( .A(n49665), .B(n36976), .Y(n49203) );
  NOR2X1 U51299 ( .A(n42893), .B(n36994), .Y(n49202) );
  NOR2X1 U51300 ( .A(n49203), .B(n49202), .Y(n49205) );
  NAND2X1 U51301 ( .A(n2264), .B(n40515), .Y(n49204) );
  NAND2X1 U51302 ( .A(n49205), .B(n49204), .Y(n49206) );
  NOR2X1 U51303 ( .A(n49207), .B(n49206), .Y(n49208) );
  NAND2X1 U51304 ( .A(n49209), .B(n49208), .Y(n49210) );
  NOR2X1 U51305 ( .A(n49211), .B(n49210), .Y(n49212) );
  NOR2X1 U51306 ( .A(n49212), .B(n42885), .Y(n49214) );
  NOR2X1 U51307 ( .A(n40847), .B(n37229), .Y(n49213) );
  NOR2X1 U51308 ( .A(n49214), .B(n49213), .Y(n49218) );
  NOR2X1 U51309 ( .A(n40277), .B(n37230), .Y(n49216) );
  NOR2X1 U51310 ( .A(n49624), .B(n37232), .Y(n49215) );
  NOR2X1 U51311 ( .A(n49216), .B(n49215), .Y(n49217) );
  NAND2X1 U51312 ( .A(n49218), .B(n49217), .Y(n49219) );
  NOR2X1 U51313 ( .A(n40406), .B(n37223), .Y(n49222) );
  NOR2X1 U51314 ( .A(n43130), .B(n40360), .Y(n49221) );
  NOR2X1 U51315 ( .A(n49222), .B(n49221), .Y(n49224) );
  NAND2X1 U51316 ( .A(writeback_exec_value_w[11]), .B(n43020), .Y(n49223) );
  NAND2X1 U51317 ( .A(n49224), .B(n49223), .Y(n49232) );
  NOR2X1 U51318 ( .A(n42909), .B(n37225), .Y(n49226) );
  NOR2X1 U51319 ( .A(n42913), .B(n37228), .Y(n49225) );
  NOR2X1 U51320 ( .A(n49226), .B(n49225), .Y(n49230) );
  NOR2X1 U51321 ( .A(n40855), .B(n37227), .Y(n49228) );
  NOR2X1 U51322 ( .A(n42917), .B(n37231), .Y(n49227) );
  NOR2X1 U51323 ( .A(n49228), .B(n49227), .Y(n49229) );
  NAND2X1 U51324 ( .A(n49230), .B(n49229), .Y(n49231) );
  NAND2X1 U51325 ( .A(n43820), .B(n72820), .Y(n49234) );
  NAND2X1 U51326 ( .A(n43866), .B(n43968), .Y(n49233) );
  NAND2X1 U51327 ( .A(n43866), .B(n43812), .Y(n49235) );
  NAND2X1 U51328 ( .A(n42084), .B(n49235), .Y(n49236) );
  NOR2X1 U51329 ( .A(n49237), .B(n49236), .Y(n49238) );
  NOR2X1 U51330 ( .A(n49239), .B(n49238), .Y(n49371) );
  NAND2X1 U51331 ( .A(n43967), .B(n43812), .Y(n49370) );
  NAND2X1 U51332 ( .A(mem_d_data_rd_i[12]), .B(n31921), .Y(n49240) );
  NAND2X1 U51333 ( .A(n34489), .B(n49240), .Y(n49241) );
  NOR2X1 U51334 ( .A(n43136), .B(n43455), .Y(n49243) );
  NOR2X1 U51335 ( .A(n43021), .B(n43139), .Y(n49242) );
  NOR2X1 U51336 ( .A(n49243), .B(n49242), .Y(n49306) );
  NAND2X1 U51337 ( .A(n2714), .B(n43361), .Y(n49245) );
  NAND2X1 U51338 ( .A(n2689), .B(n38410), .Y(n49244) );
  NAND2X1 U51339 ( .A(n49245), .B(n49244), .Y(n49249) );
  NAND2X1 U51340 ( .A(n2696), .B(n43343), .Y(n49247) );
  NAND2X1 U51341 ( .A(n2704), .B(n38602), .Y(n49246) );
  NAND2X1 U51342 ( .A(n49247), .B(n49246), .Y(n49248) );
  NOR2X1 U51343 ( .A(n49249), .B(n49248), .Y(n49257) );
  NAND2X1 U51344 ( .A(n2686), .B(n38599), .Y(n49251) );
  NAND2X1 U51345 ( .A(n2692), .B(n43033), .Y(n49250) );
  NAND2X1 U51346 ( .A(n49251), .B(n49250), .Y(n49255) );
  NAND2X1 U51347 ( .A(n2706), .B(n38534), .Y(n49253) );
  NAND2X1 U51348 ( .A(n2698), .B(n43352), .Y(n49252) );
  NAND2X1 U51349 ( .A(n49253), .B(n49252), .Y(n49254) );
  NOR2X1 U51350 ( .A(n49255), .B(n49254), .Y(n49256) );
  NAND2X1 U51351 ( .A(n49257), .B(n49256), .Y(n49273) );
  NAND2X1 U51352 ( .A(n2702), .B(n43355), .Y(n49259) );
  NAND2X1 U51353 ( .A(n2700), .B(n40169), .Y(n49258) );
  NAND2X1 U51354 ( .A(n49259), .B(n49258), .Y(n49263) );
  NAND2X1 U51355 ( .A(n1818), .B(n39807), .Y(n49261) );
  NAND2X1 U51356 ( .A(n2708), .B(n43043), .Y(n49260) );
  NAND2X1 U51357 ( .A(n49261), .B(n49260), .Y(n49262) );
  NOR2X1 U51358 ( .A(n49263), .B(n49262), .Y(n49271) );
  NAND2X1 U51359 ( .A(n2712), .B(n43359), .Y(n49265) );
  NAND2X1 U51360 ( .A(n2687), .B(n43346), .Y(n49264) );
  NAND2X1 U51361 ( .A(n49265), .B(n49264), .Y(n49269) );
  NAND2X1 U51362 ( .A(n2694), .B(n43339), .Y(n49267) );
  NAND2X1 U51363 ( .A(n2710), .B(n43366), .Y(n49266) );
  NAND2X1 U51364 ( .A(n49267), .B(n49266), .Y(n49268) );
  NOR2X1 U51365 ( .A(n49269), .B(n49268), .Y(n49270) );
  NAND2X1 U51366 ( .A(n49271), .B(n49270), .Y(n49272) );
  NOR2X1 U51367 ( .A(n49273), .B(n49272), .Y(n49303) );
  NAND2X1 U51368 ( .A(n2707), .B(n40273), .Y(n49275) );
  NAND2X1 U51369 ( .A(n2713), .B(n43048), .Y(n49274) );
  NAND2X1 U51370 ( .A(n49275), .B(n49274), .Y(n49279) );
  NAND2X1 U51371 ( .A(n2705), .B(n43050), .Y(n49277) );
  NAND2X1 U51372 ( .A(n2691), .B(n43052), .Y(n49276) );
  NAND2X1 U51373 ( .A(n49277), .B(n49276), .Y(n49278) );
  NOR2X1 U51374 ( .A(n49279), .B(n49278), .Y(n49285) );
  NOR2X1 U51375 ( .A(n43371), .B(n36928), .Y(n49283) );
  NAND2X1 U51376 ( .A(n2693), .B(n38577), .Y(n49281) );
  NAND2X1 U51377 ( .A(n2715), .B(n40026), .Y(n49280) );
  NAND2X1 U51378 ( .A(n49281), .B(n49280), .Y(n49282) );
  NOR2X1 U51379 ( .A(n49283), .B(n49282), .Y(n49284) );
  NAND2X1 U51380 ( .A(n49285), .B(n49284), .Y(n49301) );
  NAND2X1 U51381 ( .A(n2711), .B(n43061), .Y(n49287) );
  NAND2X1 U51382 ( .A(n2709), .B(n39136), .Y(n49286) );
  NAND2X1 U51383 ( .A(n49287), .B(n49286), .Y(n49291) );
  NAND2X1 U51384 ( .A(n2701), .B(n40158), .Y(n49289) );
  NAND2X1 U51385 ( .A(n2690), .B(n38573), .Y(n49288) );
  NAND2X1 U51386 ( .A(n49289), .B(n49288), .Y(n49290) );
  NOR2X1 U51387 ( .A(n49291), .B(n49290), .Y(n49299) );
  NAND2X1 U51388 ( .A(n2697), .B(n38528), .Y(n49293) );
  NAND2X1 U51389 ( .A(n2703), .B(n43350), .Y(n49292) );
  NAND2X1 U51390 ( .A(n49293), .B(n49292), .Y(n49297) );
  NAND2X1 U51391 ( .A(n2695), .B(n43069), .Y(n49295) );
  NAND2X1 U51392 ( .A(n2688), .B(n43072), .Y(n49294) );
  NAND2X1 U51393 ( .A(n49295), .B(n49294), .Y(n49296) );
  NOR2X1 U51394 ( .A(n49297), .B(n49296), .Y(n49298) );
  NAND2X1 U51395 ( .A(n49299), .B(n49298), .Y(n49300) );
  NOR2X1 U51396 ( .A(n49301), .B(n49300), .Y(n49302) );
  NAND2X1 U51397 ( .A(n49303), .B(n49302), .Y(n49304) );
  NAND2X1 U51398 ( .A(n42805), .B(n49304), .Y(n49305) );
  NOR2X1 U51399 ( .A(n49625), .B(n37194), .Y(n49308) );
  NOR2X1 U51400 ( .A(n38798), .B(n37199), .Y(n49307) );
  NOR2X1 U51401 ( .A(n49308), .B(n49307), .Y(n49310) );
  NAND2X1 U51402 ( .A(n2688), .B(n49647), .Y(n49309) );
  NAND2X1 U51403 ( .A(n49310), .B(n49309), .Y(n49357) );
  NAND2X1 U51404 ( .A(n2691), .B(n49674), .Y(n49312) );
  NAND2X1 U51405 ( .A(n2705), .B(n42627), .Y(n49311) );
  NAND2X1 U51406 ( .A(n49312), .B(n49311), .Y(n49318) );
  NOR2X1 U51407 ( .A(n45640), .B(n36914), .Y(n49314) );
  NOR2X1 U51408 ( .A(n38753), .B(n36924), .Y(n49313) );
  NOR2X1 U51409 ( .A(n49314), .B(n49313), .Y(n49316) );
  NAND2X1 U51410 ( .A(n2715), .B(n42619), .Y(n49315) );
  NAND2X1 U51411 ( .A(n49316), .B(n49315), .Y(n49317) );
  NOR2X1 U51412 ( .A(n49318), .B(n49317), .Y(n49328) );
  NAND2X1 U51413 ( .A(n2704), .B(n40426), .Y(n49320) );
  NAND2X1 U51414 ( .A(n2706), .B(n40536), .Y(n49319) );
  NAND2X1 U51415 ( .A(n49320), .B(n49319), .Y(n49326) );
  NOR2X1 U51416 ( .A(n45870), .B(n36920), .Y(n49322) );
  NOR2X1 U51417 ( .A(n42859), .B(n36929), .Y(n49321) );
  NOR2X1 U51418 ( .A(n49322), .B(n49321), .Y(n49324) );
  NAND2X1 U51419 ( .A(n2707), .B(n42679), .Y(n49323) );
  NAND2X1 U51420 ( .A(n49324), .B(n49323), .Y(n49325) );
  NOR2X1 U51421 ( .A(n49326), .B(n49325), .Y(n49327) );
  NAND2X1 U51422 ( .A(n49328), .B(n49327), .Y(n49348) );
  NAND2X1 U51423 ( .A(n2696), .B(n42778), .Y(n49330) );
  NAND2X1 U51424 ( .A(n2687), .B(n38709), .Y(n49329) );
  NAND2X1 U51425 ( .A(n49330), .B(n49329), .Y(n49336) );
  NOR2X1 U51426 ( .A(n36609), .B(n36921), .Y(n49332) );
  NOR2X1 U51427 ( .A(n45651), .B(n36928), .Y(n49331) );
  NOR2X1 U51428 ( .A(n49332), .B(n49331), .Y(n49334) );
  NAND2X1 U51429 ( .A(n2694), .B(n42675), .Y(n49333) );
  NAND2X1 U51430 ( .A(n49334), .B(n49333), .Y(n49335) );
  NOR2X1 U51431 ( .A(n49336), .B(n49335), .Y(n49346) );
  NAND2X1 U51432 ( .A(n2702), .B(n42781), .Y(n49338) );
  NAND2X1 U51433 ( .A(n2697), .B(n40537), .Y(n49337) );
  NAND2X1 U51434 ( .A(n49338), .B(n49337), .Y(n49344) );
  NOR2X1 U51435 ( .A(n40857), .B(n36930), .Y(n49340) );
  NOR2X1 U51436 ( .A(n42893), .B(n36937), .Y(n49339) );
  NOR2X1 U51437 ( .A(n49340), .B(n49339), .Y(n49342) );
  NAND2X1 U51438 ( .A(n2698), .B(n57613), .Y(n49341) );
  NAND2X1 U51439 ( .A(n49342), .B(n49341), .Y(n49343) );
  NOR2X1 U51440 ( .A(n49344), .B(n49343), .Y(n49345) );
  NAND2X1 U51441 ( .A(n49346), .B(n49345), .Y(n49347) );
  NOR2X1 U51442 ( .A(n49348), .B(n49347), .Y(n49349) );
  NOR2X1 U51443 ( .A(n49349), .B(n42886), .Y(n49351) );
  NOR2X1 U51444 ( .A(n40847), .B(n37203), .Y(n49350) );
  NOR2X1 U51445 ( .A(n49351), .B(n49350), .Y(n49355) );
  NOR2X1 U51446 ( .A(n40277), .B(n37204), .Y(n49353) );
  NOR2X1 U51447 ( .A(n42901), .B(n37206), .Y(n49352) );
  NOR2X1 U51448 ( .A(n49353), .B(n49352), .Y(n49354) );
  NAND2X1 U51449 ( .A(n49355), .B(n49354), .Y(n49356) );
  NOR2X1 U51450 ( .A(n42900), .B(n37197), .Y(n49359) );
  NOR2X1 U51451 ( .A(n43136), .B(n42899), .Y(n49358) );
  NOR2X1 U51452 ( .A(n49359), .B(n49358), .Y(n49361) );
  NAND2X1 U51453 ( .A(writeback_exec_value_w[12]), .B(n43020), .Y(n49360) );
  NAND2X1 U51454 ( .A(n49361), .B(n49360), .Y(n49369) );
  NOR2X1 U51455 ( .A(n42910), .B(n37205), .Y(n49363) );
  NOR2X1 U51456 ( .A(n42913), .B(n37213), .Y(n49362) );
  NOR2X1 U51457 ( .A(n49363), .B(n49362), .Y(n49367) );
  NOR2X1 U51458 ( .A(n40855), .B(n37210), .Y(n49365) );
  NOR2X1 U51459 ( .A(n42918), .B(n37215), .Y(n49364) );
  NOR2X1 U51460 ( .A(n49365), .B(n49364), .Y(n49366) );
  NAND2X1 U51461 ( .A(n49367), .B(n49366), .Y(n49368) );
  NAND2X1 U51462 ( .A(n43958), .B(n40461), .Y(n57801) );
  NAND2X1 U51463 ( .A(n49370), .B(n57801), .Y(n57661) );
  NOR2X1 U51464 ( .A(n49371), .B(n57661), .Y(n49497) );
  NOR2X1 U51465 ( .A(n42907), .B(n37182), .Y(n49373) );
  NOR2X1 U51466 ( .A(n40517), .B(n37183), .Y(n49372) );
  NOR2X1 U51467 ( .A(n49373), .B(n49372), .Y(n49375) );
  NAND2X1 U51468 ( .A(n2757), .B(n49647), .Y(n49374) );
  NAND2X1 U51469 ( .A(n49375), .B(n49374), .Y(n49413) );
  NOR2X1 U51470 ( .A(n45640), .B(n36838), .Y(n49377) );
  NOR2X1 U51471 ( .A(n38753), .B(n36849), .Y(n49376) );
  NOR2X1 U51472 ( .A(n49377), .B(n49376), .Y(n49379) );
  NAND2X1 U51473 ( .A(n49379), .B(n49378), .Y(n49380) );
  NAND2X1 U51474 ( .A(n2773), .B(n40425), .Y(n49383) );
  NAND2X1 U51475 ( .A(n2775), .B(n40535), .Y(n49382) );
  NAND2X1 U51476 ( .A(n49383), .B(n49382), .Y(n49389) );
  NOR2X1 U51477 ( .A(n42647), .B(n36850), .Y(n49385) );
  NOR2X1 U51478 ( .A(n42859), .B(n36855), .Y(n49384) );
  NOR2X1 U51479 ( .A(n49385), .B(n49384), .Y(n49387) );
  NAND2X1 U51480 ( .A(n2776), .B(n42678), .Y(n49386) );
  NAND2X1 U51481 ( .A(n49387), .B(n49386), .Y(n49388) );
  NAND2X1 U51482 ( .A(n2765), .B(n42778), .Y(n49391) );
  NAND2X1 U51483 ( .A(n2756), .B(n38709), .Y(n49390) );
  NAND2X1 U51484 ( .A(n49391), .B(n49390), .Y(n49397) );
  NOR2X1 U51485 ( .A(n36609), .B(n36844), .Y(n49393) );
  NOR2X1 U51486 ( .A(n42895), .B(n36853), .Y(n49392) );
  NOR2X1 U51487 ( .A(n49393), .B(n49392), .Y(n49395) );
  NAND2X1 U51488 ( .A(n2763), .B(n46174), .Y(n49394) );
  NAND2X1 U51489 ( .A(n49395), .B(n49394), .Y(n49396) );
  NAND2X1 U51490 ( .A(n2771), .B(n46177), .Y(n49399) );
  NAND2X1 U51491 ( .A(n2766), .B(n40537), .Y(n49398) );
  NAND2X1 U51492 ( .A(n49399), .B(n49398), .Y(n49402) );
  NOR2X1 U51493 ( .A(n49404), .B(n49403), .Y(n49405) );
  NOR2X1 U51494 ( .A(n49405), .B(n42887), .Y(n49407) );
  NOR2X1 U51495 ( .A(n40847), .B(n37186), .Y(n49406) );
  NOR2X1 U51496 ( .A(n49407), .B(n49406), .Y(n49411) );
  NOR2X1 U51497 ( .A(n39335), .B(n37185), .Y(n49409) );
  NOR2X1 U51498 ( .A(n42901), .B(n37189), .Y(n49408) );
  NOR2X1 U51499 ( .A(n49409), .B(n49408), .Y(n49410) );
  NAND2X1 U51500 ( .A(n49411), .B(n49410), .Y(n49412) );
  NOR2X1 U51501 ( .A(n39353), .B(n37184), .Y(n49417) );
  NAND2X1 U51502 ( .A(mem_d_data_rd_i[13]), .B(n31921), .Y(n49414) );
  NAND2X1 U51503 ( .A(n34489), .B(n49414), .Y(n49415) );
  NOR2X1 U51504 ( .A(n43086), .B(n42899), .Y(n49416) );
  NOR2X1 U51505 ( .A(n49417), .B(n49416), .Y(n49419) );
  NAND2X1 U51506 ( .A(writeback_exec_value_w[13]), .B(n43020), .Y(n49418) );
  NAND2X1 U51507 ( .A(n49419), .B(n49418), .Y(n49427) );
  NOR2X1 U51508 ( .A(n49710), .B(n37187), .Y(n49421) );
  NOR2X1 U51509 ( .A(n38932), .B(n37191), .Y(n49420) );
  NOR2X1 U51510 ( .A(n49421), .B(n49420), .Y(n49425) );
  NOR2X1 U51511 ( .A(n49637), .B(n37190), .Y(n49423) );
  NOR2X1 U51512 ( .A(n42919), .B(n37193), .Y(n49422) );
  NOR2X1 U51513 ( .A(n49423), .B(n49422), .Y(n49424) );
  NAND2X1 U51514 ( .A(n49425), .B(n49424), .Y(n49426) );
  NAND2X1 U51515 ( .A(n40476), .B(n40461), .Y(n57798) );
  INVX1 U51516 ( .A(n57798), .Y(n49495) );
  NOR2X1 U51517 ( .A(n43086), .B(n43455), .Y(n49429) );
  NOR2X1 U51518 ( .A(n43021), .B(n43089), .Y(n49428) );
  NAND2X1 U51519 ( .A(n2783), .B(n43361), .Y(n49431) );
  NAND2X1 U51520 ( .A(n2758), .B(n38412), .Y(n49430) );
  NAND2X1 U51521 ( .A(n49431), .B(n49430), .Y(n49435) );
  NAND2X1 U51522 ( .A(n2765), .B(n43342), .Y(n49433) );
  NAND2X1 U51523 ( .A(n2773), .B(n38602), .Y(n49432) );
  NAND2X1 U51524 ( .A(n49433), .B(n49432), .Y(n49434) );
  NOR2X1 U51525 ( .A(n49435), .B(n49434), .Y(n49443) );
  NAND2X1 U51526 ( .A(n2755), .B(n38599), .Y(n49437) );
  NAND2X1 U51527 ( .A(n2761), .B(n43033), .Y(n49436) );
  NAND2X1 U51528 ( .A(n49437), .B(n49436), .Y(n49441) );
  NAND2X1 U51529 ( .A(n2775), .B(n38534), .Y(n49439) );
  NAND2X1 U51530 ( .A(n2767), .B(n43352), .Y(n49438) );
  NAND2X1 U51531 ( .A(n49439), .B(n49438), .Y(n49440) );
  NOR2X1 U51532 ( .A(n49441), .B(n49440), .Y(n49442) );
  NAND2X1 U51533 ( .A(n49443), .B(n49442), .Y(n49459) );
  NAND2X1 U51534 ( .A(n2771), .B(n43354), .Y(n49445) );
  NAND2X1 U51535 ( .A(n2769), .B(n40169), .Y(n49444) );
  NAND2X1 U51536 ( .A(n49445), .B(n49444), .Y(n49449) );
  NAND2X1 U51537 ( .A(n1812), .B(n39808), .Y(n49447) );
  NAND2X1 U51538 ( .A(n2777), .B(n43043), .Y(n49446) );
  NAND2X1 U51539 ( .A(n49447), .B(n49446), .Y(n49448) );
  NOR2X1 U51540 ( .A(n49449), .B(n49448), .Y(n49457) );
  NAND2X1 U51541 ( .A(n2781), .B(n43358), .Y(n49451) );
  NAND2X1 U51542 ( .A(n2756), .B(n43346), .Y(n49450) );
  NAND2X1 U51543 ( .A(n49451), .B(n49450), .Y(n49455) );
  NAND2X1 U51544 ( .A(n2763), .B(n43339), .Y(n49453) );
  NAND2X1 U51545 ( .A(n2779), .B(n43366), .Y(n49452) );
  NAND2X1 U51546 ( .A(n49453), .B(n49452), .Y(n49454) );
  NOR2X1 U51547 ( .A(n49455), .B(n49454), .Y(n49456) );
  NAND2X1 U51548 ( .A(n49457), .B(n49456), .Y(n49458) );
  NOR2X1 U51549 ( .A(n49459), .B(n49458), .Y(n49489) );
  NAND2X1 U51550 ( .A(n2776), .B(n40273), .Y(n49461) );
  NAND2X1 U51551 ( .A(n2782), .B(n43048), .Y(n49460) );
  NAND2X1 U51552 ( .A(n49461), .B(n49460), .Y(n49465) );
  NAND2X1 U51553 ( .A(n2774), .B(n43050), .Y(n49463) );
  NAND2X1 U51554 ( .A(n2760), .B(n43052), .Y(n49462) );
  NAND2X1 U51555 ( .A(n49463), .B(n49462), .Y(n49464) );
  NOR2X1 U51556 ( .A(n49465), .B(n49464), .Y(n49471) );
  NOR2X1 U51557 ( .A(n43371), .B(n36853), .Y(n49469) );
  NAND2X1 U51558 ( .A(n2762), .B(n38577), .Y(n49467) );
  NAND2X1 U51559 ( .A(n2784), .B(n40026), .Y(n49466) );
  NAND2X1 U51560 ( .A(n49467), .B(n49466), .Y(n49468) );
  NOR2X1 U51561 ( .A(n49469), .B(n49468), .Y(n49470) );
  NAND2X1 U51562 ( .A(n49471), .B(n49470), .Y(n49487) );
  NAND2X1 U51563 ( .A(n2780), .B(n43061), .Y(n49473) );
  NAND2X1 U51564 ( .A(n2778), .B(n39138), .Y(n49472) );
  NAND2X1 U51565 ( .A(n49473), .B(n49472), .Y(n49477) );
  NAND2X1 U51566 ( .A(n2770), .B(n40158), .Y(n49475) );
  NAND2X1 U51567 ( .A(n2759), .B(n38573), .Y(n49474) );
  NAND2X1 U51568 ( .A(n49475), .B(n49474), .Y(n49476) );
  NOR2X1 U51569 ( .A(n49477), .B(n49476), .Y(n49485) );
  NAND2X1 U51570 ( .A(n2766), .B(n38528), .Y(n49479) );
  NAND2X1 U51571 ( .A(n2772), .B(n43349), .Y(n49478) );
  NAND2X1 U51572 ( .A(n49479), .B(n49478), .Y(n49483) );
  NAND2X1 U51573 ( .A(n2764), .B(n43069), .Y(n49481) );
  NAND2X1 U51574 ( .A(n2757), .B(n43072), .Y(n49480) );
  NAND2X1 U51575 ( .A(n49481), .B(n49480), .Y(n49482) );
  NOR2X1 U51576 ( .A(n49483), .B(n49482), .Y(n49484) );
  NAND2X1 U51577 ( .A(n49485), .B(n49484), .Y(n49486) );
  NOR2X1 U51578 ( .A(n49487), .B(n49486), .Y(n49488) );
  NAND2X1 U51579 ( .A(n49489), .B(n49488), .Y(n49490) );
  NAND2X1 U51580 ( .A(n43875), .B(n40468), .Y(n49492) );
  NAND2X1 U51581 ( .A(n43958), .B(n40475), .Y(n49491) );
  NAND2X1 U51582 ( .A(n49492), .B(n49491), .Y(n57800) );
  INVX1 U51583 ( .A(n57800), .Y(n49493) );
  NAND2X1 U51584 ( .A(n43875), .B(n43957), .Y(n57797) );
  NAND2X1 U51585 ( .A(n49493), .B(n57797), .Y(n49494) );
  NOR2X1 U51586 ( .A(n49495), .B(n49494), .Y(n49496) );
  NOR2X1 U51587 ( .A(n49497), .B(n49496), .Y(n49499) );
  NAND2X1 U51588 ( .A(n43885), .B(n40488), .Y(n57808) );
  INVX1 U51589 ( .A(n57808), .Y(n49498) );
  NOR2X1 U51590 ( .A(n49499), .B(n49498), .Y(n49500) );
  NAND2X1 U51591 ( .A(n43875), .B(n40470), .Y(n57809) );
  NAND2X1 U51592 ( .A(n49500), .B(n57809), .Y(n49501) );
  NAND2X1 U51593 ( .A(n73435), .B(n49501), .Y(n49502) );
  NAND2X1 U51594 ( .A(n57828), .B(n49502), .Y(n49503) );
  NOR2X1 U51595 ( .A(n57637), .B(n49503), .Y(n49504) );
  NAND2X1 U51596 ( .A(n43726), .B(n43899), .Y(n57831) );
  INVX1 U51597 ( .A(n57831), .Y(n57665) );
  NOR2X1 U51598 ( .A(n49504), .B(n57665), .Y(n49505) );
  NAND2X1 U51599 ( .A(n43908), .B(n42643), .Y(n57629) );
  INVX1 U51600 ( .A(n57629), .Y(n57840) );
  NOR2X1 U51601 ( .A(n49505), .B(n57840), .Y(n49506) );
  NOR2X1 U51602 ( .A(n57833), .B(n49506), .Y(n49646) );
  INVX1 U51603 ( .A(mem_d_data_rd_i[18]), .Y(n73551) );
  NAND2X1 U51604 ( .A(n40935), .B(n73551), .Y(n49507) );
  NOR2X1 U51605 ( .A(n43454), .B(n43160), .Y(n49509) );
  NOR2X1 U51606 ( .A(n43021), .B(n43163), .Y(n49508) );
  NOR2X1 U51607 ( .A(n49509), .B(n49508), .Y(n49572) );
  NAND2X1 U51608 ( .A(n2680), .B(n43361), .Y(n49511) );
  NAND2X1 U51609 ( .A(n2655), .B(n38408), .Y(n49510) );
  NAND2X1 U51610 ( .A(n49511), .B(n49510), .Y(n49515) );
  NAND2X1 U51611 ( .A(n2662), .B(n43342), .Y(n49513) );
  NAND2X1 U51612 ( .A(n2670), .B(n38602), .Y(n49512) );
  NAND2X1 U51613 ( .A(n49513), .B(n49512), .Y(n49514) );
  NOR2X1 U51614 ( .A(n49515), .B(n49514), .Y(n49523) );
  NAND2X1 U51615 ( .A(n2652), .B(n38599), .Y(n49517) );
  NAND2X1 U51616 ( .A(n2658), .B(n43034), .Y(n49516) );
  NAND2X1 U51617 ( .A(n49517), .B(n49516), .Y(n49521) );
  NAND2X1 U51618 ( .A(n2672), .B(n38534), .Y(n49519) );
  NAND2X1 U51619 ( .A(n2664), .B(n43352), .Y(n49518) );
  NAND2X1 U51620 ( .A(n49519), .B(n49518), .Y(n49520) );
  NOR2X1 U51621 ( .A(n49521), .B(n49520), .Y(n49522) );
  NAND2X1 U51622 ( .A(n49523), .B(n49522), .Y(n49539) );
  NAND2X1 U51623 ( .A(n2668), .B(n43355), .Y(n49525) );
  NAND2X1 U51624 ( .A(n2666), .B(n40169), .Y(n49524) );
  NAND2X1 U51625 ( .A(n49525), .B(n49524), .Y(n49529) );
  NAND2X1 U51626 ( .A(n1819), .B(n39804), .Y(n49527) );
  NAND2X1 U51627 ( .A(n2674), .B(n43043), .Y(n49526) );
  NAND2X1 U51628 ( .A(n49527), .B(n49526), .Y(n49528) );
  NOR2X1 U51629 ( .A(n49529), .B(n49528), .Y(n49537) );
  NAND2X1 U51630 ( .A(n2678), .B(n43358), .Y(n49531) );
  NAND2X1 U51631 ( .A(n2653), .B(n43347), .Y(n49530) );
  NAND2X1 U51632 ( .A(n49531), .B(n49530), .Y(n49535) );
  NAND2X1 U51633 ( .A(n2660), .B(n43340), .Y(n49533) );
  NAND2X1 U51634 ( .A(n2676), .B(n43367), .Y(n49532) );
  NAND2X1 U51635 ( .A(n49533), .B(n49532), .Y(n49534) );
  NOR2X1 U51636 ( .A(n49535), .B(n49534), .Y(n49536) );
  NAND2X1 U51637 ( .A(n49537), .B(n49536), .Y(n49538) );
  NOR2X1 U51638 ( .A(n49539), .B(n49538), .Y(n49569) );
  NAND2X1 U51639 ( .A(n2673), .B(n40273), .Y(n49541) );
  NAND2X1 U51640 ( .A(n2679), .B(n43048), .Y(n49540) );
  NAND2X1 U51641 ( .A(n49541), .B(n49540), .Y(n49545) );
  NAND2X1 U51642 ( .A(n2671), .B(n43050), .Y(n49543) );
  NAND2X1 U51643 ( .A(n2656), .B(n43053), .Y(n49542) );
  NAND2X1 U51644 ( .A(n49543), .B(n49542), .Y(n49544) );
  NOR2X1 U51645 ( .A(n49545), .B(n49544), .Y(n49551) );
  NOR2X1 U51646 ( .A(n43370), .B(n37315), .Y(n49549) );
  NAND2X1 U51647 ( .A(n2659), .B(n38577), .Y(n49547) );
  NAND2X1 U51648 ( .A(n2681), .B(n40026), .Y(n49546) );
  NAND2X1 U51649 ( .A(n49547), .B(n49546), .Y(n49548) );
  NOR2X1 U51650 ( .A(n49549), .B(n49548), .Y(n49550) );
  NAND2X1 U51651 ( .A(n49551), .B(n49550), .Y(n49567) );
  NAND2X1 U51652 ( .A(n2677), .B(n43062), .Y(n49553) );
  NAND2X1 U51653 ( .A(n2675), .B(n39134), .Y(n49552) );
  NAND2X1 U51654 ( .A(n49553), .B(n49552), .Y(n49557) );
  NAND2X1 U51655 ( .A(n2667), .B(n40158), .Y(n49555) );
  NAND2X1 U51656 ( .A(n2657), .B(n38573), .Y(n49554) );
  NAND2X1 U51657 ( .A(n49555), .B(n49554), .Y(n49556) );
  NOR2X1 U51658 ( .A(n49557), .B(n49556), .Y(n49565) );
  NAND2X1 U51659 ( .A(n2663), .B(n38528), .Y(n49559) );
  NAND2X1 U51660 ( .A(n2669), .B(n43349), .Y(n49558) );
  NAND2X1 U51661 ( .A(n49559), .B(n49558), .Y(n49563) );
  NAND2X1 U51662 ( .A(n2661), .B(n43069), .Y(n49561) );
  NAND2X1 U51663 ( .A(n2654), .B(n43073), .Y(n49560) );
  NAND2X1 U51664 ( .A(n49561), .B(n49560), .Y(n49562) );
  NOR2X1 U51665 ( .A(n49563), .B(n49562), .Y(n49564) );
  NAND2X1 U51666 ( .A(n49565), .B(n49564), .Y(n49566) );
  NOR2X1 U51667 ( .A(n49567), .B(n49566), .Y(n49568) );
  NAND2X1 U51668 ( .A(n49569), .B(n49568), .Y(n49570) );
  NAND2X1 U51669 ( .A(n42802), .B(n49570), .Y(n49571) );
  NAND2X1 U51670 ( .A(n49572), .B(n49571), .Y(n73232) );
  NOR2X1 U51671 ( .A(n46903), .B(n37124), .Y(n49575) );
  NOR2X1 U51672 ( .A(n42914), .B(n37129), .Y(n49574) );
  NOR2X1 U51673 ( .A(n49575), .B(n49574), .Y(n49623) );
  NOR2X1 U51674 ( .A(n42682), .B(n36906), .Y(n49581) );
  NOR2X1 U51675 ( .A(n40508), .B(n39195), .Y(n49577) );
  NAND2X1 U51676 ( .A(n49577), .B(n2679), .Y(n49579) );
  NAND2X1 U51677 ( .A(n46929), .B(n2658), .Y(n49578) );
  NAND2X1 U51678 ( .A(n49579), .B(n49578), .Y(n49580) );
  NOR2X1 U51679 ( .A(n49581), .B(n49580), .Y(n49586) );
  NOR2X1 U51680 ( .A(n45244), .B(n36908), .Y(n49584) );
  NOR2X1 U51681 ( .A(n40428), .B(n36918), .Y(n49583) );
  NOR2X1 U51682 ( .A(n49584), .B(n49583), .Y(n49585) );
  NOR2X1 U51683 ( .A(n42623), .B(n36912), .Y(n49592) );
  NAND2X1 U51684 ( .A(n46167), .B(n2678), .Y(n49590) );
  NAND2X1 U51685 ( .A(n46772), .B(n2680), .Y(n49589) );
  NAND2X1 U51686 ( .A(n49590), .B(n49589), .Y(n49591) );
  NOR2X1 U51687 ( .A(n49592), .B(n49591), .Y(n49598) );
  NOR2X1 U51688 ( .A(n42629), .B(n36919), .Y(n49596) );
  NOR2X1 U51689 ( .A(n39654), .B(n36926), .Y(n49595) );
  NOR2X1 U51690 ( .A(n49596), .B(n49595), .Y(n49597) );
  NOR2X1 U51691 ( .A(n49599), .B(n36911), .Y(n49603) );
  NAND2X1 U51692 ( .A(n2655), .B(n57621), .Y(n49601) );
  NAND2X1 U51693 ( .A(n46178), .B(n2676), .Y(n49600) );
  NAND2X1 U51694 ( .A(n49601), .B(n49600), .Y(n49602) );
  NOR2X1 U51695 ( .A(n49603), .B(n49602), .Y(n49609) );
  NOR2X1 U51696 ( .A(n49604), .B(n36917), .Y(n49607) );
  NOR2X1 U51697 ( .A(n38701), .B(n36927), .Y(n49606) );
  NOR2X1 U51698 ( .A(n49607), .B(n49606), .Y(n49608) );
  NAND2X1 U51699 ( .A(n49609), .B(n49608), .Y(n49619) );
  NAND2X1 U51700 ( .A(n2665), .B(n42821), .Y(n49613) );
  NAND2X1 U51701 ( .A(n2659), .B(n49611), .Y(n49612) );
  NOR2X1 U51702 ( .A(n38711), .B(n36931), .Y(n49615) );
  NOR2X1 U51703 ( .A(n42775), .B(n36939), .Y(n49614) );
  NOR2X1 U51704 ( .A(n49615), .B(n49614), .Y(n49616) );
  NAND2X1 U51705 ( .A(n49617), .B(n49616), .Y(n49618) );
  NAND2X1 U51706 ( .A(n40490), .B(n49620), .Y(n49622) );
  NAND2X1 U51707 ( .A(n49623), .B(n49622), .Y(n49629) );
  NOR2X1 U51708 ( .A(n49629), .B(n49628), .Y(n49645) );
  NOR2X1 U51709 ( .A(n40406), .B(n37125), .Y(n49632) );
  NOR2X1 U51710 ( .A(n43162), .B(n42899), .Y(n49631) );
  NOR2X1 U51711 ( .A(n49632), .B(n49631), .Y(n49634) );
  NAND2X1 U51712 ( .A(writeback_exec_value_w[18]), .B(n43020), .Y(n49633) );
  NAND2X1 U51713 ( .A(n49634), .B(n49633), .Y(n49643) );
  NOR2X1 U51714 ( .A(n42909), .B(n37121), .Y(n49636) );
  NOR2X1 U51715 ( .A(n46382), .B(n37126), .Y(n49635) );
  NOR2X1 U51716 ( .A(n49636), .B(n49635), .Y(n49641) );
  NOR2X1 U51717 ( .A(n40855), .B(n37123), .Y(n49639) );
  NOR2X1 U51718 ( .A(n42917), .B(n37128), .Y(n49638) );
  NOR2X1 U51719 ( .A(n49639), .B(n49638), .Y(n49640) );
  NAND2X1 U51720 ( .A(n49641), .B(n49640), .Y(n49642) );
  NOR2X1 U51721 ( .A(n49642), .B(n49643), .Y(n49644) );
  NAND2X1 U51722 ( .A(n43915), .B(n40259), .Y(n57630) );
  INVX1 U51723 ( .A(n57630), .Y(n57856) );
  NOR2X1 U51724 ( .A(n49646), .B(n57856), .Y(n49793) );
  NAND2X1 U51725 ( .A(n2288), .B(n42707), .Y(n49650) );
  NAND2X1 U51726 ( .A(n2311), .B(n49648), .Y(n49649) );
  NAND2X1 U51727 ( .A(n49650), .B(n49649), .Y(n49654) );
  NAND2X1 U51728 ( .A(n2308), .B(n42830), .Y(n49652) );
  NAND2X1 U51729 ( .A(n2295), .B(n40531), .Y(n49651) );
  NAND2X1 U51730 ( .A(n49652), .B(n49651), .Y(n49653) );
  NAND2X1 U51731 ( .A(n2296), .B(n42778), .Y(n49656) );
  NAND2X1 U51732 ( .A(n2287), .B(n38709), .Y(n49655) );
  NAND2X1 U51733 ( .A(n49656), .B(n49655), .Y(n49662) );
  NOR2X1 U51734 ( .A(n42891), .B(n36881), .Y(n49658) );
  NOR2X1 U51735 ( .A(n45651), .B(n36887), .Y(n49657) );
  NOR2X1 U51736 ( .A(n49658), .B(n49657), .Y(n49660) );
  NAND2X1 U51737 ( .A(n2294), .B(n42675), .Y(n49659) );
  NAND2X1 U51738 ( .A(n49660), .B(n49659), .Y(n49661) );
  NOR2X1 U51739 ( .A(n49662), .B(n49661), .Y(n49673) );
  NAND2X1 U51740 ( .A(n2302), .B(n40943), .Y(n49664) );
  NAND2X1 U51741 ( .A(n2297), .B(n39319), .Y(n49663) );
  NAND2X1 U51742 ( .A(n49664), .B(n49663), .Y(n49671) );
  NOR2X1 U51743 ( .A(n36884), .B(n45507), .Y(n49667) );
  NOR2X1 U51744 ( .A(n40497), .B(n36892), .Y(n49666) );
  NOR2X1 U51745 ( .A(n49667), .B(n49666), .Y(n49669) );
  NAND2X1 U51746 ( .A(n2298), .B(n40514), .Y(n49668) );
  NAND2X1 U51747 ( .A(n49669), .B(n49668), .Y(n49670) );
  NOR2X1 U51748 ( .A(n49671), .B(n49670), .Y(n49672) );
  NAND2X1 U51749 ( .A(n49673), .B(n49672), .Y(n49698) );
  NAND2X1 U51750 ( .A(n2290), .B(n40520), .Y(n49676) );
  NAND2X1 U51751 ( .A(n2305), .B(n42626), .Y(n49675) );
  NAND2X1 U51752 ( .A(n49676), .B(n49675), .Y(n49684) );
  NOR2X1 U51753 ( .A(n36886), .B(n42902), .Y(n49680) );
  NOR2X1 U51754 ( .A(n36891), .B(n42904), .Y(n49679) );
  NOR2X1 U51755 ( .A(n49680), .B(n49679), .Y(n49682) );
  NAND2X1 U51756 ( .A(n2315), .B(n42621), .Y(n49681) );
  NAND2X1 U51757 ( .A(n49682), .B(n49681), .Y(n49683) );
  NOR2X1 U51758 ( .A(n49684), .B(n49683), .Y(n49696) );
  NAND2X1 U51759 ( .A(n2304), .B(n40426), .Y(n49687) );
  NAND2X1 U51760 ( .A(n2306), .B(n40535), .Y(n49686) );
  NAND2X1 U51761 ( .A(n49687), .B(n49686), .Y(n49694) );
  NOR2X1 U51762 ( .A(n42647), .B(n36894), .Y(n49690) );
  NAND2X1 U51763 ( .A(n39197), .B(n40513), .Y(n49688) );
  NOR2X1 U51764 ( .A(n36896), .B(n49688), .Y(n49689) );
  NOR2X1 U51765 ( .A(n49690), .B(n49689), .Y(n49692) );
  NAND2X1 U51766 ( .A(n2307), .B(n42681), .Y(n49691) );
  NAND2X1 U51767 ( .A(n49692), .B(n49691), .Y(n49693) );
  NOR2X1 U51768 ( .A(n49694), .B(n49693), .Y(n49695) );
  NAND2X1 U51769 ( .A(n49696), .B(n49695), .Y(n49697) );
  NOR2X1 U51770 ( .A(n49698), .B(n49697), .Y(n49700) );
  NOR2X1 U51771 ( .A(n49700), .B(n42889), .Y(n49704) );
  NAND2X1 U51772 ( .A(n2301), .B(n41741), .Y(n49702) );
  NAND2X1 U51773 ( .A(n2309), .B(n40521), .Y(n49701) );
  NAND2X1 U51774 ( .A(n49702), .B(n49701), .Y(n49703) );
  NAND2X1 U51775 ( .A(n2291), .B(n49705), .Y(n49708) );
  NAND2X1 U51776 ( .A(n2286), .B(n49706), .Y(n49707) );
  NAND2X1 U51777 ( .A(n49708), .B(n49707), .Y(n49714) );
  NAND2X1 U51778 ( .A(n1834), .B(n49709), .Y(n49712) );
  NAND2X1 U51779 ( .A(n49712), .B(n49711), .Y(n49713) );
  NOR2X1 U51780 ( .A(n49715), .B(n43169), .Y(n49723) );
  INVX1 U51781 ( .A(mem_d_data_rd_i[19]), .Y(n73550) );
  NAND2X1 U51782 ( .A(n40935), .B(n73550), .Y(n49716) );
  INVX1 U51783 ( .A(n40360), .Y(n49718) );
  NAND2X1 U51784 ( .A(n37354), .B(n49718), .Y(n49721) );
  NAND2X1 U51785 ( .A(n2300), .B(n49719), .Y(n49720) );
  NAND2X1 U51786 ( .A(n49721), .B(n49720), .Y(n49722) );
  NAND2X1 U51787 ( .A(n42339), .B(n42344), .Y(n72815) );
  NAND2X1 U51788 ( .A(n43798), .B(n43772), .Y(n57852) );
  INVX1 U51789 ( .A(n57852), .Y(n49791) );
  NOR2X1 U51790 ( .A(n43454), .B(n43166), .Y(n49725) );
  NOR2X1 U51791 ( .A(n43021), .B(n43170), .Y(n49724) );
  NAND2X1 U51792 ( .A(n2314), .B(n43361), .Y(n49727) );
  NAND2X1 U51793 ( .A(n2289), .B(n38409), .Y(n49726) );
  NAND2X1 U51794 ( .A(n49727), .B(n49726), .Y(n49731) );
  NAND2X1 U51795 ( .A(n2296), .B(n38401), .Y(n49729) );
  NAND2X1 U51796 ( .A(n2304), .B(n38602), .Y(n49728) );
  NAND2X1 U51797 ( .A(n49729), .B(n49728), .Y(n49730) );
  NOR2X1 U51798 ( .A(n49731), .B(n49730), .Y(n49739) );
  NAND2X1 U51799 ( .A(n2286), .B(n38599), .Y(n49733) );
  NAND2X1 U51800 ( .A(n2292), .B(n43034), .Y(n49732) );
  NAND2X1 U51801 ( .A(n49733), .B(n49732), .Y(n49737) );
  NAND2X1 U51802 ( .A(n2306), .B(n38534), .Y(n49735) );
  NAND2X1 U51803 ( .A(n49735), .B(n49734), .Y(n49736) );
  NOR2X1 U51804 ( .A(n49737), .B(n49736), .Y(n49738) );
  NAND2X1 U51805 ( .A(n49739), .B(n49738), .Y(n49755) );
  NAND2X1 U51806 ( .A(n2302), .B(n43354), .Y(n49741) );
  NAND2X1 U51807 ( .A(n2300), .B(n40169), .Y(n49740) );
  NAND2X1 U51808 ( .A(n49741), .B(n49740), .Y(n49745) );
  NAND2X1 U51809 ( .A(n1834), .B(n39805), .Y(n49743) );
  NAND2X1 U51810 ( .A(n2308), .B(n43043), .Y(n49742) );
  NAND2X1 U51811 ( .A(n49743), .B(n49742), .Y(n49744) );
  NOR2X1 U51812 ( .A(n49745), .B(n49744), .Y(n49753) );
  NAND2X1 U51813 ( .A(n2312), .B(n38389), .Y(n49747) );
  NAND2X1 U51814 ( .A(n2287), .B(n43347), .Y(n49746) );
  NAND2X1 U51815 ( .A(n49747), .B(n49746), .Y(n49751) );
  NAND2X1 U51816 ( .A(n2294), .B(n43340), .Y(n49749) );
  NAND2X1 U51817 ( .A(n2310), .B(n43367), .Y(n49748) );
  NAND2X1 U51818 ( .A(n49749), .B(n49748), .Y(n49750) );
  NOR2X1 U51819 ( .A(n49751), .B(n49750), .Y(n49752) );
  NAND2X1 U51820 ( .A(n49753), .B(n49752), .Y(n49754) );
  NOR2X1 U51821 ( .A(n49755), .B(n49754), .Y(n49785) );
  NAND2X1 U51822 ( .A(n2307), .B(n40273), .Y(n49757) );
  NAND2X1 U51823 ( .A(n2313), .B(n43048), .Y(n49756) );
  NAND2X1 U51824 ( .A(n49757), .B(n49756), .Y(n49761) );
  NAND2X1 U51825 ( .A(n2305), .B(n43050), .Y(n49759) );
  NAND2X1 U51826 ( .A(n2290), .B(n43053), .Y(n49758) );
  NAND2X1 U51827 ( .A(n49759), .B(n49758), .Y(n49760) );
  NOR2X1 U51828 ( .A(n49761), .B(n49760), .Y(n49767) );
  NOR2X1 U51829 ( .A(n43371), .B(n36887), .Y(n49765) );
  NAND2X1 U51830 ( .A(n2293), .B(n38577), .Y(n49763) );
  NAND2X1 U51831 ( .A(n2315), .B(n40026), .Y(n49762) );
  NAND2X1 U51832 ( .A(n49763), .B(n49762), .Y(n49764) );
  NOR2X1 U51833 ( .A(n49765), .B(n49764), .Y(n49766) );
  NAND2X1 U51834 ( .A(n49767), .B(n49766), .Y(n49783) );
  NAND2X1 U51835 ( .A(n2311), .B(n43062), .Y(n49769) );
  NAND2X1 U51836 ( .A(n2309), .B(n39135), .Y(n49768) );
  NAND2X1 U51837 ( .A(n49769), .B(n49768), .Y(n49773) );
  NAND2X1 U51838 ( .A(n2301), .B(n40158), .Y(n49771) );
  NAND2X1 U51839 ( .A(n2291), .B(n38573), .Y(n49770) );
  NAND2X1 U51840 ( .A(n49771), .B(n49770), .Y(n49772) );
  NOR2X1 U51841 ( .A(n49773), .B(n49772), .Y(n49781) );
  NAND2X1 U51842 ( .A(n2303), .B(n43350), .Y(n49774) );
  NAND2X1 U51843 ( .A(n49775), .B(n49774), .Y(n49779) );
  NAND2X1 U51844 ( .A(n2295), .B(n43070), .Y(n49777) );
  NAND2X1 U51845 ( .A(n2288), .B(n43073), .Y(n49776) );
  NAND2X1 U51846 ( .A(n49777), .B(n49776), .Y(n49778) );
  NOR2X1 U51847 ( .A(n49779), .B(n49778), .Y(n49780) );
  NAND2X1 U51848 ( .A(n49781), .B(n49780), .Y(n49782) );
  NOR2X1 U51849 ( .A(n49783), .B(n49782), .Y(n49784) );
  NAND2X1 U51850 ( .A(n49785), .B(n49784), .Y(n49786) );
  NAND2X1 U51851 ( .A(n43923), .B(n43772), .Y(n49788) );
  NAND2X1 U51852 ( .A(n43915), .B(n43798), .Y(n49787) );
  NAND2X1 U51853 ( .A(n49788), .B(n49787), .Y(n57854) );
  INVX1 U51854 ( .A(n57854), .Y(n49789) );
  NAND2X1 U51855 ( .A(n43922), .B(n43915), .Y(n57851) );
  NAND2X1 U51856 ( .A(n49789), .B(n57851), .Y(n49790) );
  NOR2X1 U51857 ( .A(n49791), .B(n49790), .Y(n49792) );
  NOR2X1 U51858 ( .A(n49793), .B(n49792), .Y(n49794) );
  NAND2X1 U51859 ( .A(n43931), .B(n42658), .Y(n57863) );
  INVX1 U51860 ( .A(n57863), .Y(n57874) );
  NOR2X1 U51861 ( .A(n49794), .B(n57874), .Y(n49795) );
  NAND2X1 U51862 ( .A(n43922), .B(n43799), .Y(n57864) );
  NAND2X1 U51863 ( .A(n49795), .B(n57864), .Y(n49796) );
  NAND2X1 U51864 ( .A(n49797), .B(n49796), .Y(n49798) );
  NAND2X1 U51865 ( .A(n73436), .B(n49798), .Y(n49799) );
  NAND2X1 U51866 ( .A(n43988), .B(n43479), .Y(n57718) );
  NAND2X1 U51867 ( .A(n43978), .B(n43776), .Y(n49801) );
  NAND2X1 U51868 ( .A(n57718), .B(n49801), .Y(n31152) );
  NAND2X1 U51869 ( .A(n43490), .B(n43999), .Y(n57678) );
  NAND2X1 U51870 ( .A(n49804), .B(n57678), .Y(n49805) );
  NAND2X1 U51871 ( .A(n43495), .B(n49805), .Y(n49875) );
  NOR2X1 U51872 ( .A(n43454), .B(n43210), .Y(n49808) );
  NOR2X1 U51873 ( .A(n43021), .B(n43215), .Y(n49807) );
  NOR2X1 U51874 ( .A(n49808), .B(n49807), .Y(n49872) );
  NAND2X1 U51875 ( .A(n2814), .B(n43361), .Y(n49810) );
  NAND2X1 U51876 ( .A(n2789), .B(n38407), .Y(n49809) );
  NAND2X1 U51877 ( .A(n49810), .B(n49809), .Y(n49814) );
  NAND2X1 U51878 ( .A(n2796), .B(n43344), .Y(n49812) );
  NAND2X1 U51879 ( .A(n49812), .B(n49811), .Y(n49813) );
  NOR2X1 U51880 ( .A(n49814), .B(n49813), .Y(n49822) );
  NAND2X1 U51881 ( .A(n2786), .B(n38599), .Y(n49816) );
  NAND2X1 U51882 ( .A(n2791), .B(n43032), .Y(n49815) );
  NAND2X1 U51883 ( .A(n49816), .B(n49815), .Y(n49820) );
  NAND2X1 U51884 ( .A(n2806), .B(n38534), .Y(n49818) );
  NAND2X1 U51885 ( .A(n2798), .B(n43351), .Y(n49817) );
  NAND2X1 U51886 ( .A(n49818), .B(n49817), .Y(n49819) );
  NOR2X1 U51887 ( .A(n49820), .B(n49819), .Y(n49821) );
  NAND2X1 U51888 ( .A(n49822), .B(n49821), .Y(n49838) );
  NAND2X1 U51889 ( .A(n2802), .B(n43355), .Y(n49824) );
  NAND2X1 U51890 ( .A(n2800), .B(n40169), .Y(n49823) );
  NAND2X1 U51891 ( .A(n49824), .B(n49823), .Y(n49828) );
  NAND2X1 U51892 ( .A(n1811), .B(n39801), .Y(n49826) );
  NAND2X1 U51893 ( .A(n49826), .B(n49825), .Y(n49827) );
  NOR2X1 U51894 ( .A(n49828), .B(n49827), .Y(n49836) );
  NAND2X1 U51895 ( .A(n2812), .B(n43360), .Y(n49830) );
  NAND2X1 U51896 ( .A(n2787), .B(n43345), .Y(n49829) );
  NAND2X1 U51897 ( .A(n49830), .B(n49829), .Y(n49834) );
  NAND2X1 U51898 ( .A(n2794), .B(n43338), .Y(n49832) );
  NAND2X1 U51899 ( .A(n2810), .B(n43365), .Y(n49831) );
  NAND2X1 U51900 ( .A(n49832), .B(n49831), .Y(n49833) );
  NOR2X1 U51901 ( .A(n49834), .B(n49833), .Y(n49835) );
  NAND2X1 U51902 ( .A(n49836), .B(n49835), .Y(n49837) );
  NOR2X1 U51903 ( .A(n49838), .B(n49837), .Y(n49869) );
  NAND2X1 U51904 ( .A(n49840), .B(n49839), .Y(n49845) );
  NAND2X1 U51905 ( .A(n2790), .B(n43051), .Y(n49842) );
  NAND2X1 U51906 ( .A(n49843), .B(n49842), .Y(n49844) );
  NOR2X1 U51907 ( .A(n49845), .B(n49844), .Y(n49851) );
  NOR2X1 U51908 ( .A(n43371), .B(n37323), .Y(n49849) );
  NAND2X1 U51909 ( .A(n2792), .B(n38577), .Y(n49847) );
  NAND2X1 U51910 ( .A(n2815), .B(n40026), .Y(n49846) );
  NAND2X1 U51911 ( .A(n49847), .B(n49846), .Y(n49848) );
  NOR2X1 U51912 ( .A(n49849), .B(n49848), .Y(n49850) );
  NAND2X1 U51913 ( .A(n49851), .B(n49850), .Y(n49867) );
  NAND2X1 U51914 ( .A(n2811), .B(n43060), .Y(n49853) );
  NAND2X1 U51915 ( .A(n2809), .B(n39133), .Y(n49852) );
  NAND2X1 U51916 ( .A(n49853), .B(n49852), .Y(n49857) );
  NAND2X1 U51917 ( .A(n2801), .B(n43065), .Y(n49855) );
  NAND2X1 U51918 ( .A(n2793), .B(n38573), .Y(n49854) );
  NAND2X1 U51919 ( .A(n49855), .B(n49854), .Y(n49856) );
  NOR2X1 U51920 ( .A(n49857), .B(n49856), .Y(n49865) );
  NAND2X1 U51921 ( .A(n2797), .B(n43372), .Y(n49859) );
  NAND2X1 U51922 ( .A(n2803), .B(n43349), .Y(n49858) );
  NAND2X1 U51923 ( .A(n49859), .B(n49858), .Y(n49863) );
  NAND2X1 U51924 ( .A(n2795), .B(n43070), .Y(n49861) );
  NAND2X1 U51925 ( .A(n2788), .B(n43071), .Y(n49860) );
  NAND2X1 U51926 ( .A(n49861), .B(n49860), .Y(n49862) );
  NOR2X1 U51927 ( .A(n49863), .B(n49862), .Y(n49864) );
  NAND2X1 U51928 ( .A(n49865), .B(n49864), .Y(n49866) );
  NOR2X1 U51929 ( .A(n49867), .B(n49866), .Y(n49868) );
  NAND2X1 U51930 ( .A(n49869), .B(n49868), .Y(n49870) );
  NAND2X1 U51931 ( .A(n42805), .B(n49870), .Y(n49871) );
  NAND2X1 U51932 ( .A(n49872), .B(n49871), .Y(n73311) );
  NAND2X1 U51933 ( .A(n49873), .B(n44007), .Y(n49874) );
  NAND2X1 U51934 ( .A(n49875), .B(n49874), .Y(n49876) );
  NAND2X1 U51935 ( .A(n44021), .B(n43496), .Y(n57697) );
  NAND2X1 U51936 ( .A(n49876), .B(n57697), .Y(n49877) );
  NAND2X1 U51937 ( .A(n57695), .B(n49877), .Y(n49882) );
  NOR2X1 U51938 ( .A(n44024), .B(n49882), .Y(n49879) );
  NOR2X1 U51939 ( .A(n49879), .B(n49878), .Y(n49881) );
  NAND2X1 U51940 ( .A(n36706), .B(n44047), .Y(n49897) );
  NAND2X1 U51941 ( .A(n49897), .B(n58159), .Y(n49880) );
  NOR2X1 U51942 ( .A(n49881), .B(n49880), .Y(n49888) );
  INVX1 U51943 ( .A(n58159), .Y(n57676) );
  NOR2X1 U51944 ( .A(n57676), .B(n49882), .Y(n49884) );
  INVX1 U51945 ( .A(n49897), .Y(n57887) );
  NOR2X1 U51946 ( .A(n43504), .B(n57887), .Y(n49883) );
  NAND2X1 U51947 ( .A(n49884), .B(n49883), .Y(n49886) );
  NAND2X1 U51948 ( .A(n49886), .B(n49885), .Y(n49887) );
  NOR2X1 U51949 ( .A(n49890), .B(n49889), .Y(n49892) );
  INVX1 U51950 ( .A(n50040), .Y(n49891) );
  MX2X1 U51951 ( .A(n49892), .B(n49891), .S0(opcode_instr_w_24), .Y(n49893) );
  AND2X1 U51952 ( .A(n54897), .B(n49893), .Y(n50038) );
  NAND2X1 U51953 ( .A(n57676), .B(n49894), .Y(n49895) );
  NAND2X1 U51954 ( .A(n49897), .B(n49896), .Y(n49900) );
  NAND2X1 U51955 ( .A(n49898), .B(n50028), .Y(n49899) );
  NOR2X1 U51956 ( .A(n49900), .B(n49899), .Y(n50031) );
  NAND2X1 U51957 ( .A(n44634), .B(n39653), .Y(n49901) );
  NAND2X1 U51958 ( .A(n44833), .B(n40930), .Y(n50017) );
  NAND2X1 U51959 ( .A(n49901), .B(n42924), .Y(n50026) );
  NAND2X1 U51960 ( .A(n44634), .B(n39960), .Y(n49902) );
  XNOR2X1 U51961 ( .A(n44636), .B(n44053), .Y(n50251) );
  XNOR2X1 U51962 ( .A(n44638), .B(n44021), .Y(n50469) );
  XNOR2X1 U51963 ( .A(n44638), .B(n44013), .Y(n50115) );
  XNOR2X1 U51964 ( .A(n44637), .B(n43996), .Y(n50131) );
  XNOR2X1 U51965 ( .A(n44637), .B(n43989), .Y(n50411) );
  XNOR2X1 U51966 ( .A(n44637), .B(n43979), .Y(n50397) );
  XNOR2X1 U51967 ( .A(n44637), .B(n43949), .Y(n50268) );
  XNOR2X1 U51968 ( .A(n44637), .B(n43939), .Y(n50425) );
  XNOR2X1 U51969 ( .A(n44637), .B(n43932), .Y(n50168) );
  XNOR2X1 U51970 ( .A(n44636), .B(n43915), .Y(n50355) );
  XNOR2X1 U51971 ( .A(n44637), .B(n43902), .Y(n50151) );
  XNOR2X1 U51972 ( .A(n44637), .B(n43886), .Y(n50291) );
  XNOR2X1 U51973 ( .A(n44637), .B(n43876), .Y(n50375) );
  XNOR2X1 U51974 ( .A(n44637), .B(n43959), .Y(n50311) );
  XNOR2X1 U51975 ( .A(n44637), .B(n43969), .Y(n54971) );
  XNOR2X1 U51976 ( .A(n44637), .B(n43865), .Y(n54899) );
  XNOR2X1 U51977 ( .A(n44637), .B(n43856), .Y(n54781) );
  XNOR2X1 U51978 ( .A(n44637), .B(n44041), .Y(n54823) );
  XNOR2X1 U51979 ( .A(n44637), .B(n38385), .Y(n54721) );
  XNOR2X1 U51980 ( .A(n44637), .B(n43846), .Y(n54658) );
  XNOR2X1 U51981 ( .A(n44637), .B(n39945), .Y(n54598) );
  XNOR2X1 U51982 ( .A(n44637), .B(n43470), .Y(n54458) );
  XNOR2X1 U51983 ( .A(n44637), .B(n43475), .Y(n54514) );
  XNOR2X1 U51984 ( .A(n44636), .B(n40627), .Y(n54394) );
  NOR2X1 U51985 ( .A(n62458), .B(n39116), .Y(n49903) );
  NAND2X1 U51986 ( .A(n43734), .B(n73384), .Y(n57635) );
  MX2X1 U51987 ( .A(n49903), .B(n57635), .S0(n44636), .Y(n51926) );
  XNOR2X1 U51988 ( .A(n44636), .B(n38518), .Y(n51924) );
  INVX1 U51989 ( .A(n51924), .Y(n49905) );
  INVX1 U51990 ( .A(n51926), .Y(n49904) );
  NAND2X1 U51991 ( .A(n49905), .B(n49904), .Y(n49906) );
  MX2X1 U51992 ( .A(n40453), .B(n43753), .S0(n44635), .Y(n51923) );
  NAND2X1 U51993 ( .A(n54394), .B(n54395), .Y(n49910) );
  INVX1 U51994 ( .A(n54394), .Y(n49907) );
  NAND2X1 U51995 ( .A(n37939), .B(n49907), .Y(n49908) );
  MX2X1 U51996 ( .A(n36599), .B(n43814), .S0(n44636), .Y(n54393) );
  NAND2X1 U51997 ( .A(n49908), .B(n54393), .Y(n49909) );
  NAND2X1 U51998 ( .A(n49910), .B(n49909), .Y(n54516) );
  INVX1 U51999 ( .A(n54514), .Y(n49911) );
  NAND2X1 U52000 ( .A(n37942), .B(n49911), .Y(n49912) );
  MX2X1 U52001 ( .A(n42759), .B(n43805), .S0(n44636), .Y(n54513) );
  NAND2X1 U52002 ( .A(n54458), .B(n54460), .Y(n49917) );
  INVX1 U52003 ( .A(n54460), .Y(n49914) );
  INVX1 U52004 ( .A(n54458), .Y(n49913) );
  NAND2X1 U52005 ( .A(n49914), .B(n49913), .Y(n49915) );
  MX2X1 U52006 ( .A(n42747), .B(n43766), .S0(n44636), .Y(n54457) );
  NAND2X1 U52007 ( .A(n49915), .B(n54457), .Y(n49916) );
  NAND2X1 U52008 ( .A(n49917), .B(n49916), .Y(n54600) );
  NAND2X1 U52009 ( .A(n54598), .B(n54600), .Y(n49921) );
  INVX1 U52010 ( .A(n54598), .Y(n49918) );
  NAND2X1 U52011 ( .A(n37952), .B(n49918), .Y(n49919) );
  MX2X1 U52012 ( .A(opcode_opcode_w[25]), .B(n43744), .S0(n44636), .Y(n54597)
         );
  NAND2X1 U52013 ( .A(n49919), .B(n54597), .Y(n49920) );
  NAND2X1 U52014 ( .A(n49921), .B(n49920), .Y(n49922) );
  INVX1 U52015 ( .A(n49922), .Y(n54660) );
  INVX1 U52016 ( .A(n54658), .Y(n49923) );
  NAND2X1 U52017 ( .A(n54660), .B(n49923), .Y(n49924) );
  MX2X1 U52018 ( .A(opcode_opcode_w[26]), .B(n43792), .S0(n44636), .Y(n54657)
         );
  NAND2X1 U52019 ( .A(n54721), .B(n49925), .Y(n49929) );
  INVX1 U52020 ( .A(n54721), .Y(n49926) );
  NAND2X1 U52021 ( .A(n37893), .B(n49926), .Y(n49927) );
  MX2X1 U52022 ( .A(opcode_opcode_w[27]), .B(n43780), .S0(n44636), .Y(n54720)
         );
  NAND2X1 U52023 ( .A(n49927), .B(n54720), .Y(n49928) );
  NAND2X1 U52024 ( .A(n49929), .B(n49928), .Y(n49930) );
  INVX1 U52025 ( .A(n49930), .Y(n54825) );
  INVX1 U52026 ( .A(n54823), .Y(n49931) );
  NAND2X1 U52027 ( .A(n54825), .B(n49931), .Y(n49932) );
  MX2X1 U52028 ( .A(opcode_opcode_w[28]), .B(n43738), .S0(n44636), .Y(n54822)
         );
  NAND2X1 U52029 ( .A(n54781), .B(n49933), .Y(n49937) );
  INVX1 U52030 ( .A(n54781), .Y(n49934) );
  NAND2X1 U52031 ( .A(n37898), .B(n49934), .Y(n49935) );
  MX2X1 U52032 ( .A(opcode_opcode_w[29]), .B(n43758), .S0(n44636), .Y(n54780)
         );
  NAND2X1 U52033 ( .A(n49935), .B(n54780), .Y(n49936) );
  NAND2X1 U52034 ( .A(n49937), .B(n49936), .Y(n49938) );
  INVX1 U52035 ( .A(n49938), .Y(n54901) );
  INVX1 U52036 ( .A(n54899), .Y(n49939) );
  NAND2X1 U52037 ( .A(n54901), .B(n49939), .Y(n49940) );
  MX2X1 U52038 ( .A(opcode_opcode_w[30]), .B(n43821), .S0(n44635), .Y(n54898)
         );
  INVX1 U52039 ( .A(n54972), .Y(n49942) );
  INVX1 U52040 ( .A(n54971), .Y(n49941) );
  NAND2X1 U52041 ( .A(n49942), .B(n49941), .Y(n49944) );
  NAND2X1 U52042 ( .A(n44635), .B(n43812), .Y(n49943) );
  NAND2X1 U52043 ( .A(n49943), .B(n42925), .Y(n54970) );
  INVX1 U52044 ( .A(n50311), .Y(n49945) );
  NAND2X1 U52045 ( .A(n37984), .B(n49945), .Y(n49947) );
  NAND2X1 U52046 ( .A(n44635), .B(n40466), .Y(n49946) );
  NAND2X1 U52047 ( .A(n49946), .B(n42926), .Y(n50310) );
  INVX1 U52048 ( .A(n50377), .Y(n49949) );
  INVX1 U52049 ( .A(n50375), .Y(n49948) );
  NAND2X1 U52050 ( .A(n49949), .B(n49948), .Y(n49951) );
  NAND2X1 U52051 ( .A(n44635), .B(n40472), .Y(n49950) );
  NAND2X1 U52052 ( .A(n49950), .B(n42927), .Y(n50374) );
  INVX1 U52053 ( .A(n50293), .Y(n49953) );
  INVX1 U52054 ( .A(n50291), .Y(n49952) );
  NAND2X1 U52055 ( .A(n49953), .B(n49952), .Y(n49955) );
  NAND2X1 U52056 ( .A(n44635), .B(n40487), .Y(n49954) );
  NAND2X1 U52057 ( .A(n49954), .B(n42923), .Y(n50290) );
  INVX1 U52058 ( .A(n50328), .Y(n49956) );
  NAND2X1 U52059 ( .A(n37989), .B(n49956), .Y(n49958) );
  NAND2X1 U52060 ( .A(n44634), .B(n43787), .Y(n49957) );
  NAND2X1 U52061 ( .A(n49957), .B(n42928), .Y(n50327) );
  NAND2X1 U52062 ( .A(n50151), .B(n50152), .Y(n49964) );
  INVX1 U52063 ( .A(n50152), .Y(n49960) );
  INVX1 U52064 ( .A(n50151), .Y(n49959) );
  NAND2X1 U52065 ( .A(n49960), .B(n49959), .Y(n49962) );
  NAND2X1 U52066 ( .A(n44635), .B(n43724), .Y(n49961) );
  NAND2X1 U52067 ( .A(n49961), .B(n42922), .Y(n50150) );
  NAND2X1 U52068 ( .A(n49962), .B(n50150), .Y(n49963) );
  NAND2X1 U52069 ( .A(n49964), .B(n49963), .Y(n49965) );
  INVX1 U52070 ( .A(n49965), .Y(n50080) );
  INVX1 U52071 ( .A(n49966), .Y(n50079) );
  NAND2X1 U52072 ( .A(n50080), .B(n50079), .Y(n49968) );
  NAND2X1 U52073 ( .A(n44635), .B(n42636), .Y(n49967) );
  NAND2X1 U52074 ( .A(n49967), .B(n42923), .Y(n50078) );
  INVX1 U52075 ( .A(n50355), .Y(n49969) );
  NAND2X1 U52076 ( .A(n37959), .B(n49969), .Y(n49971) );
  NAND2X1 U52077 ( .A(n44635), .B(n40259), .Y(n49970) );
  NAND2X1 U52078 ( .A(n49970), .B(n42928), .Y(n50354) );
  INVX1 U52079 ( .A(n50451), .Y(n49973) );
  INVX1 U52080 ( .A(n50449), .Y(n49972) );
  NAND2X1 U52081 ( .A(n49973), .B(n49972), .Y(n49975) );
  NAND2X1 U52082 ( .A(n44634), .B(n43798), .Y(n49974) );
  NAND2X1 U52083 ( .A(n49974), .B(n42922), .Y(n50448) );
  NAND2X1 U52084 ( .A(n50168), .B(n50169), .Y(n49980) );
  INVX1 U52085 ( .A(n50168), .Y(n49976) );
  NAND2X1 U52086 ( .A(n37995), .B(n49976), .Y(n49978) );
  NAND2X1 U52087 ( .A(n44635), .B(n42652), .Y(n49977) );
  NAND2X1 U52088 ( .A(n49977), .B(n42923), .Y(n50167) );
  NAND2X1 U52089 ( .A(n49978), .B(n50167), .Y(n49979) );
  NAND2X1 U52090 ( .A(n49980), .B(n49979), .Y(n49981) );
  INVX1 U52091 ( .A(n49981), .Y(n50427) );
  INVX1 U52092 ( .A(n50425), .Y(n49982) );
  NAND2X1 U52093 ( .A(n50427), .B(n49982), .Y(n49984) );
  NAND2X1 U52094 ( .A(n44634), .B(n42712), .Y(n49983) );
  NAND2X1 U52095 ( .A(n49983), .B(n42924), .Y(n50424) );
  NAND2X1 U52096 ( .A(n50268), .B(n49985), .Y(n49990) );
  INVX1 U52097 ( .A(n50268), .Y(n49986) );
  NAND2X1 U52098 ( .A(n44634), .B(n43795), .Y(n49987) );
  NAND2X1 U52099 ( .A(n49987), .B(n42924), .Y(n50267) );
  NAND2X1 U52100 ( .A(n49988), .B(n50267), .Y(n49989) );
  NAND2X1 U52101 ( .A(n49990), .B(n49989), .Y(n49991) );
  INVX1 U52102 ( .A(n49991), .Y(n50399) );
  INVX1 U52103 ( .A(n50397), .Y(n49992) );
  NAND2X1 U52104 ( .A(n50399), .B(n49992), .Y(n49994) );
  NAND2X1 U52105 ( .A(n44634), .B(n43776), .Y(n49993) );
  NAND2X1 U52106 ( .A(n49993), .B(n42924), .Y(n50396) );
  INVX1 U52107 ( .A(n49995), .Y(n50413) );
  INVX1 U52108 ( .A(n50411), .Y(n49996) );
  NAND2X1 U52109 ( .A(n50413), .B(n49996), .Y(n49998) );
  NAND2X1 U52110 ( .A(n44634), .B(n43479), .Y(n49997) );
  NAND2X1 U52111 ( .A(n49997), .B(n42924), .Y(n50410) );
  INVX1 U52112 ( .A(n49999), .Y(n50133) );
  INVX1 U52113 ( .A(n50131), .Y(n50000) );
  NAND2X1 U52114 ( .A(n50133), .B(n50000), .Y(n50002) );
  NAND2X1 U52115 ( .A(n44634), .B(n38312), .Y(n50001) );
  NAND2X1 U52116 ( .A(n50001), .B(n42925), .Y(n50130) );
  INVX1 U52117 ( .A(n50003), .Y(n50215) );
  INVX1 U52118 ( .A(n50213), .Y(n50004) );
  NAND2X1 U52119 ( .A(n50215), .B(n50004), .Y(n50006) );
  NAND2X1 U52120 ( .A(n44634), .B(n43487), .Y(n50005) );
  NAND2X1 U52121 ( .A(n50005), .B(n42924), .Y(n50212) );
  INVX1 U52122 ( .A(n50117), .Y(n50008) );
  INVX1 U52123 ( .A(n50115), .Y(n50007) );
  NAND2X1 U52124 ( .A(n50008), .B(n50007), .Y(n50010) );
  NAND2X1 U52125 ( .A(n44634), .B(n43493), .Y(n50009) );
  NAND2X1 U52126 ( .A(n50009), .B(n42925), .Y(n50114) );
  INVX1 U52127 ( .A(n50471), .Y(n50012) );
  INVX1 U52128 ( .A(n50469), .Y(n50011) );
  NAND2X1 U52129 ( .A(n50012), .B(n50011), .Y(n50014) );
  NAND2X1 U52130 ( .A(n44634), .B(n43497), .Y(n50013) );
  NAND2X1 U52131 ( .A(n50013), .B(n42926), .Y(n50468) );
  INVX1 U52132 ( .A(n50199), .Y(n50016) );
  INVX1 U52133 ( .A(n50197), .Y(n50015) );
  NAND2X1 U52134 ( .A(n50016), .B(n50015), .Y(n50019) );
  NAND2X1 U52135 ( .A(n44635), .B(n43502), .Y(n50018) );
  NAND2X1 U52136 ( .A(n50018), .B(n42927), .Y(n50196) );
  NOR2X1 U52137 ( .A(n50251), .B(n50253), .Y(n50020) );
  NOR2X1 U52138 ( .A(n42298), .B(n50020), .Y(n50024) );
  INVX1 U52139 ( .A(n50253), .Y(n50022) );
  INVX1 U52140 ( .A(n50251), .Y(n50021) );
  NOR2X1 U52141 ( .A(n50022), .B(n50021), .Y(n50023) );
  NOR2X1 U52142 ( .A(n50024), .B(n50023), .Y(n50025) );
  XNOR2X1 U52143 ( .A(n50026), .B(n50025), .Y(n50027) );
  INVX1 U52144 ( .A(n50229), .Y(n50029) );
  NAND2X1 U52145 ( .A(opcode_instr_w_26), .B(n50028), .Y(n50034) );
  NOR2X1 U52146 ( .A(n50029), .B(n50034), .Y(n50030) );
  NOR2X1 U52147 ( .A(n50031), .B(n50030), .Y(n50032) );
  NOR2X1 U52148 ( .A(opcode_instr_w_24), .B(n50034), .Y(n50035) );
  NOR2X1 U52149 ( .A(n1888), .B(n50035), .Y(n50036) );
  NOR2X1 U52150 ( .A(n42873), .B(n50039), .Y(n50041) );
  NAND2X1 U52151 ( .A(n8696), .B(n50042), .Y(n54382) );
  NAND2X1 U52152 ( .A(n50044), .B(n37413), .Y(n8443) );
  INVX1 U52153 ( .A(rst_i), .Y(n73547) );
  INVX1 U52154 ( .A(mem_i_inst_i[19]), .Y(n50054) );
  NOR2X1 U52155 ( .A(n50045), .B(n57427), .Y(n50049) );
  INVX1 U52156 ( .A(n28934), .Y(n50047) );
  NOR2X1 U52157 ( .A(n50047), .B(n50046), .Y(n50048) );
  NAND2X1 U52158 ( .A(n50049), .B(n50048), .Y(n50499) );
  NAND2X1 U52159 ( .A(n8696), .B(n50499), .Y(n73387) );
  INVX1 U52160 ( .A(n73387), .Y(n50052) );
  NOR2X1 U52161 ( .A(mem_i_valid_i), .B(n58511), .Y(n50050) );
  NAND2X1 U52162 ( .A(n50050), .B(n50534), .Y(n50051) );
  NAND2X1 U52163 ( .A(n38002), .B(n50051), .Y(n57559) );
  INVX1 U52164 ( .A(n57559), .Y(n73390) );
  NAND2X1 U52165 ( .A(n50052), .B(n73390), .Y(n57280) );
  INVX1 U52166 ( .A(mem_i_error_i), .Y(n50053) );
  NAND2X1 U52167 ( .A(n50534), .B(n50053), .Y(n58506) );
  INVX1 U52168 ( .A(n58506), .Y(n50496) );
  NOR2X1 U52169 ( .A(n50054), .B(n43404), .Y(net2361) );
  NAND2X1 U52170 ( .A(n43319), .B(n58511), .Y(n50055) );
  NAND2X1 U52171 ( .A(n50055), .B(n44858), .Y(n54437) );
  NAND2X1 U52172 ( .A(challenge[105]), .B(n44848), .Y(n50056) );
  NAND2X1 U52173 ( .A(n54437), .B(n50056), .Y(n17313) );
  NAND2X1 U52174 ( .A(n29680), .B(u_mmu_itlb_entry_q_3), .Y(n50057) );
  NAND2X1 U52175 ( .A(n44073), .B(n50057), .Y(n58126) );
  NOR2X1 U52176 ( .A(n2162), .B(n43305), .Y(n50110) );
  NAND2X1 U52177 ( .A(n43307), .B(n55361), .Y(n50109) );
  XNOR2X1 U52178 ( .A(opcode_pc_w[17]), .B(n42851), .Y(n50076) );
  NAND2X1 U52179 ( .A(opcode_pc_w[16]), .B(n44836), .Y(n50075) );
  NAND2X1 U52180 ( .A(n44841), .B(n58319), .Y(n50073) );
  NAND2X1 U52181 ( .A(opcode_pc_w[15]), .B(n44836), .Y(n50072) );
  NAND2X1 U52182 ( .A(n44842), .B(n58312), .Y(n50070) );
  NAND2X1 U52183 ( .A(opcode_pc_w[14]), .B(n44836), .Y(n50069) );
  NAND2X1 U52184 ( .A(n44844), .B(n58305), .Y(n50067) );
  NAND2X1 U52185 ( .A(opcode_pc_w[13]), .B(n44836), .Y(n50066) );
  NAND2X1 U52186 ( .A(n44839), .B(n58298), .Y(n50064) );
  NAND2X1 U52187 ( .A(opcode_pc_w[12]), .B(n44836), .Y(n50063) );
  NAND2X1 U52188 ( .A(n44839), .B(n58291), .Y(n50061) );
  NAND2X1 U52189 ( .A(opcode_pc_w[11]), .B(opcode_opcode_w[7]), .Y(n50060) );
  NAND2X1 U52190 ( .A(n50700), .B(n58286), .Y(n50058) );
  NAND2X1 U52191 ( .A(opcode_pc_w[10]), .B(opcode_opcode_w[30]), .Y(n29942) );
  NAND2X1 U52192 ( .A(n30771), .B(n29942), .Y(n54968) );
  NAND2X1 U52193 ( .A(n50058), .B(n54968), .Y(n50059) );
  NAND2X1 U52194 ( .A(n50060), .B(n50059), .Y(n50308) );
  NAND2X1 U52195 ( .A(n50061), .B(n50308), .Y(n50062) );
  NAND2X1 U52196 ( .A(n50063), .B(n50062), .Y(n50372) );
  NAND2X1 U52197 ( .A(n50064), .B(n50372), .Y(n50065) );
  NAND2X1 U52198 ( .A(n50066), .B(n50065), .Y(n50288) );
  NAND2X1 U52199 ( .A(n50067), .B(n50288), .Y(n50068) );
  NAND2X1 U52200 ( .A(n50069), .B(n50068), .Y(n50325) );
  NAND2X1 U52201 ( .A(n50070), .B(n50325), .Y(n50071) );
  NAND2X1 U52202 ( .A(n50072), .B(n50071), .Y(n50148) );
  NAND2X1 U52203 ( .A(n50073), .B(n50148), .Y(n50074) );
  NAND2X1 U52204 ( .A(n50075), .B(n50074), .Y(n50349) );
  NOR2X1 U52205 ( .A(n50077), .B(n42874), .Y(n50084) );
  XNOR2X1 U52206 ( .A(n50081), .B(n50080), .Y(n50082) );
  NOR2X1 U52207 ( .A(n50082), .B(n42929), .Y(n50083) );
  NOR2X1 U52208 ( .A(n50084), .B(n50083), .Y(n50107) );
  NAND2X1 U52209 ( .A(opcode_pc_w[16]), .B(n42722), .Y(n50102) );
  NAND2X1 U52210 ( .A(n42725), .B(n58319), .Y(n50100) );
  NAND2X1 U52211 ( .A(opcode_pc_w[15]), .B(n42728), .Y(n50099) );
  NAND2X1 U52212 ( .A(n42730), .B(n58312), .Y(n50097) );
  NAND2X1 U52213 ( .A(opcode_opcode_w[14]), .B(opcode_pc_w[14]), .Y(n50096) );
  NAND2X1 U52214 ( .A(n58305), .B(n56876), .Y(n50094) );
  NAND2X1 U52215 ( .A(opcode_opcode_w[13]), .B(opcode_pc_w[13]), .Y(n50093) );
  NAND2X1 U52216 ( .A(n58298), .B(n56868), .Y(n50091) );
  NAND2X1 U52217 ( .A(opcode_opcode_w[12]), .B(opcode_pc_w[12]), .Y(n50090) );
  NAND2X1 U52218 ( .A(n58291), .B(n56860), .Y(n50088) );
  NAND2X1 U52219 ( .A(opcode_pc_w[11]), .B(n39115), .Y(n50087) );
  NAND2X1 U52220 ( .A(n39116), .B(n58286), .Y(n50085) );
  NAND2X1 U52221 ( .A(n30820), .B(n29942), .Y(n54976) );
  NAND2X1 U52222 ( .A(n50085), .B(n54976), .Y(n50086) );
  NAND2X1 U52223 ( .A(n50087), .B(n50086), .Y(n50316) );
  NAND2X1 U52224 ( .A(n50088), .B(n50316), .Y(n50089) );
  NAND2X1 U52225 ( .A(n50090), .B(n50089), .Y(n50381) );
  NAND2X1 U52226 ( .A(n50091), .B(n50381), .Y(n50092) );
  NAND2X1 U52227 ( .A(n50093), .B(n50092), .Y(n50297) );
  NAND2X1 U52228 ( .A(n50094), .B(n50297), .Y(n50095) );
  NAND2X1 U52229 ( .A(n50096), .B(n50095), .Y(n50334) );
  NAND2X1 U52230 ( .A(n50097), .B(n50334), .Y(n50098) );
  NAND2X1 U52231 ( .A(n50099), .B(n50098), .Y(n50156) );
  NAND2X1 U52232 ( .A(n50100), .B(n50156), .Y(n50101) );
  NAND2X1 U52233 ( .A(n50102), .B(n50101), .Y(n50171) );
  INVX1 U52234 ( .A(n50171), .Y(n50104) );
  XNOR2X1 U52235 ( .A(n42688), .B(opcode_pc_w[17]), .Y(n50103) );
  XNOR2X1 U52236 ( .A(n50104), .B(n50103), .Y(n50105) );
  INVX1 U52237 ( .A(n43013), .Y(n54979) );
  NAND2X1 U52238 ( .A(n50105), .B(n54979), .Y(n50106) );
  NAND2X1 U52239 ( .A(n50107), .B(n50106), .Y(n55360) );
  NAND2X1 U52240 ( .A(n43313), .B(n55360), .Y(n50108) );
  NAND2X1 U52241 ( .A(n50109), .B(n50108), .Y(n55365) );
  NOR2X1 U52242 ( .A(n50110), .B(n55365), .Y(n50112) );
  OR2X1 U52243 ( .A(n1775), .B(n42846), .Y(n50111) );
  NAND2X1 U52244 ( .A(n50112), .B(n50111), .Y(n6) );
  INVX1 U52245 ( .A(n6), .Y(n55416) );
  XNOR2X1 U52246 ( .A(n2883), .B(n55416), .Y(n50147) );
  NOR2X1 U52247 ( .A(n1938), .B(n43305), .Y(n50127) );
  NAND2X1 U52248 ( .A(n43309), .B(n55989), .Y(n50126) );
  NAND2X1 U52249 ( .A(n44839), .B(n58389), .Y(n30414) );
  NAND2X1 U52250 ( .A(opcode_pc_w[27]), .B(n44836), .Y(n50475) );
  NAND2X1 U52251 ( .A(n30414), .B(n50475), .Y(n50121) );
  NAND2X1 U52252 ( .A(opcode_pc_w[26]), .B(n44836), .Y(n30546) );
  NAND2X1 U52253 ( .A(n30547), .B(n30546), .Y(n30403) );
  XOR2X1 U52254 ( .A(n50121), .B(n30403), .Y(n50113) );
  NOR2X1 U52255 ( .A(n50113), .B(n42872), .Y(n50120) );
  XNOR2X1 U52256 ( .A(n50115), .B(n50114), .Y(n50116) );
  XOR2X1 U52257 ( .A(n50117), .B(n50116), .Y(n50118) );
  NOR2X1 U52258 ( .A(n50118), .B(n42929), .Y(n50119) );
  NOR2X1 U52259 ( .A(n50120), .B(n50119), .Y(n50124) );
  NAND2X1 U52260 ( .A(n30560), .B(n30546), .Y(n30413) );
  XNOR2X1 U52261 ( .A(n50121), .B(n30413), .Y(n50122) );
  NAND2X1 U52262 ( .A(n50122), .B(n54979), .Y(n50123) );
  NAND2X1 U52263 ( .A(n50124), .B(n50123), .Y(n55988) );
  NAND2X1 U52264 ( .A(n43311), .B(n55988), .Y(n50125) );
  NAND2X1 U52265 ( .A(n50126), .B(n50125), .Y(n55995) );
  NOR2X1 U52266 ( .A(n50127), .B(n55995), .Y(n50129) );
  OR2X1 U52267 ( .A(n1785), .B(n43314), .Y(n50128) );
  NAND2X1 U52268 ( .A(n50129), .B(n50128), .Y(n19) );
  XNOR2X1 U52269 ( .A(n19), .B(u_mmu_itlb_va_addr_q[27]), .Y(n50145) );
  NOR2X1 U52270 ( .A(n2186), .B(n43305), .Y(n50141) );
  NAND2X1 U52271 ( .A(n43309), .B(n55766), .Y(n50140) );
  NOR2X1 U52272 ( .A(n30327), .B(n37342), .Y(n50138) );
  NAND2X1 U52273 ( .A(n30317), .B(n54897), .Y(n50136) );
  INVX1 U52274 ( .A(n42929), .Y(n54903) );
  XNOR2X1 U52275 ( .A(n50133), .B(n50132), .Y(n50134) );
  NAND2X1 U52276 ( .A(n54903), .B(n50134), .Y(n50135) );
  NAND2X1 U52277 ( .A(n50136), .B(n50135), .Y(n50137) );
  OR2X1 U52278 ( .A(n50138), .B(n50137), .Y(n55765) );
  NAND2X1 U52279 ( .A(n43311), .B(n55765), .Y(n50139) );
  NAND2X1 U52280 ( .A(n50140), .B(n50139), .Y(n55770) );
  NOR2X1 U52281 ( .A(n50141), .B(n55770), .Y(n50143) );
  OR2X1 U52282 ( .A(n1783), .B(n43314), .Y(n50142) );
  NAND2X1 U52283 ( .A(n50143), .B(n50142), .Y(n23) );
  XNOR2X1 U52284 ( .A(n23), .B(u_mmu_itlb_va_addr_q[25]), .Y(n50144) );
  NAND2X1 U52285 ( .A(n50145), .B(n50144), .Y(n50146) );
  NOR2X1 U52286 ( .A(n50147), .B(n50146), .Y(n50194) );
  NOR2X1 U52287 ( .A(n2159), .B(n43305), .Y(n50164) );
  NAND2X1 U52288 ( .A(n43309), .B(n55301), .Y(n50163) );
  NOR2X1 U52289 ( .A(n50149), .B(n42873), .Y(n50155) );
  NOR2X1 U52290 ( .A(n50153), .B(n42929), .Y(n50154) );
  NOR2X1 U52291 ( .A(n50155), .B(n50154), .Y(n50161) );
  INVX1 U52292 ( .A(n50156), .Y(n50158) );
  XNOR2X1 U52293 ( .A(n42722), .B(opcode_pc_w[16]), .Y(n50157) );
  XOR2X1 U52294 ( .A(n50158), .B(n50157), .Y(n50159) );
  NAND2X1 U52295 ( .A(n50159), .B(n54979), .Y(n50160) );
  NAND2X1 U52296 ( .A(n50161), .B(n50160), .Y(n55300) );
  NAND2X1 U52297 ( .A(n43311), .B(n55300), .Y(n50162) );
  NAND2X1 U52298 ( .A(n50163), .B(n50162), .Y(n55314) );
  NOR2X1 U52299 ( .A(n50164), .B(n55314), .Y(n50166) );
  OR2X1 U52300 ( .A(n1774), .B(n43314), .Y(n50165) );
  NAND2X1 U52301 ( .A(n50166), .B(n50165), .Y(n8) );
  INVX1 U52302 ( .A(n8), .Y(n55305) );
  XNOR2X1 U52303 ( .A(n2517), .B(n55305), .Y(n50192) );
  NOR2X1 U52304 ( .A(n2171), .B(n43305), .Y(n50188) );
  NAND2X1 U52305 ( .A(n43309), .B(n55519), .Y(n50187) );
  NOR2X1 U52306 ( .A(n50170), .B(n42929), .Y(n50183) );
  NAND2X1 U52307 ( .A(opcode_pc_w[19]), .B(n42792), .Y(n50180) );
  NAND2X1 U52308 ( .A(n42790), .B(n58338), .Y(n50178) );
  NAND2X1 U52309 ( .A(opcode_pc_w[18]), .B(opcode_opcode_w[18]), .Y(n50177) );
  NAND2X1 U52310 ( .A(n42662), .B(n58331), .Y(n50175) );
  NAND2X1 U52311 ( .A(opcode_pc_w[17]), .B(n42686), .Y(n50174) );
  NAND2X1 U52312 ( .A(n42688), .B(n58324), .Y(n50172) );
  NAND2X1 U52313 ( .A(n50172), .B(n50171), .Y(n50173) );
  NAND2X1 U52314 ( .A(n50174), .B(n50173), .Y(n50361) );
  NAND2X1 U52315 ( .A(n50175), .B(n50361), .Y(n50176) );
  NAND2X1 U52316 ( .A(n50177), .B(n50176), .Y(n50455) );
  NAND2X1 U52317 ( .A(n50178), .B(n50455), .Y(n50179) );
  NAND2X1 U52318 ( .A(n50180), .B(n50179), .Y(n30637) );
  XOR2X1 U52319 ( .A(n30709), .B(n30637), .Y(n50181) );
  NOR2X1 U52320 ( .A(n43013), .B(n50181), .Y(n50182) );
  NOR2X1 U52321 ( .A(n50183), .B(n50182), .Y(n50185) );
  NAND2X1 U52322 ( .A(n30708), .B(n54897), .Y(n50184) );
  NAND2X1 U52323 ( .A(n50185), .B(n50184), .Y(n55518) );
  NAND2X1 U52324 ( .A(n43313), .B(n55518), .Y(n50186) );
  NAND2X1 U52325 ( .A(n50187), .B(n50186), .Y(n55524) );
  NOR2X1 U52326 ( .A(n50188), .B(n55524), .Y(n50190) );
  OR2X1 U52327 ( .A(n1778), .B(n43314), .Y(n50189) );
  NAND2X1 U52328 ( .A(n50190), .B(n50189), .Y(n7) );
  INVX1 U52329 ( .A(n7), .Y(n55522) );
  XNOR2X1 U52330 ( .A(n2384), .B(n55522), .Y(n50191) );
  NOR2X1 U52331 ( .A(n50192), .B(n50191), .Y(n50193) );
  NAND2X1 U52332 ( .A(n50194), .B(n50193), .Y(n50287) );
  NOR2X1 U52333 ( .A(n1934), .B(n43306), .Y(n50209) );
  NAND2X1 U52334 ( .A(n43309), .B(n56349), .Y(n50208) );
  NAND2X1 U52335 ( .A(n44840), .B(n58403), .Y(n30494) );
  NAND2X1 U52336 ( .A(opcode_pc_w[29]), .B(n44835), .Y(n50257) );
  NAND2X1 U52337 ( .A(n30494), .B(n50257), .Y(n50203) );
  NAND2X1 U52338 ( .A(opcode_pc_w[28]), .B(n44835), .Y(n50466) );
  NAND2X1 U52339 ( .A(n30544), .B(n50466), .Y(n30495) );
  XOR2X1 U52340 ( .A(n50203), .B(n30495), .Y(n50195) );
  NOR2X1 U52341 ( .A(n50195), .B(n42874), .Y(n50202) );
  XNOR2X1 U52342 ( .A(n50197), .B(n50196), .Y(n50198) );
  XOR2X1 U52343 ( .A(n50199), .B(n50198), .Y(n50200) );
  NOR2X1 U52344 ( .A(n50200), .B(n42931), .Y(n50201) );
  NOR2X1 U52345 ( .A(n50202), .B(n50201), .Y(n50206) );
  NAND2X1 U52346 ( .A(n30558), .B(n50466), .Y(n30505) );
  XNOR2X1 U52347 ( .A(n50203), .B(n30505), .Y(n50204) );
  NAND2X1 U52348 ( .A(n50204), .B(n54979), .Y(n50205) );
  NAND2X1 U52349 ( .A(n50206), .B(n50205), .Y(n56348) );
  NAND2X1 U52350 ( .A(n43313), .B(n56348), .Y(n50207) );
  NAND2X1 U52351 ( .A(n50208), .B(n50207), .Y(n56181) );
  NOR2X1 U52352 ( .A(n50209), .B(n56181), .Y(n50211) );
  OR2X1 U52353 ( .A(n1787), .B(n43314), .Y(n50210) );
  NAND2X1 U52354 ( .A(n50211), .B(n50210), .Y(n14) );
  INVX1 U52355 ( .A(n14), .Y(n56352) );
  XNOR2X1 U52356 ( .A(u_mmu_itlb_va_addr_q[29]), .B(n56352), .Y(n50228) );
  NOR2X1 U52357 ( .A(n2189), .B(n43306), .Y(n50223) );
  NAND2X1 U52358 ( .A(n43309), .B(n55812), .Y(n50222) );
  NOR2X1 U52359 ( .A(n30583), .B(n43014), .Y(n50220) );
  NAND2X1 U52360 ( .A(n30569), .B(n54897), .Y(n50218) );
  XNOR2X1 U52361 ( .A(n50215), .B(n50214), .Y(n50216) );
  NAND2X1 U52362 ( .A(n54903), .B(n50216), .Y(n50217) );
  NAND2X1 U52363 ( .A(n50218), .B(n50217), .Y(n50219) );
  OR2X1 U52364 ( .A(n50220), .B(n50219), .Y(n55811) );
  NAND2X1 U52365 ( .A(n43313), .B(n55811), .Y(n50221) );
  NAND2X1 U52366 ( .A(n50222), .B(n50221), .Y(n54370) );
  NOR2X1 U52367 ( .A(n50223), .B(n54370), .Y(n50225) );
  OR2X1 U52368 ( .A(n1784), .B(n43314), .Y(n50224) );
  NAND2X1 U52369 ( .A(n50225), .B(n50224), .Y(n13) );
  XNOR2X1 U52370 ( .A(n13), .B(u_mmu_itlb_va_addr_q[26]), .Y(n50226) );
  NAND2X1 U52371 ( .A(u_mmu_itlb_valid_q), .B(n50226), .Y(n50227) );
  NOR2X1 U52372 ( .A(n50228), .B(n50227), .Y(n50285) );
  NOR2X1 U52373 ( .A(n2916), .B(n43306), .Y(n50246) );
  NAND2X1 U52374 ( .A(n43308), .B(n56613), .Y(n50245) );
  NAND2X1 U52375 ( .A(n54903), .B(n50229), .Y(n50243) );
  NAND2X1 U52376 ( .A(opcode_pc_w[30]), .B(n44836), .Y(n50249) );
  INVX1 U52377 ( .A(n50249), .Y(n50231) );
  OR2X1 U52378 ( .A(n30426), .B(n50231), .Y(n50235) );
  INVX1 U52379 ( .A(n50235), .Y(n50230) );
  NOR2X1 U52380 ( .A(n50230), .B(n42872), .Y(n50234) );
  OR2X1 U52381 ( .A(n30435), .B(n50231), .Y(n50236) );
  INVX1 U52382 ( .A(n50236), .Y(n50232) );
  NOR2X1 U52383 ( .A(n43013), .B(n50232), .Y(n50233) );
  NOR2X1 U52384 ( .A(n50234), .B(n50233), .Y(n50241) );
  NOR2X1 U52385 ( .A(n42874), .B(n50235), .Y(n50238) );
  NOR2X1 U52386 ( .A(n43014), .B(n50236), .Y(n50237) );
  NOR2X1 U52387 ( .A(n50238), .B(n50237), .Y(n50240) );
  XNOR2X1 U52388 ( .A(n44845), .B(opcode_pc_w[31]), .Y(n50239) );
  MX2X1 U52389 ( .A(n50241), .B(n50240), .S0(n50239), .Y(n50242) );
  NAND2X1 U52390 ( .A(n50243), .B(n50242), .Y(n56612) );
  NAND2X1 U52391 ( .A(n43313), .B(n56612), .Y(n50244) );
  NAND2X1 U52392 ( .A(n50245), .B(n50244), .Y(n56568) );
  NOR2X1 U52393 ( .A(n50246), .B(n56568), .Y(n50248) );
  OR2X1 U52394 ( .A(n1757), .B(n43314), .Y(n50247) );
  NAND2X1 U52395 ( .A(n50248), .B(n50247), .Y(\mmu_ifetch_pc_w[31] ) );
  INVX1 U52396 ( .A(\mmu_ifetch_pc_w[31] ), .Y(n56619) );
  XNOR2X1 U52397 ( .A(u_mmu_itlb_va_addr_q[31]), .B(n56619), .Y(n50283) );
  NOR2X1 U52398 ( .A(n2221), .B(n43305), .Y(n50264) );
  NAND2X1 U52399 ( .A(n43309), .B(n56542), .Y(n50263) );
  NAND2X1 U52400 ( .A(n44840), .B(n58409), .Y(n57891) );
  NAND2X1 U52401 ( .A(n57891), .B(n50249), .Y(n50258) );
  XNOR2X1 U52402 ( .A(n50258), .B(n42437), .Y(n50250) );
  NOR2X1 U52403 ( .A(n50250), .B(n42873), .Y(n50256) );
  XNOR2X1 U52404 ( .A(n50251), .B(n42298), .Y(n50252) );
  XNOR2X1 U52405 ( .A(n50253), .B(n50252), .Y(n50254) );
  NOR2X1 U52406 ( .A(n50254), .B(n42930), .Y(n50255) );
  NOR2X1 U52407 ( .A(n50256), .B(n50255), .Y(n50261) );
  NAND2X1 U52408 ( .A(n30504), .B(n50257), .Y(n57892) );
  XNOR2X1 U52409 ( .A(n57892), .B(n50258), .Y(n50259) );
  NAND2X1 U52410 ( .A(n50259), .B(n54979), .Y(n50260) );
  NAND2X1 U52411 ( .A(n50261), .B(n50260), .Y(n56541) );
  NAND2X1 U52412 ( .A(n43311), .B(n56541), .Y(n50262) );
  NAND2X1 U52413 ( .A(n50263), .B(n50262), .Y(n56372) );
  NOR2X1 U52414 ( .A(n50264), .B(n56372), .Y(n50266) );
  OR2X1 U52415 ( .A(n1788), .B(n43314), .Y(n50265) );
  NAND2X1 U52416 ( .A(n50266), .B(n50265), .Y(n16) );
  XNOR2X1 U52417 ( .A(n16), .B(u_mmu_itlb_va_addr_q[30]), .Y(n50281) );
  NOR2X1 U52418 ( .A(n2177), .B(n43305), .Y(n50277) );
  NAND2X1 U52419 ( .A(n43309), .B(n55620), .Y(n50276) );
  NOR2X1 U52420 ( .A(n30479), .B(n37342), .Y(n50274) );
  NAND2X1 U52421 ( .A(n30469), .B(n54897), .Y(n50272) );
  XNOR2X1 U52422 ( .A(n37998), .B(n50269), .Y(n50270) );
  NAND2X1 U52423 ( .A(n54903), .B(n50270), .Y(n50271) );
  NAND2X1 U52424 ( .A(n50272), .B(n50271), .Y(n50273) );
  OR2X1 U52425 ( .A(n50274), .B(n50273), .Y(n55619) );
  NAND2X1 U52426 ( .A(n43311), .B(n55619), .Y(n50275) );
  NAND2X1 U52427 ( .A(n50276), .B(n50275), .Y(n55626) );
  NOR2X1 U52428 ( .A(n50277), .B(n55626), .Y(n50279) );
  OR2X1 U52429 ( .A(n1780), .B(n43314), .Y(n50278) );
  NAND2X1 U52430 ( .A(n50279), .B(n50278), .Y(n17) );
  XNOR2X1 U52431 ( .A(n17), .B(u_mmu_itlb_va_addr_q[22]), .Y(n50280) );
  NAND2X1 U52432 ( .A(n50281), .B(n50280), .Y(n50282) );
  NOR2X1 U52433 ( .A(n50283), .B(n50282), .Y(n50284) );
  NAND2X1 U52434 ( .A(n50285), .B(n50284), .Y(n50286) );
  NOR2X1 U52435 ( .A(n50287), .B(n50286), .Y(n50492) );
  NOR2X1 U52436 ( .A(n2151), .B(n43306), .Y(n50305) );
  NAND2X1 U52437 ( .A(n43308), .B(n55188), .Y(n50304) );
  NOR2X1 U52438 ( .A(n50289), .B(n42874), .Y(n50296) );
  XNOR2X1 U52439 ( .A(n50291), .B(n50290), .Y(n50292) );
  XOR2X1 U52440 ( .A(n50293), .B(n50292), .Y(n50294) );
  NOR2X1 U52441 ( .A(n50294), .B(n42931), .Y(n50295) );
  NOR2X1 U52442 ( .A(n50296), .B(n50295), .Y(n50302) );
  INVX1 U52443 ( .A(n50297), .Y(n50299) );
  XNOR2X1 U52444 ( .A(opcode_pc_w[14]), .B(opcode_opcode_w[14]), .Y(n50298) );
  XOR2X1 U52445 ( .A(n50299), .B(n50298), .Y(n50300) );
  NAND2X1 U52446 ( .A(n50300), .B(n54979), .Y(n50301) );
  NAND2X1 U52447 ( .A(n50302), .B(n50301), .Y(n55187) );
  NAND2X1 U52448 ( .A(n43311), .B(n55187), .Y(n50303) );
  NAND2X1 U52449 ( .A(n50304), .B(n50303), .Y(n55193) );
  NOR2X1 U52450 ( .A(n50305), .B(n55193), .Y(n50307) );
  OR2X1 U52451 ( .A(n1772), .B(n43314), .Y(n50306) );
  NAND2X1 U52452 ( .A(n50307), .B(n50306), .Y(n24) );
  XNOR2X1 U52453 ( .A(n24), .B(n17100), .Y(n50348) );
  NOR2X1 U52454 ( .A(n2145), .B(n43305), .Y(n50324) );
  NAND2X1 U52455 ( .A(n43308), .B(n55084), .Y(n50323) );
  NOR2X1 U52456 ( .A(n50309), .B(n42872), .Y(n50315) );
  NOR2X1 U52457 ( .A(n50313), .B(n42930), .Y(n50314) );
  NOR2X1 U52458 ( .A(n50315), .B(n50314), .Y(n50321) );
  INVX1 U52459 ( .A(n50316), .Y(n50318) );
  XNOR2X1 U52460 ( .A(opcode_pc_w[12]), .B(opcode_opcode_w[12]), .Y(n50317) );
  XOR2X1 U52461 ( .A(n50318), .B(n50317), .Y(n50319) );
  NAND2X1 U52462 ( .A(n50319), .B(n54979), .Y(n50320) );
  NAND2X1 U52463 ( .A(n50321), .B(n50320), .Y(n55083) );
  NAND2X1 U52464 ( .A(n43313), .B(n55083), .Y(n50322) );
  NAND2X1 U52465 ( .A(n50323), .B(n50322), .Y(n55088) );
  XNOR2X1 U52466 ( .A(n21), .B(n2684), .Y(n50346) );
  NOR2X1 U52467 ( .A(n2155), .B(n43306), .Y(n50342) );
  NAND2X1 U52468 ( .A(n43308), .B(n55248), .Y(n50341) );
  NOR2X1 U52469 ( .A(n50326), .B(n42873), .Y(n50333) );
  XNOR2X1 U52470 ( .A(n50328), .B(n50327), .Y(n50329) );
  XOR2X1 U52471 ( .A(n50330), .B(n50329), .Y(n50331) );
  NOR2X1 U52472 ( .A(n50331), .B(n42931), .Y(n50332) );
  NOR2X1 U52473 ( .A(n50333), .B(n50332), .Y(n50339) );
  INVX1 U52474 ( .A(n50334), .Y(n50336) );
  XNOR2X1 U52475 ( .A(n42729), .B(opcode_pc_w[15]), .Y(n50335) );
  XOR2X1 U52476 ( .A(n50336), .B(n50335), .Y(n50337) );
  NAND2X1 U52477 ( .A(n50337), .B(n54979), .Y(n50338) );
  NAND2X1 U52478 ( .A(n50339), .B(n50338), .Y(n55247) );
  NAND2X1 U52479 ( .A(n43311), .B(n55247), .Y(n50340) );
  NAND2X1 U52480 ( .A(n50341), .B(n50340), .Y(n55254) );
  NOR2X1 U52481 ( .A(n50342), .B(n55254), .Y(n50344) );
  OR2X1 U52482 ( .A(n1773), .B(n42845), .Y(n50343) );
  NAND2X1 U52483 ( .A(n50344), .B(n50343), .Y(n22) );
  XNOR2X1 U52484 ( .A(n22), .B(n2157), .Y(n50345) );
  NAND2X1 U52485 ( .A(n50346), .B(n50345), .Y(n50347) );
  NOR2X1 U52486 ( .A(n50348), .B(n50347), .Y(n50395) );
  NOR2X1 U52487 ( .A(n2165), .B(n43306), .Y(n50369) );
  NAND2X1 U52488 ( .A(n43308), .B(n55413), .Y(n50368) );
  NAND2X1 U52489 ( .A(opcode_pc_w[17]), .B(n44835), .Y(n50352) );
  NAND2X1 U52490 ( .A(n44840), .B(n58324), .Y(n50350) );
  NAND2X1 U52491 ( .A(n50350), .B(n50349), .Y(n50351) );
  NAND2X1 U52492 ( .A(n50352), .B(n50351), .Y(n50442) );
  NOR2X1 U52493 ( .A(n50353), .B(n42874), .Y(n50360) );
  XNOR2X1 U52494 ( .A(n50355), .B(n50354), .Y(n50356) );
  XOR2X1 U52495 ( .A(n50357), .B(n50356), .Y(n50358) );
  NOR2X1 U52496 ( .A(n50358), .B(n42930), .Y(n50359) );
  NOR2X1 U52497 ( .A(n50360), .B(n50359), .Y(n50366) );
  INVX1 U52498 ( .A(n50361), .Y(n50363) );
  XNOR2X1 U52499 ( .A(n42668), .B(opcode_pc_w[18]), .Y(n50362) );
  XOR2X1 U52500 ( .A(n50363), .B(n50362), .Y(n50364) );
  NAND2X1 U52501 ( .A(n50364), .B(n54979), .Y(n50365) );
  NAND2X1 U52502 ( .A(n50366), .B(n50365), .Y(n55412) );
  NAND2X1 U52503 ( .A(n43311), .B(n55412), .Y(n50367) );
  NAND2X1 U52504 ( .A(n50368), .B(n50367), .Y(n55419) );
  NOR2X1 U52505 ( .A(n50369), .B(n55419), .Y(n50371) );
  OR2X1 U52506 ( .A(n1776), .B(n42847), .Y(n50370) );
  NAND2X1 U52507 ( .A(n50371), .B(n50370), .Y(n10) );
  XNOR2X1 U52508 ( .A(n10), .B(n17102), .Y(n50393) );
  NOR2X1 U52509 ( .A(n2148), .B(n43305), .Y(n50389) );
  NAND2X1 U52510 ( .A(n43308), .B(n55133), .Y(n50388) );
  NOR2X1 U52511 ( .A(n50373), .B(n42872), .Y(n50380) );
  XNOR2X1 U52512 ( .A(n50375), .B(n50374), .Y(n50376) );
  XOR2X1 U52513 ( .A(n50377), .B(n50376), .Y(n50378) );
  NOR2X1 U52514 ( .A(n50378), .B(n42931), .Y(n50379) );
  NOR2X1 U52515 ( .A(n50380), .B(n50379), .Y(n50386) );
  INVX1 U52516 ( .A(n50381), .Y(n50383) );
  XNOR2X1 U52517 ( .A(opcode_pc_w[13]), .B(opcode_opcode_w[13]), .Y(n50382) );
  XOR2X1 U52518 ( .A(n50383), .B(n50382), .Y(n50384) );
  NAND2X1 U52519 ( .A(n50384), .B(n54979), .Y(n50385) );
  NAND2X1 U52520 ( .A(n50386), .B(n50385), .Y(n55132) );
  NAND2X1 U52521 ( .A(n43313), .B(n55132), .Y(n50387) );
  NAND2X1 U52522 ( .A(n50388), .B(n50387), .Y(n55137) );
  NOR2X1 U52523 ( .A(n50389), .B(n55137), .Y(n50391) );
  OR2X1 U52524 ( .A(n1771), .B(n42846), .Y(n50390) );
  NAND2X1 U52525 ( .A(n50391), .B(n50390), .Y(n9) );
  XNOR2X1 U52526 ( .A(n9), .B(n16237), .Y(n50392) );
  NOR2X1 U52527 ( .A(n50393), .B(n50392), .Y(n50394) );
  NAND2X1 U52528 ( .A(n50395), .B(n50394), .Y(n50490) );
  NOR2X1 U52529 ( .A(n2180), .B(n43306), .Y(n50407) );
  NAND2X1 U52530 ( .A(n43308), .B(n55667), .Y(n50406) );
  NOR2X1 U52531 ( .A(n30523), .B(n43014), .Y(n50404) );
  NAND2X1 U52532 ( .A(n30513), .B(n54897), .Y(n50402) );
  XNOR2X1 U52533 ( .A(n50399), .B(n50398), .Y(n50400) );
  NAND2X1 U52534 ( .A(n54903), .B(n50400), .Y(n50401) );
  NAND2X1 U52535 ( .A(n50402), .B(n50401), .Y(n50403) );
  OR2X1 U52536 ( .A(n50404), .B(n50403), .Y(n55666) );
  NAND2X1 U52537 ( .A(n43313), .B(n55666), .Y(n50405) );
  NAND2X1 U52538 ( .A(n50406), .B(n50405), .Y(n55674) );
  NOR2X1 U52539 ( .A(n50407), .B(n55674), .Y(n50409) );
  OR2X1 U52540 ( .A(n1781), .B(n42847), .Y(n50408) );
  NAND2X1 U52541 ( .A(n50409), .B(n50408), .Y(n15) );
  INVX1 U52542 ( .A(n15), .Y(n55672) );
  XNOR2X1 U52543 ( .A(u_mmu_itlb_va_addr_q[23]), .B(n55672), .Y(n50441) );
  NOR2X1 U52544 ( .A(n2183), .B(n43305), .Y(n50421) );
  NAND2X1 U52545 ( .A(n43308), .B(n55718), .Y(n50420) );
  NOR2X1 U52546 ( .A(n30632), .B(n37342), .Y(n50418) );
  NAND2X1 U52547 ( .A(n30616), .B(n54897), .Y(n50416) );
  XNOR2X1 U52548 ( .A(n50413), .B(n50412), .Y(n50414) );
  NAND2X1 U52549 ( .A(n54903), .B(n50414), .Y(n50415) );
  NAND2X1 U52550 ( .A(n50416), .B(n50415), .Y(n50417) );
  OR2X1 U52551 ( .A(n50418), .B(n50417), .Y(n55717) );
  NAND2X1 U52552 ( .A(n43313), .B(n55717), .Y(n50419) );
  NAND2X1 U52553 ( .A(n50420), .B(n50419), .Y(n55722) );
  NOR2X1 U52554 ( .A(n50421), .B(n55722), .Y(n50423) );
  OR2X1 U52555 ( .A(n1782), .B(n42846), .Y(n50422) );
  NAND2X1 U52556 ( .A(n50423), .B(n50422), .Y(n11) );
  XNOR2X1 U52557 ( .A(n11), .B(u_mmu_itlb_va_addr_q[24]), .Y(n50439) );
  NOR2X1 U52558 ( .A(n2174), .B(n43306), .Y(n50435) );
  NAND2X1 U52559 ( .A(n43308), .B(n55572), .Y(n50434) );
  NOR2X1 U52560 ( .A(n30604), .B(n43014), .Y(n50432) );
  NAND2X1 U52561 ( .A(n30594), .B(n54897), .Y(n50430) );
  XNOR2X1 U52562 ( .A(n50427), .B(n50426), .Y(n50428) );
  NAND2X1 U52563 ( .A(n54903), .B(n50428), .Y(n50429) );
  NAND2X1 U52564 ( .A(n50430), .B(n50429), .Y(n50431) );
  OR2X1 U52565 ( .A(n50432), .B(n50431), .Y(n55571) );
  NAND2X1 U52566 ( .A(n43311), .B(n55571), .Y(n50433) );
  NAND2X1 U52567 ( .A(n50434), .B(n50433), .Y(n55576) );
  NOR2X1 U52568 ( .A(n50435), .B(n55576), .Y(n50437) );
  OR2X1 U52569 ( .A(n1779), .B(n42846), .Y(n50436) );
  NAND2X1 U52570 ( .A(n50437), .B(n50436), .Y(n12) );
  XNOR2X1 U52571 ( .A(n12), .B(u_mmu_itlb_va_addr_q[21]), .Y(n50438) );
  NAND2X1 U52572 ( .A(n50439), .B(n50438), .Y(n50440) );
  NOR2X1 U52573 ( .A(n50441), .B(n50440), .Y(n50488) );
  NOR2X1 U52574 ( .A(n2168), .B(n43305), .Y(n50463) );
  NAND2X1 U52575 ( .A(n43308), .B(n55464), .Y(n50462) );
  NAND2X1 U52576 ( .A(opcode_pc_w[18]), .B(n44835), .Y(n50445) );
  NAND2X1 U52577 ( .A(n44841), .B(n58331), .Y(n50443) );
  NAND2X1 U52578 ( .A(n50443), .B(n50442), .Y(n50444) );
  NAND2X1 U52579 ( .A(n50445), .B(n50444), .Y(n57890) );
  XNOR2X1 U52580 ( .A(n42852), .B(opcode_pc_w[19]), .Y(n50446) );
  XOR2X1 U52581 ( .A(n57890), .B(n50446), .Y(n50447) );
  NOR2X1 U52582 ( .A(n50447), .B(n42873), .Y(n50454) );
  XNOR2X1 U52583 ( .A(n50449), .B(n50448), .Y(n50450) );
  XOR2X1 U52584 ( .A(n50451), .B(n50450), .Y(n50452) );
  NOR2X1 U52585 ( .A(n50452), .B(n42930), .Y(n50453) );
  NOR2X1 U52586 ( .A(n50454), .B(n50453), .Y(n50460) );
  INVX1 U52587 ( .A(n50455), .Y(n50457) );
  XNOR2X1 U52588 ( .A(n42793), .B(opcode_pc_w[19]), .Y(n50456) );
  XOR2X1 U52589 ( .A(n50457), .B(n50456), .Y(n50458) );
  NAND2X1 U52590 ( .A(n50458), .B(n54979), .Y(n50459) );
  NAND2X1 U52591 ( .A(n50460), .B(n50459), .Y(n55463) );
  NAND2X1 U52592 ( .A(n43313), .B(n55463), .Y(n50461) );
  NAND2X1 U52593 ( .A(n50462), .B(n50461), .Y(n55471) );
  NOR2X1 U52594 ( .A(n50463), .B(n55471), .Y(n50465) );
  OR2X1 U52595 ( .A(n1777), .B(n42847), .Y(n50464) );
  NAND2X1 U52596 ( .A(n50465), .B(n50464), .Y(n20) );
  INVX1 U52597 ( .A(n20), .Y(n55469) );
  XNOR2X1 U52598 ( .A(n2284), .B(n55469), .Y(n50486) );
  NOR2X1 U52599 ( .A(n1936), .B(n43306), .Y(n50482) );
  NAND2X1 U52600 ( .A(n43308), .B(n56166), .Y(n50481) );
  NAND2X1 U52601 ( .A(n44841), .B(n58396), .Y(n30456) );
  NAND2X1 U52602 ( .A(n30456), .B(n50466), .Y(n50476) );
  NAND2X1 U52603 ( .A(n30545), .B(n50475), .Y(n30445) );
  XOR2X1 U52604 ( .A(n50476), .B(n30445), .Y(n50467) );
  NOR2X1 U52605 ( .A(n50467), .B(n42874), .Y(n50474) );
  XNOR2X1 U52606 ( .A(n50469), .B(n50468), .Y(n50470) );
  XOR2X1 U52607 ( .A(n50471), .B(n50470), .Y(n50472) );
  NOR2X1 U52608 ( .A(n50472), .B(n42931), .Y(n50473) );
  NOR2X1 U52609 ( .A(n50474), .B(n50473), .Y(n50479) );
  NAND2X1 U52610 ( .A(n30559), .B(n50475), .Y(n30455) );
  XNOR2X1 U52611 ( .A(n50476), .B(n30455), .Y(n50477) );
  NAND2X1 U52612 ( .A(n50477), .B(n54979), .Y(n50478) );
  NAND2X1 U52613 ( .A(n50479), .B(n50478), .Y(n56165) );
  NAND2X1 U52614 ( .A(n43311), .B(n56165), .Y(n50480) );
  NAND2X1 U52615 ( .A(n50481), .B(n50480), .Y(n56171) );
  NOR2X1 U52616 ( .A(n50482), .B(n56171), .Y(n50484) );
  OR2X1 U52617 ( .A(n1786), .B(n42846), .Y(n50483) );
  NAND2X1 U52618 ( .A(n50484), .B(n50483), .Y(n18) );
  INVX1 U52619 ( .A(n18), .Y(n56169) );
  XNOR2X1 U52620 ( .A(u_mmu_itlb_va_addr_q[28]), .B(n56169), .Y(n50485) );
  NOR2X1 U52621 ( .A(n50486), .B(n50485), .Y(n50487) );
  NAND2X1 U52622 ( .A(n50488), .B(n50487), .Y(n50489) );
  NOR2X1 U52623 ( .A(n50490), .B(n50489), .Y(n50491) );
  NAND2X1 U52624 ( .A(n50492), .B(n50491), .Y(n52002) );
  NAND2X1 U52625 ( .A(n44073), .B(n52002), .Y(n58127) );
  NAND2X1 U52626 ( .A(n50493), .B(n58127), .Y(n55306) );
  INVX1 U52627 ( .A(mem_i_valid_i), .Y(n50494) );
  NAND2X1 U52628 ( .A(u_fetch_icache_fetch_q), .B(n50494), .Y(n57557) );
  NAND2X1 U52629 ( .A(n57557), .B(n73387), .Y(n55308) );
  INVX1 U52630 ( .A(n55308), .Y(n50495) );
  NAND2X1 U52631 ( .A(u_fetch_active_q), .B(n50495), .Y(n29013) );
  INVX1 U52632 ( .A(n29013), .Y(n55307) );
  NOR2X1 U52633 ( .A(n58126), .B(n51998), .Y(u_fetch_N157) );
  NAND2X1 U52634 ( .A(n8801), .B(n50496), .Y(n57600) );
  INVX1 U52635 ( .A(n57600), .Y(n73545) );
  NAND2X1 U52636 ( .A(mem_i_inst_i[19]), .B(n44085), .Y(n50498) );
  NAND2X1 U52637 ( .A(u_fetch_skid_buffer_q[19]), .B(n43407), .Y(n50497) );
  INVX1 U52638 ( .A(n50499), .Y(n50500) );
  NOR2X1 U52639 ( .A(n37561), .B(n42932), .Y(u_decode_N341) );
  NAND2X1 U52640 ( .A(n38001), .B(n42932), .Y(n50537) );
  NAND2X1 U52641 ( .A(n50537), .B(n44863), .Y(n54381) );
  NAND2X1 U52642 ( .A(challenge[33]), .B(n44855), .Y(n50501) );
  NAND2X1 U52643 ( .A(n54381), .B(n50501), .Y(n17241) );
  INVX1 U52644 ( .A(mem_i_inst_i[16]), .Y(n50502) );
  NOR2X1 U52645 ( .A(n50502), .B(n43405), .Y(net2358) );
  NOR2X1 U52646 ( .A(n8801), .B(n50503), .Y(n50505) );
  NOR2X1 U52647 ( .A(n57600), .B(n50502), .Y(n50504) );
  NOR2X1 U52648 ( .A(n50505), .B(n50504), .Y(n24517) );
  NOR2X1 U52649 ( .A(n24517), .B(n42932), .Y(u_decode_N338) );
  INVX1 U52650 ( .A(mem_i_inst_i[17]), .Y(n50506) );
  NOR2X1 U52651 ( .A(n43404), .B(n50506), .Y(net2359) );
  NAND2X1 U52652 ( .A(u_fetch_skid_buffer_q[17]), .B(n58511), .Y(n50508) );
  NAND2X1 U52653 ( .A(mem_i_inst_i[17]), .B(n44086), .Y(n50507) );
  NAND2X1 U52654 ( .A(n50508), .B(n50507), .Y(n24515) );
  INVX1 U52655 ( .A(n24515), .Y(n50509) );
  NOR2X1 U52656 ( .A(n50509), .B(n42934), .Y(u_decode_N339) );
  INVX1 U52657 ( .A(mem_i_inst_i[7]), .Y(n50510) );
  NOR2X1 U52658 ( .A(n50510), .B(n43405), .Y(net2344) );
  NAND2X1 U52659 ( .A(challenge[104]), .B(n44855), .Y(n50511) );
  NAND2X1 U52660 ( .A(n54437), .B(n50511), .Y(n17312) );
  NOR2X1 U52661 ( .A(n8801), .B(n50512), .Y(n50514) );
  NOR2X1 U52662 ( .A(n57600), .B(n50510), .Y(n50513) );
  NOR2X1 U52663 ( .A(n50514), .B(n50513), .Y(n24454) );
  NOR2X1 U52664 ( .A(n24454), .B(n42933), .Y(u_decode_N329) );
  INVX1 U52665 ( .A(mem_i_inst_i[11]), .Y(n50515) );
  NOR2X1 U52666 ( .A(n50515), .B(n43405), .Y(net2348) );
  NAND2X1 U52667 ( .A(u_fetch_skid_buffer_q[11]), .B(n58511), .Y(n50517) );
  NAND2X1 U52668 ( .A(mem_i_inst_i[11]), .B(n44086), .Y(n50516) );
  NAND2X1 U52669 ( .A(n50517), .B(n50516), .Y(n24519) );
  INVX1 U52670 ( .A(n24519), .Y(n621) );
  NOR2X1 U52671 ( .A(n621), .B(n42934), .Y(u_decode_N333) );
  INVX1 U52672 ( .A(mem_i_inst_i[10]), .Y(n50518) );
  NOR2X1 U52673 ( .A(n43404), .B(n50518), .Y(net2347) );
  NAND2X1 U52674 ( .A(u_fetch_skid_buffer_q[10]), .B(n58511), .Y(n50520) );
  NAND2X1 U52675 ( .A(mem_i_inst_i[10]), .B(n73545), .Y(n50519) );
  NAND2X1 U52676 ( .A(n50520), .B(n50519), .Y(n24528) );
  INVX1 U52677 ( .A(n24528), .Y(n50521) );
  NOR2X1 U52678 ( .A(n50521), .B(n42933), .Y(u_decode_N332) );
  INVX1 U52679 ( .A(mem_i_inst_i[8]), .Y(n50522) );
  NOR2X1 U52680 ( .A(n43404), .B(n50522), .Y(net2345) );
  NAND2X1 U52681 ( .A(u_fetch_skid_buffer_q[8]), .B(n58511), .Y(n50524) );
  NAND2X1 U52682 ( .A(mem_i_inst_i[8]), .B(n44086), .Y(n50523) );
  NAND2X1 U52683 ( .A(n50524), .B(n50523), .Y(n24530) );
  INVX1 U52684 ( .A(n24530), .Y(n50525) );
  NOR2X1 U52685 ( .A(n50525), .B(n42934), .Y(u_decode_N330) );
  INVX1 U52686 ( .A(mem_i_inst_i[9]), .Y(n50526) );
  NOR2X1 U52687 ( .A(n43404), .B(n50526), .Y(net2346) );
  NAND2X1 U52688 ( .A(u_fetch_skid_buffer_q[9]), .B(n43407), .Y(n50528) );
  NAND2X1 U52689 ( .A(mem_i_inst_i[9]), .B(n44086), .Y(n50527) );
  NAND2X1 U52690 ( .A(n50528), .B(n50527), .Y(n24529) );
  INVX1 U52691 ( .A(n24529), .Y(n50529) );
  NOR2X1 U52692 ( .A(n50529), .B(n42933), .Y(u_decode_N331) );
  NAND2X1 U52693 ( .A(n50530), .B(n28934), .Y(n28034) );
  INVX1 U52694 ( .A(n28034), .Y(n73544) );
  NAND2X1 U52695 ( .A(n29640), .B(n73544), .Y(n27326) );
  INVX1 U52696 ( .A(mem_i_inst_i[27]), .Y(n50531) );
  NOR2X1 U52697 ( .A(mem_i_error_i), .B(n50531), .Y(n50532) );
  NOR2X1 U52698 ( .A(u_fetch_fetch_page_fault_q), .B(n50532), .Y(n50533) );
  NOR2X1 U52699 ( .A(n50533), .B(n43317), .Y(net2370) );
  MX2X1 U52700 ( .A(n1836), .B(n50534), .S0(n8801), .Y(n50536) );
  NAND2X1 U52701 ( .A(mem_i_inst_i[27]), .B(n44086), .Y(n50535) );
  NAND2X1 U52702 ( .A(n50536), .B(n50535), .Y(n24469) );
  INVX1 U52703 ( .A(n50537), .Y(n50585) );
  NAND2X1 U52704 ( .A(n50585), .B(opcode_opcode_w[27]), .Y(n50539) );
  INVX1 U52705 ( .A(n42932), .Y(n57593) );
  NAND2X1 U52706 ( .A(n57593), .B(n24469), .Y(n50538) );
  NAND2X1 U52707 ( .A(n50539), .B(n50538), .Y(n8516) );
  INVX1 U52708 ( .A(mem_i_inst_i[28]), .Y(n50540) );
  NOR2X1 U52709 ( .A(n50540), .B(n43405), .Y(net2371) );
  NAND2X1 U52710 ( .A(u_fetch_skid_buffer_q[28]), .B(n43407), .Y(n50542) );
  NAND2X1 U52711 ( .A(mem_i_inst_i[28]), .B(n73545), .Y(n50541) );
  NAND2X1 U52712 ( .A(n50542), .B(n50541), .Y(n24436) );
  NAND2X1 U52713 ( .A(n50585), .B(opcode_opcode_w[28]), .Y(n50544) );
  NAND2X1 U52714 ( .A(n57593), .B(n24436), .Y(n50543) );
  NAND2X1 U52715 ( .A(n50544), .B(n50543), .Y(n8517) );
  INVX1 U52716 ( .A(mem_i_inst_i[31]), .Y(n50545) );
  NOR2X1 U52717 ( .A(n43404), .B(n50545), .Y(net2374) );
  NAND2X1 U52718 ( .A(u_fetch_skid_buffer_q[31]), .B(n43407), .Y(n50547) );
  NAND2X1 U52719 ( .A(mem_i_inst_i[31]), .B(n44085), .Y(n50546) );
  NAND2X1 U52720 ( .A(n50547), .B(n50546), .Y(n24557) );
  NAND2X1 U52721 ( .A(n50585), .B(n44835), .Y(n50549) );
  NAND2X1 U52722 ( .A(n57593), .B(n24557), .Y(n50548) );
  NAND2X1 U52723 ( .A(n50549), .B(n50548), .Y(n8538) );
  INVX1 U52724 ( .A(mem_i_inst_i[30]), .Y(n50550) );
  NOR2X1 U52725 ( .A(n43404), .B(n50550), .Y(net2373) );
  NAND2X1 U52726 ( .A(u_fetch_skid_buffer_q[30]), .B(n43407), .Y(n50552) );
  NAND2X1 U52727 ( .A(mem_i_inst_i[30]), .B(n44086), .Y(n50551) );
  NAND2X1 U52728 ( .A(n50552), .B(n50551), .Y(n24384) );
  NAND2X1 U52729 ( .A(n50585), .B(opcode_opcode_w[30]), .Y(n50554) );
  NAND2X1 U52730 ( .A(n57593), .B(n24384), .Y(n50553) );
  NAND2X1 U52731 ( .A(n50554), .B(n50553), .Y(n8519) );
  INVX1 U52732 ( .A(mem_i_inst_i[24]), .Y(n50555) );
  NOR2X1 U52733 ( .A(n43404), .B(n50555), .Y(net2366) );
  NAND2X1 U52734 ( .A(u_fetch_skid_buffer_q[24]), .B(n43407), .Y(n50557) );
  NAND2X1 U52735 ( .A(mem_i_inst_i[24]), .B(n44086), .Y(n50556) );
  NAND2X1 U52736 ( .A(n50557), .B(n50556), .Y(n24525) );
  NAND2X1 U52737 ( .A(n50585), .B(n42747), .Y(n50559) );
  NAND2X1 U52738 ( .A(n57593), .B(n24525), .Y(n50558) );
  NAND2X1 U52739 ( .A(n50559), .B(n50558), .Y(n8513) );
  INVX1 U52740 ( .A(mem_i_inst_i[26]), .Y(n50560) );
  NOR2X1 U52741 ( .A(n43404), .B(n50560), .Y(net2368) );
  NAND2X1 U52742 ( .A(u_fetch_skid_buffer_q[26]), .B(n43407), .Y(n50562) );
  NAND2X1 U52743 ( .A(mem_i_inst_i[26]), .B(n44086), .Y(n50561) );
  NAND2X1 U52744 ( .A(n50562), .B(n50561), .Y(n24556) );
  NAND2X1 U52745 ( .A(n50585), .B(opcode_opcode_w[26]), .Y(n50564) );
  NAND2X1 U52746 ( .A(n57593), .B(n24556), .Y(n50563) );
  NAND2X1 U52747 ( .A(n50564), .B(n50563), .Y(n8515) );
  INVX1 U52748 ( .A(mem_i_inst_i[22]), .Y(n58512) );
  NOR2X1 U52749 ( .A(n58512), .B(n43405), .Y(net2364) );
  NAND2X1 U52750 ( .A(u_fetch_skid_buffer_q[22]), .B(n43407), .Y(n24464) );
  NAND2X1 U52751 ( .A(mem_i_inst_i[22]), .B(n73545), .Y(n24435) );
  NAND2X1 U52752 ( .A(n24464), .B(n24435), .Y(n50565) );
  NAND2X1 U52753 ( .A(n57593), .B(n50565), .Y(n50567) );
  NAND2X1 U52754 ( .A(n50585), .B(n38064), .Y(n50566) );
  NAND2X1 U52755 ( .A(n50567), .B(n50566), .Y(n8511) );
  INVX1 U52756 ( .A(mem_i_inst_i[20]), .Y(n73558) );
  NOR2X1 U52757 ( .A(n73558), .B(n43405), .Y(net2362) );
  NAND2X1 U52758 ( .A(u_fetch_skid_buffer_q[20]), .B(n43407), .Y(n51401) );
  NAND2X1 U52759 ( .A(n73545), .B(mem_i_inst_i[20]), .Y(n50568) );
  NAND2X1 U52760 ( .A(n51401), .B(n50568), .Y(n24437) );
  INVX1 U52761 ( .A(n24437), .Y(n51960) );
  NOR2X1 U52762 ( .A(n51960), .B(n42934), .Y(u_decode_N342) );
  INVX1 U52763 ( .A(mem_i_inst_i[21]), .Y(n50569) );
  NOR2X1 U52764 ( .A(n50569), .B(n43405), .Y(net2363) );
  NAND2X1 U52765 ( .A(u_fetch_skid_buffer_q[21]), .B(n43407), .Y(n50571) );
  NAND2X1 U52766 ( .A(mem_i_inst_i[21]), .B(n44085), .Y(n50570) );
  NAND2X1 U52767 ( .A(n50571), .B(n50570), .Y(n58514) );
  NAND2X1 U52768 ( .A(n57593), .B(n58514), .Y(n51958) );
  INVX1 U52769 ( .A(n51958), .Y(n73540) );
  INVX1 U52770 ( .A(mem_i_inst_i[29]), .Y(n50572) );
  NOR2X1 U52771 ( .A(n43404), .B(n50572), .Y(net2372) );
  NAND2X1 U52772 ( .A(u_fetch_skid_buffer_q[29]), .B(n43407), .Y(n50574) );
  NAND2X1 U52773 ( .A(mem_i_inst_i[29]), .B(n44085), .Y(n50573) );
  NAND2X1 U52774 ( .A(n50574), .B(n50573), .Y(n24445) );
  NAND2X1 U52775 ( .A(n50585), .B(opcode_opcode_w[29]), .Y(n50576) );
  NAND2X1 U52776 ( .A(n57593), .B(n24445), .Y(n50575) );
  NAND2X1 U52777 ( .A(n50576), .B(n50575), .Y(n8518) );
  INVX1 U52778 ( .A(mem_i_inst_i[23]), .Y(n50577) );
  NOR2X1 U52779 ( .A(n43404), .B(n50577), .Y(net2365) );
  NAND2X1 U52780 ( .A(u_fetch_skid_buffer_q[23]), .B(n43407), .Y(n50579) );
  NAND2X1 U52781 ( .A(mem_i_inst_i[23]), .B(n44085), .Y(n50578) );
  NAND2X1 U52782 ( .A(n50579), .B(n50578), .Y(n24524) );
  NAND2X1 U52783 ( .A(n50585), .B(n40454), .Y(n50581) );
  NAND2X1 U52784 ( .A(n57593), .B(n24524), .Y(n50580) );
  NAND2X1 U52785 ( .A(n50581), .B(n50580), .Y(n8512) );
  INVX1 U52786 ( .A(mem_i_inst_i[25]), .Y(n50582) );
  NOR2X1 U52787 ( .A(n50582), .B(n43405), .Y(net2367) );
  NAND2X1 U52788 ( .A(u_fetch_skid_buffer_q[25]), .B(n43406), .Y(n50584) );
  NAND2X1 U52789 ( .A(mem_i_inst_i[25]), .B(n44085), .Y(n50583) );
  NAND2X1 U52790 ( .A(n50584), .B(n50583), .Y(n24455) );
  NAND2X1 U52791 ( .A(n50585), .B(opcode_opcode_w[25]), .Y(n50587) );
  NAND2X1 U52792 ( .A(n57593), .B(n24455), .Y(n50586) );
  NAND2X1 U52793 ( .A(n50587), .B(n50586), .Y(n8514) );
  NOR2X1 U52794 ( .A(n28765), .B(n57380), .Y(n50588) );
  NAND2X1 U52795 ( .A(n50588), .B(n37550), .Y(n57918) );
  NAND2X1 U52796 ( .A(u_mmu_state_q[1]), .B(n57380), .Y(n57915) );
  NAND2X1 U52797 ( .A(n57918), .B(n57915), .Y(n8556) );
  OR2X1 U52798 ( .A(n28765), .B(n57915), .Y(n50590) );
  INVX1 U52799 ( .A(n57918), .Y(n57395) );
  NAND2X1 U52800 ( .A(n30273), .B(n28796), .Y(n57394) );
  NAND2X1 U52801 ( .A(n57395), .B(n57394), .Y(n50589) );
  NAND2X1 U52802 ( .A(n50590), .B(n50589), .Y(n28797) );
  INVX1 U52803 ( .A(mem_i_inst_i[5]), .Y(n50591) );
  NOR2X1 U52804 ( .A(n50591), .B(n43405), .Y(net2342) );
  NAND2X1 U52805 ( .A(n43319), .B(n58506), .Y(n58510) );
  NAND2X1 U52806 ( .A(mem_i_inst_i[4]), .B(n43319), .Y(n50592) );
  NAND2X1 U52807 ( .A(n58510), .B(n50592), .Y(net2341) );
  NAND2X1 U52808 ( .A(u_fetch_skid_buffer_q[4]), .B(n43406), .Y(n50593) );
  NAND2X1 U52809 ( .A(n24839), .B(n50593), .Y(n24535) );
  NAND2X1 U52810 ( .A(u_fetch_skid_buffer_q[5]), .B(n43406), .Y(n50595) );
  NAND2X1 U52811 ( .A(mem_i_inst_i[5]), .B(n44085), .Y(n50594) );
  NAND2X1 U52812 ( .A(n50595), .B(n50594), .Y(n51121) );
  NOR2X1 U52813 ( .A(n51121), .B(n37565), .Y(n50596) );
  INVX1 U52814 ( .A(n24535), .Y(n50648) );
  NAND2X1 U52815 ( .A(n50596), .B(n50648), .Y(n24389) );
  INVX1 U52816 ( .A(mem_i_inst_i[14]), .Y(n50597) );
  NOR2X1 U52817 ( .A(n50597), .B(n43405), .Y(net2351) );
  INVX1 U52818 ( .A(mem_i_inst_i[13]), .Y(n50598) );
  NOR2X1 U52819 ( .A(n50598), .B(n43405), .Y(net2350) );
  INVX1 U52820 ( .A(mem_i_inst_i[12]), .Y(n50599) );
  NOR2X1 U52821 ( .A(n50599), .B(n43405), .Y(net2349) );
  NAND2X1 U52822 ( .A(u_fetch_skid_buffer_q[12]), .B(n43406), .Y(n50601) );
  NAND2X1 U52823 ( .A(mem_i_inst_i[12]), .B(n44085), .Y(n50600) );
  NAND2X1 U52824 ( .A(n50601), .B(n50600), .Y(n50634) );
  INVX1 U52825 ( .A(n50634), .Y(n57411) );
  NAND2X1 U52826 ( .A(mem_i_inst_i[13]), .B(n44085), .Y(n50603) );
  NAND2X1 U52827 ( .A(u_fetch_skid_buffer_q[13]), .B(n43406), .Y(n50602) );
  NAND2X1 U52828 ( .A(n50603), .B(n50602), .Y(n50633) );
  INVX1 U52829 ( .A(n50633), .Y(n73536) );
  NAND2X1 U52830 ( .A(n57411), .B(n73536), .Y(n24388) );
  NAND2X1 U52831 ( .A(u_fetch_skid_buffer_q[14]), .B(n43406), .Y(n50605) );
  NAND2X1 U52832 ( .A(mem_i_inst_i[14]), .B(n44085), .Y(n50604) );
  NAND2X1 U52833 ( .A(n50605), .B(n50604), .Y(n57579) );
  INVX1 U52834 ( .A(n24388), .Y(n50609) );
  NAND2X1 U52835 ( .A(n42424), .B(n50609), .Y(n57405) );
  NOR2X1 U52836 ( .A(n24389), .B(n57405), .Y(u_decode_N768) );
  NAND2X1 U52837 ( .A(challenge[31]), .B(n44855), .Y(n50606) );
  NAND2X1 U52838 ( .A(n54381), .B(n50606), .Y(n17239) );
  INVX1 U52839 ( .A(n57579), .Y(n73537) );
  NAND2X1 U52840 ( .A(n37570), .B(n73537), .Y(n24416) );
  INVX1 U52841 ( .A(n24416), .Y(n50607) );
  NAND2X1 U52842 ( .A(n57593), .B(n50607), .Y(n55035) );
  NOR2X1 U52843 ( .A(n24389), .B(n55035), .Y(u_decode_N767) );
  NAND2X1 U52844 ( .A(challenge[30]), .B(n44855), .Y(n50608) );
  NAND2X1 U52845 ( .A(n54381), .B(n50608), .Y(n17238) );
  NAND2X1 U52846 ( .A(n73536), .B(n50634), .Y(n57580) );
  INVX1 U52847 ( .A(n57580), .Y(n73535) );
  NAND2X1 U52848 ( .A(n73535), .B(n73537), .Y(n73388) );
  INVX1 U52849 ( .A(n73388), .Y(n73534) );
  NAND2X1 U52850 ( .A(n57593), .B(n73534), .Y(n57414) );
  NOR2X1 U52851 ( .A(n24389), .B(n57414), .Y(u_decode_N766) );
  NAND2X1 U52852 ( .A(n73537), .B(n50609), .Y(n57567) );
  INVX1 U52853 ( .A(n57567), .Y(n73533) );
  NAND2X1 U52854 ( .A(n57593), .B(n73533), .Y(n57415) );
  NOR2X1 U52855 ( .A(n24389), .B(n57415), .Y(u_decode_N765) );
  NOR2X1 U52856 ( .A(n1855), .B(n1853), .Y(n50610) );
  NAND2X1 U52857 ( .A(n50610), .B(n73363), .Y(n28949) );
  NAND2X1 U52858 ( .A(n37570), .B(n42424), .Y(n57404) );
  NOR2X1 U52859 ( .A(n24389), .B(n57404), .Y(u_decode_N770) );
  NAND2X1 U52860 ( .A(n42424), .B(n73535), .Y(n57407) );
  NOR2X1 U52861 ( .A(n24389), .B(n57407), .Y(u_decode_N769) );
  NOR2X1 U52862 ( .A(n28949), .B(n50611), .Y(n50613) );
  NOR2X1 U52863 ( .A(n1849), .B(n1850), .Y(n50612) );
  NAND2X1 U52864 ( .A(n50613), .B(n50612), .Y(n15219) );
  NAND2X1 U52865 ( .A(opcode_instr_w_41), .B(n57351), .Y(n57902) );
  NAND2X1 U52866 ( .A(n57351), .B(n15219), .Y(n50619) );
  INVX1 U52867 ( .A(n50619), .Y(n54286) );
  MX2X1 U52868 ( .A(n50700), .B(n42740), .S0(n54286), .Y(n50615) );
  NOR2X1 U52869 ( .A(n43376), .B(n50615), .Y(n50614) );
  XNOR2X1 U52870 ( .A(n39625), .B(n50614), .Y(n73431) );
  INVX1 U52871 ( .A(n73431), .Y(n57364) );
  MX2X1 U52872 ( .A(n57429), .B(n42762), .S0(n54286), .Y(n54274) );
  INVX1 U52873 ( .A(n54274), .Y(n54273) );
  XNOR2X1 U52874 ( .A(n42296), .B(n54273), .Y(n50616) );
  NOR2X1 U52875 ( .A(n43377), .B(n50616), .Y(n50617) );
  XNOR2X1 U52876 ( .A(n43461), .B(n50617), .Y(n73430) );
  INVX1 U52877 ( .A(n73430), .Y(n57365) );
  NAND2X1 U52878 ( .A(n57364), .B(n57365), .Y(n57350) );
  NAND2X1 U52879 ( .A(n57351), .B(n57350), .Y(n50618) );
  OR2X1 U52880 ( .A(n15318), .B(n50618), .Y(n57560) );
  INVX1 U52881 ( .A(n57560), .Y(n57353) );
  NOR2X1 U52882 ( .A(n57353), .B(n50619), .Y(u_lsu_N103) );
  NOR2X1 U52883 ( .A(n24535), .B(n37565), .Y(n50620) );
  NAND2X1 U52884 ( .A(n50620), .B(n51121), .Y(n58517) );
  NOR2X1 U52885 ( .A(n57415), .B(n58517), .Y(u_decode_N771) );
  INVX1 U52886 ( .A(n24533), .Y(n50621) );
  NAND2X1 U52887 ( .A(n24535), .B(n50621), .Y(n606) );
  NAND2X1 U52888 ( .A(mem_i_inst_i[6]), .B(n43319), .Y(n50622) );
  NAND2X1 U52889 ( .A(n58510), .B(n50622), .Y(net2343) );
  NAND2X1 U52890 ( .A(u_fetch_skid_buffer_q[6]), .B(n43406), .Y(n50623) );
  NAND2X1 U52891 ( .A(n24845), .B(n50623), .Y(n24473) );
  INVX1 U52892 ( .A(n606), .Y(n50636) );
  NAND2X1 U52893 ( .A(n37558), .B(n24473), .Y(n24422) );
  NOR2X1 U52894 ( .A(n24422), .B(n57414), .Y(u_decode_N777) );
  NOR2X1 U52895 ( .A(n24473), .B(n24384), .Y(n50626) );
  INVX1 U52896 ( .A(n24448), .Y(n50624) );
  NOR2X1 U52897 ( .A(n24455), .B(n50624), .Y(n50625) );
  NAND2X1 U52898 ( .A(n50625), .B(n37558), .Y(n51959) );
  INVX1 U52899 ( .A(n51959), .Y(n73529) );
  NAND2X1 U52900 ( .A(n24552), .B(n73529), .Y(n50628) );
  INVX1 U52901 ( .A(n50628), .Y(n57581) );
  NAND2X1 U52902 ( .A(n50626), .B(n57581), .Y(n24409) );
  NOR2X1 U52903 ( .A(n24409), .B(n57404), .Y(u_decode_N752) );
  NOR2X1 U52904 ( .A(n24409), .B(n57415), .Y(u_decode_N747) );
  NAND2X1 U52905 ( .A(challenge[29]), .B(n44855), .Y(n50627) );
  NAND2X1 U52906 ( .A(n54381), .B(n50627), .Y(n17237) );
  NAND2X1 U52907 ( .A(n37572), .B(n42424), .Y(n57406) );
  NOR2X1 U52908 ( .A(n24409), .B(n57406), .Y(u_decode_N753) );
  NOR2X1 U52909 ( .A(n24409), .B(n57407), .Y(u_decode_N755) );
  NOR2X1 U52910 ( .A(n24473), .B(n57567), .Y(n50630) );
  INVX1 U52911 ( .A(n24384), .Y(n51119) );
  NOR2X1 U52912 ( .A(n51119), .B(n50628), .Y(n50629) );
  NAND2X1 U52913 ( .A(n50630), .B(n50629), .Y(n24410) );
  NOR2X1 U52914 ( .A(n24410), .B(n42933), .Y(u_decode_N748) );
  INVX1 U52915 ( .A(n57407), .Y(n50642) );
  NAND2X1 U52916 ( .A(n50642), .B(n24384), .Y(n50632) );
  INVX1 U52917 ( .A(n24473), .Y(n51408) );
  NAND2X1 U52918 ( .A(n57581), .B(n51408), .Y(n50631) );
  NOR2X1 U52919 ( .A(n50632), .B(n50631), .Y(u_decode_N756) );
  NOR2X1 U52920 ( .A(n24409), .B(n57414), .Y(u_decode_N754) );
  NAND2X1 U52921 ( .A(n42425), .B(n73537), .Y(n57413) );
  INVX1 U52922 ( .A(n57413), .Y(n50635) );
  NAND2X1 U52923 ( .A(n50635), .B(n50634), .Y(n58129) );
  NOR2X1 U52924 ( .A(n24409), .B(n58129), .Y(u_decode_N750) );
  NOR2X1 U52925 ( .A(n24409), .B(n57405), .Y(u_decode_N751) );
  NOR2X1 U52926 ( .A(n24409), .B(n55035), .Y(u_decode_N749) );
  INVX1 U52927 ( .A(n51121), .Y(n57401) );
  NAND2X1 U52928 ( .A(n37568), .B(n50636), .Y(n24378) );
  NOR2X1 U52929 ( .A(n24378), .B(n57406), .Y(u_decode_N736) );
  NOR2X1 U52930 ( .A(n24378), .B(n57415), .Y(u_decode_N737) );
  NOR2X1 U52931 ( .A(n24378), .B(n57405), .Y(u_decode_N741) );
  NOR2X1 U52932 ( .A(n24378), .B(n57404), .Y(u_decode_N740) );
  INVX1 U52933 ( .A(n24378), .Y(n50637) );
  NAND2X1 U52934 ( .A(n57411), .B(n50637), .Y(n50638) );
  NOR2X1 U52935 ( .A(n57413), .B(n50638), .Y(u_decode_N738) );
  NOR2X1 U52936 ( .A(n24378), .B(n58129), .Y(u_decode_N739) );
  NOR2X1 U52937 ( .A(n1851), .B(opcode_instr_w[5]), .Y(n50640) );
  NOR2X1 U52938 ( .A(n1890), .B(n1854), .Y(n50639) );
  NAND2X1 U52939 ( .A(n50640), .B(n50639), .Y(n17938) );
  NAND2X1 U52940 ( .A(n24488), .B(n57401), .Y(n24385) );
  INVX1 U52941 ( .A(n24385), .Y(n73528) );
  NAND2X1 U52942 ( .A(n50642), .B(n73528), .Y(n50641) );
  NOR2X1 U52943 ( .A(n51119), .B(n50641), .Y(u_decode_N744) );
  NAND2X1 U52944 ( .A(n50642), .B(n51119), .Y(n50643) );
  NOR2X1 U52945 ( .A(n24385), .B(n50643), .Y(u_decode_N743) );
  NAND2X1 U52946 ( .A(n51119), .B(n73528), .Y(n50644) );
  NOR2X1 U52947 ( .A(n57414), .B(n50644), .Y(u_decode_N742) );
  INVX1 U52948 ( .A(mem_i_inst_i[3]), .Y(n50645) );
  NOR2X1 U52949 ( .A(n50645), .B(n43405), .Y(net2340) );
  NAND2X1 U52950 ( .A(u_fetch_skid_buffer_q[3]), .B(n43406), .Y(n50647) );
  NAND2X1 U52951 ( .A(mem_i_inst_i[3]), .B(n44085), .Y(n50646) );
  NAND2X1 U52952 ( .A(n50647), .B(n50646), .Y(n24429) );
  NOR2X1 U52953 ( .A(n24429), .B(n24473), .Y(n50650) );
  NOR2X1 U52954 ( .A(n24539), .B(n50648), .Y(n50649) );
  NAND2X1 U52955 ( .A(n50650), .B(n50649), .Y(n24405) );
  INVX1 U52956 ( .A(n24405), .Y(n50651) );
  NAND2X1 U52957 ( .A(n57593), .B(n50651), .Y(n50652) );
  NOR2X1 U52958 ( .A(n57401), .B(n50652), .Y(u_decode_N745) );
  AND2X1 U52959 ( .A(n24538), .B(n51121), .Y(n50653) );
  NAND2X1 U52960 ( .A(n50653), .B(n24473), .Y(n57561) );
  OR2X1 U52961 ( .A(n57561), .B(n57415), .Y(n50654) );
  NOR2X1 U52962 ( .A(n24429), .B(n50654), .Y(u_decode_N758) );
  INVX1 U52963 ( .A(n57561), .Y(n50655) );
  NAND2X1 U52964 ( .A(n57593), .B(n57401), .Y(n50656) );
  NOR2X1 U52965 ( .A(n24405), .B(n50656), .Y(u_decode_N746) );
  NAND2X1 U52966 ( .A(n50658), .B(n50657), .Y(n1009) );
  INVX1 U52967 ( .A(n17938), .Y(n50659) );
  NAND2X1 U52968 ( .A(n42434), .B(n50659), .Y(n50844) );
  INVX1 U52969 ( .A(n50844), .Y(n50664) );
  NAND2X1 U52970 ( .A(n50682), .B(n50678), .Y(n50854) );
  NOR2X1 U52971 ( .A(opcode_instr_w_18), .B(opcode_instr_w_16), .Y(n50660) );
  NAND2X1 U52972 ( .A(n50660), .B(n50856), .Y(n50689) );
  NAND2X1 U52973 ( .A(n50661), .B(n50858), .Y(n50673) );
  NOR2X1 U52974 ( .A(n50689), .B(n50673), .Y(n50662) );
  NAND2X1 U52975 ( .A(n50662), .B(n50850), .Y(n50681) );
  NOR2X1 U52976 ( .A(n50854), .B(n50681), .Y(n50663) );
  NAND2X1 U52977 ( .A(n50663), .B(n58540), .Y(n58556) );
  NAND2X1 U52978 ( .A(n50664), .B(n43412), .Y(n50695) );
  NAND2X1 U52979 ( .A(n50665), .B(n57095), .Y(n50671) );
  INVX1 U52980 ( .A(n50671), .Y(n50666) );
  NAND2X1 U52981 ( .A(n50666), .B(n57096), .Y(n50845) );
  NOR2X1 U52982 ( .A(n50695), .B(n50845), .Y(n50667) );
  NAND2X1 U52983 ( .A(n50667), .B(n50694), .Y(n50669) );
  INVX1 U52984 ( .A(n50669), .Y(n50668) );
  NAND2X1 U52985 ( .A(opcode_instr_w[10]), .B(n50668), .Y(n56998) );
  NAND2X1 U52986 ( .A(n56998), .B(n56824), .Y(n56852) );
  NOR2X1 U52987 ( .A(n1851), .B(n1926), .Y(n50670) );
  NAND2X1 U52988 ( .A(n50670), .B(n57096), .Y(n50693) );
  INVX1 U52989 ( .A(n50695), .Y(n57099) );
  NAND2X1 U52990 ( .A(n57099), .B(n50671), .Y(n50672) );
  NOR2X1 U52991 ( .A(opcode_instr_w[6]), .B(n50672), .Y(n50676) );
  INVX1 U52992 ( .A(n50673), .Y(n50674) );
  NOR2X1 U52993 ( .A(n50674), .B(n50689), .Y(n50675) );
  NOR2X1 U52994 ( .A(n50676), .B(n50675), .Y(n50688) );
  NOR2X1 U52995 ( .A(n1890), .B(n1009), .Y(n50677) );
  NOR2X1 U52996 ( .A(opcode_instr_w_1), .B(n50677), .Y(n50680) );
  NAND2X1 U52997 ( .A(n58540), .B(n50678), .Y(n50679) );
  NOR2X1 U52998 ( .A(n50680), .B(n50679), .Y(n50684) );
  INVX1 U52999 ( .A(n50681), .Y(n57094) );
  NAND2X1 U53000 ( .A(n57094), .B(n50682), .Y(n50683) );
  NOR2X1 U53001 ( .A(n50684), .B(n50683), .Y(n50686) );
  NOR2X1 U53002 ( .A(opcode_instr_w[11]), .B(n50850), .Y(n50685) );
  NOR2X1 U53003 ( .A(n50686), .B(n50685), .Y(n50687) );
  NAND2X1 U53004 ( .A(n50688), .B(n50687), .Y(n58544) );
  NOR2X1 U53005 ( .A(n50689), .B(n58544), .Y(n50691) );
  NOR2X1 U53006 ( .A(opcode_instr_w[5]), .B(opcode_instr_w_1), .Y(n50690) );
  NAND2X1 U53007 ( .A(n50691), .B(n50690), .Y(n50692) );
  NOR2X1 U53008 ( .A(n40679), .B(n43269), .Y(n50698) );
  NOR2X1 U53009 ( .A(n50695), .B(n50694), .Y(n50697) );
  INVX1 U53010 ( .A(n50845), .Y(n50696) );
  NAND2X1 U53011 ( .A(n50697), .B(n50696), .Y(n56993) );
  NAND2X1 U53012 ( .A(n50698), .B(n56993), .Y(n50699) );
  NAND2X1 U53013 ( .A(n42439), .B(n50699), .Y(n50701) );
  NOR2X1 U53014 ( .A(n57436), .B(n50701), .Y(u_exec_N240) );
  NOR2X1 U53015 ( .A(n54586), .B(n50701), .Y(u_exec_N242) );
  NOR2X1 U53016 ( .A(n57429), .B(n50701), .Y(u_exec_N239) );
  NOR2X1 U53017 ( .A(n50700), .B(n50701), .Y(u_exec_N238) );
  NOR2X1 U53018 ( .A(n54447), .B(n50701), .Y(u_exec_N241) );
  NOR2X1 U53019 ( .A(n15716), .B(n15717), .Y(n50703) );
  NOR2X1 U53020 ( .A(n15761), .B(n15762), .Y(n50702) );
  NAND2X1 U53021 ( .A(n50703), .B(n50702), .Y(u_exec_alu_p_w[3]) );
  NOR2X1 U53022 ( .A(n44364), .B(n43074), .Y(n50705) );
  NOR2X1 U53023 ( .A(n44361), .B(n43077), .Y(n50704) );
  NOR2X1 U53024 ( .A(n50705), .B(n50704), .Y(n50707) );
  NOR2X1 U53025 ( .A(n22856), .B(n22855), .Y(n50706) );
  NAND2X1 U53026 ( .A(n50707), .B(n50706), .Y(u_decode_u_regfile_N1213) );
  NOR2X1 U53027 ( .A(n44442), .B(n43076), .Y(n50709) );
  NOR2X1 U53028 ( .A(n44439), .B(n37664), .Y(n50708) );
  NOR2X1 U53029 ( .A(n50709), .B(n50708), .Y(n50711) );
  NOR2X1 U53030 ( .A(n21616), .B(n21615), .Y(n50710) );
  NAND2X1 U53031 ( .A(n50711), .B(n50710), .Y(u_decode_u_regfile_N325) );
  NOR2X1 U53032 ( .A(n44382), .B(n43076), .Y(n50713) );
  NOR2X1 U53033 ( .A(n44379), .B(n37664), .Y(n50712) );
  NOR2X1 U53034 ( .A(n50713), .B(n50712), .Y(n50715) );
  NOR2X1 U53035 ( .A(n22596), .B(n22595), .Y(n50714) );
  NAND2X1 U53036 ( .A(n50715), .B(n50714), .Y(u_decode_u_regfile_N140) );
  NOR2X1 U53037 ( .A(n44304), .B(n43076), .Y(n50717) );
  NOR2X1 U53038 ( .A(n44301), .B(n37664), .Y(n50716) );
  NOR2X1 U53039 ( .A(n50717), .B(n50716), .Y(n50719) );
  NOR2X1 U53040 ( .A(n23950), .B(n23949), .Y(n50718) );
  NAND2X1 U53041 ( .A(n50719), .B(n50718), .Y(u_decode_u_regfile_N1028) );
  NOR2X1 U53042 ( .A(n44406), .B(n43076), .Y(n50722) );
  NOR2X1 U53043 ( .A(n44403), .B(n43078), .Y(n50721) );
  NOR2X1 U53044 ( .A(n50722), .B(n50721), .Y(n50724) );
  NOR2X1 U53045 ( .A(n22204), .B(n22203), .Y(n50723) );
  NAND2X1 U53046 ( .A(n50724), .B(n50723), .Y(u_decode_u_regfile_N214) );
  NAND2X1 U53047 ( .A(writeback_exec_idx_w[4]), .B(n39766), .Y(n50791) );
  INVX1 U53048 ( .A(n50791), .Y(n50753) );
  NOR2X1 U53049 ( .A(n44559), .B(n43075), .Y(n50726) );
  NOR2X1 U53050 ( .A(n44556), .B(n43078), .Y(n50725) );
  NOR2X1 U53051 ( .A(n50726), .B(n50725), .Y(n50728) );
  NOR2X1 U53052 ( .A(n19454), .B(n19453), .Y(n50727) );
  NAND2X1 U53053 ( .A(n50728), .B(n50727), .Y(u_decode_u_regfile_N732) );
  NOR2X1 U53054 ( .A(n44328), .B(n43075), .Y(n50730) );
  NOR2X1 U53055 ( .A(n44325), .B(n43078), .Y(n50729) );
  NOR2X1 U53056 ( .A(n50730), .B(n50729), .Y(n50732) );
  NOR2X1 U53057 ( .A(n23510), .B(n23509), .Y(n50731) );
  NAND2X1 U53058 ( .A(n50732), .B(n50731), .Y(u_decode_u_regfile_N1102) );
  NOR2X1 U53059 ( .A(n44430), .B(n43075), .Y(n50734) );
  NOR2X1 U53060 ( .A(n44427), .B(n43078), .Y(n50733) );
  NOR2X1 U53061 ( .A(n50734), .B(n50733), .Y(n50736) );
  NOR2X1 U53062 ( .A(n21812), .B(n21811), .Y(n50735) );
  NAND2X1 U53063 ( .A(n50736), .B(n50735), .Y(u_decode_u_regfile_N288) );
  NOR2X1 U53064 ( .A(n44418), .B(n43075), .Y(n50738) );
  NOR2X1 U53065 ( .A(n44415), .B(n43078), .Y(n50737) );
  NOR2X1 U53066 ( .A(n50738), .B(n50737), .Y(n50740) );
  NOR2X1 U53067 ( .A(n22008), .B(n22007), .Y(n50739) );
  NAND2X1 U53068 ( .A(n50740), .B(n50739), .Y(u_decode_u_regfile_N251) );
  NOR2X1 U53069 ( .A(n44472), .B(n43075), .Y(n50742) );
  NOR2X1 U53070 ( .A(n44469), .B(n43078), .Y(n50741) );
  NOR2X1 U53071 ( .A(n50742), .B(n50741), .Y(n50744) );
  NOR2X1 U53072 ( .A(n21026), .B(n21025), .Y(n50743) );
  NAND2X1 U53073 ( .A(n50744), .B(n50743), .Y(u_decode_u_regfile_N436) );
  NOR2X1 U53074 ( .A(n44583), .B(n43075), .Y(n50746) );
  NOR2X1 U53075 ( .A(n44580), .B(n43078), .Y(n50745) );
  NOR2X1 U53076 ( .A(n50746), .B(n50745), .Y(n50748) );
  NOR2X1 U53077 ( .A(n18670), .B(n18669), .Y(n50747) );
  NAND2X1 U53078 ( .A(n50748), .B(n50747), .Y(u_decode_u_regfile_N880) );
  NOR2X1 U53079 ( .A(n44571), .B(n43075), .Y(n50750) );
  NOR2X1 U53080 ( .A(n44568), .B(n43078), .Y(n50749) );
  NOR2X1 U53081 ( .A(n50750), .B(n50749), .Y(n50752) );
  NOR2X1 U53082 ( .A(n19062), .B(n19061), .Y(n50751) );
  NAND2X1 U53083 ( .A(n50752), .B(n50751), .Y(u_decode_u_regfile_N806) );
  NOR2X1 U53084 ( .A(n44592), .B(n43075), .Y(n50755) );
  NOR2X1 U53085 ( .A(n44589), .B(n43078), .Y(n50754) );
  NOR2X1 U53086 ( .A(n50755), .B(n50754), .Y(n50757) );
  NOR2X1 U53087 ( .A(n18476), .B(n18475), .Y(n50756) );
  NAND2X1 U53088 ( .A(n50757), .B(n50756), .Y(u_decode_u_regfile_N917) );
  NOR2X1 U53089 ( .A(n44502), .B(n43075), .Y(n50759) );
  NOR2X1 U53090 ( .A(n44499), .B(n43078), .Y(n50758) );
  NOR2X1 U53091 ( .A(n50759), .B(n50758), .Y(n50761) );
  NOR2X1 U53092 ( .A(n20438), .B(n20437), .Y(n50760) );
  NAND2X1 U53093 ( .A(n50761), .B(n50760), .Y(u_decode_u_regfile_N547) );
  NOR2X1 U53094 ( .A(n44340), .B(n43075), .Y(n50763) );
  NOR2X1 U53095 ( .A(n44337), .B(n43078), .Y(n50762) );
  NOR2X1 U53096 ( .A(n50763), .B(n50762), .Y(n50765) );
  NOR2X1 U53097 ( .A(n23296), .B(n23295), .Y(n50764) );
  NAND2X1 U53098 ( .A(n50765), .B(n50764), .Y(u_decode_u_regfile_N1139) );
  NOR2X1 U53099 ( .A(n44352), .B(n43075), .Y(n50767) );
  NOR2X1 U53100 ( .A(n44349), .B(n43078), .Y(n50766) );
  NOR2X1 U53101 ( .A(n50767), .B(n50766), .Y(n50769) );
  NOR2X1 U53102 ( .A(n23076), .B(n23075), .Y(n50768) );
  NAND2X1 U53103 ( .A(n50769), .B(n50768), .Y(u_decode_u_regfile_N1176) );
  NOR2X1 U53104 ( .A(n44577), .B(n43075), .Y(n50771) );
  NOR2X1 U53105 ( .A(n44574), .B(n43078), .Y(n50770) );
  NOR2X1 U53106 ( .A(n50771), .B(n50770), .Y(n50773) );
  NOR2X1 U53107 ( .A(n18866), .B(n18865), .Y(n50772) );
  NAND2X1 U53108 ( .A(n50773), .B(n50772), .Y(u_decode_u_regfile_N843) );
  NOR2X1 U53109 ( .A(n44526), .B(n43075), .Y(n50775) );
  NOR2X1 U53110 ( .A(n44523), .B(n43077), .Y(n50774) );
  NOR2X1 U53111 ( .A(n50775), .B(n50774), .Y(n50777) );
  NOR2X1 U53112 ( .A(n20046), .B(n20045), .Y(n50776) );
  NAND2X1 U53113 ( .A(n50777), .B(n50776), .Y(u_decode_u_regfile_N621) );
  NOR2X1 U53114 ( .A(n44514), .B(n43074), .Y(n50779) );
  NOR2X1 U53115 ( .A(n44511), .B(n43077), .Y(n50778) );
  NOR2X1 U53116 ( .A(n50779), .B(n50778), .Y(n50781) );
  NOR2X1 U53117 ( .A(n20242), .B(n20241), .Y(n50780) );
  NAND2X1 U53118 ( .A(n50781), .B(n50780), .Y(u_decode_u_regfile_N584) );
  INVX1 U53119 ( .A(n58156), .Y(n50782) );
  NAND2X1 U53120 ( .A(n50782), .B(n43383), .Y(n57209) );
  NOR2X1 U53121 ( .A(n43074), .B(n43276), .Y(n50784) );
  NOR2X1 U53122 ( .A(n43077), .B(n43383), .Y(n50783) );
  NOR2X1 U53123 ( .A(n50784), .B(n50783), .Y(n50786) );
  NOR2X1 U53124 ( .A(n20634), .B(n20633), .Y(n50785) );
  NAND2X1 U53125 ( .A(n50786), .B(n50785), .Y(u_decode_u_regfile_N510) );
  INVX1 U53126 ( .A(n50792), .Y(n50831) );
  NAND2X1 U53127 ( .A(writeback_exec_idx_w[3]), .B(n50831), .Y(n50837) );
  INVX1 U53128 ( .A(n50837), .Y(n50825) );
  NOR2X1 U53129 ( .A(n44460), .B(n43074), .Y(n50788) );
  NOR2X1 U53130 ( .A(n44457), .B(n43077), .Y(n50787) );
  NOR2X1 U53131 ( .A(n50788), .B(n50787), .Y(n50790) );
  NOR2X1 U53132 ( .A(n21222), .B(n21221), .Y(n50789) );
  NAND2X1 U53133 ( .A(n50790), .B(n50789), .Y(u_decode_u_regfile_N399) );
  NOR2X1 U53134 ( .A(n50792), .B(n50791), .Y(n50793) );
  NOR2X1 U53135 ( .A(n19678), .B(n43074), .Y(n50795) );
  NOR2X1 U53136 ( .A(n44535), .B(n43077), .Y(n50794) );
  NOR2X1 U53137 ( .A(n50795), .B(n50794), .Y(n50797) );
  NOR2X1 U53138 ( .A(n19849), .B(n19848), .Y(n50796) );
  NAND2X1 U53139 ( .A(n50797), .B(n50796), .Y(u_decode_u_regfile_N658) );
  NOR2X1 U53140 ( .A(n44550), .B(n43075), .Y(n50799) );
  NOR2X1 U53141 ( .A(n44547), .B(n43077), .Y(n50798) );
  NOR2X1 U53142 ( .A(n50799), .B(n50798), .Y(n50801) );
  NOR2X1 U53143 ( .A(n19652), .B(n19651), .Y(n50800) );
  NAND2X1 U53144 ( .A(n50801), .B(n50800), .Y(u_decode_u_regfile_N695) );
  NOR2X1 U53145 ( .A(n44565), .B(n43074), .Y(n50804) );
  NOR2X1 U53146 ( .A(n44562), .B(n43077), .Y(n50803) );
  NOR2X1 U53147 ( .A(n50804), .B(n50803), .Y(n50806) );
  NOR2X1 U53148 ( .A(n19258), .B(n19257), .Y(n50805) );
  NAND2X1 U53149 ( .A(n50806), .B(n50805), .Y(u_decode_u_regfile_N769) );
  NOR2X1 U53150 ( .A(n44394), .B(n43074), .Y(n50808) );
  NOR2X1 U53151 ( .A(n44391), .B(n43078), .Y(n50807) );
  NOR2X1 U53152 ( .A(n50808), .B(n50807), .Y(n50810) );
  NOR2X1 U53153 ( .A(n22400), .B(n22399), .Y(n50809) );
  NAND2X1 U53154 ( .A(n50810), .B(n50809), .Y(u_decode_u_regfile_N177) );
  NOR2X1 U53155 ( .A(n44316), .B(n43074), .Y(n50812) );
  NOR2X1 U53156 ( .A(n44313), .B(n43077), .Y(n50811) );
  NOR2X1 U53157 ( .A(n50812), .B(n50811), .Y(n50814) );
  NOR2X1 U53158 ( .A(n23730), .B(n23729), .Y(n50813) );
  NAND2X1 U53159 ( .A(n50814), .B(n50813), .Y(u_decode_u_regfile_N1065) );
  NOR2X1 U53160 ( .A(n44484), .B(n43074), .Y(n50816) );
  NOR2X1 U53161 ( .A(n44481), .B(n43077), .Y(n50815) );
  NOR2X1 U53162 ( .A(n50816), .B(n50815), .Y(n50818) );
  NOR2X1 U53163 ( .A(n20830), .B(n20829), .Y(n50817) );
  NAND2X1 U53164 ( .A(n50818), .B(n50817), .Y(u_decode_u_regfile_N473) );
  NOR2X1 U53165 ( .A(n50838), .B(n50837), .Y(n50819) );
  NOR2X1 U53166 ( .A(n44601), .B(n43074), .Y(n50821) );
  NOR2X1 U53167 ( .A(n44598), .B(n43077), .Y(n50820) );
  NOR2X1 U53168 ( .A(n50821), .B(n50820), .Y(n50823) );
  NOR2X1 U53169 ( .A(n18277), .B(n18276), .Y(n50822) );
  NAND2X1 U53170 ( .A(n50823), .B(n50822), .Y(u_decode_u_regfile_N954) );
  NOR2X1 U53171 ( .A(n50838), .B(n50824), .Y(n50826) );
  NOR2X1 U53172 ( .A(n44607), .B(n43074), .Y(n50828) );
  NOR2X1 U53173 ( .A(n44604), .B(n43077), .Y(n50827) );
  NOR2X1 U53174 ( .A(n50828), .B(n50827), .Y(n50830) );
  NOR2X1 U53175 ( .A(n18060), .B(n18058), .Y(n50829) );
  NAND2X1 U53176 ( .A(n50830), .B(n50829), .Y(u_decode_u_regfile_N991) );
  NAND2X1 U53177 ( .A(n40841), .B(n35922), .Y(n24109) );
  INVX1 U53178 ( .A(n24109), .Y(n50832) );
  NAND2X1 U53179 ( .A(n43389), .B(n50832), .Y(n57144) );
  NOR2X1 U53180 ( .A(n43074), .B(n43273), .Y(n50834) );
  NOR2X1 U53181 ( .A(n43077), .B(n43389), .Y(n50833) );
  NOR2X1 U53182 ( .A(n50834), .B(n50833), .Y(n50836) );
  NOR2X1 U53183 ( .A(n23938), .B(n23937), .Y(n50835) );
  NAND2X1 U53184 ( .A(n50836), .B(n50835), .Y(u_decode_u_regfile_N103) );
  NAND2X1 U53185 ( .A(n57515), .B(n35922), .Y(n21437) );
  INVX1 U53186 ( .A(n21437), .Y(n50839) );
  NAND2X1 U53187 ( .A(n43386), .B(n50839), .Y(n57131) );
  NOR2X1 U53188 ( .A(n43074), .B(n43270), .Y(n50841) );
  NOR2X1 U53189 ( .A(n43077), .B(n43386), .Y(n50840) );
  NOR2X1 U53190 ( .A(n50841), .B(n50840), .Y(n50843) );
  NOR2X1 U53191 ( .A(n21419), .B(n21418), .Y(n50842) );
  NAND2X1 U53192 ( .A(n50843), .B(n50842), .Y(u_decode_u_regfile_N362) );
  NAND2X1 U53193 ( .A(n43408), .B(n43804), .Y(n50848) );
  NAND2X1 U53194 ( .A(n43412), .B(n50844), .Y(n58548) );
  NAND2X1 U53195 ( .A(n57099), .B(n50845), .Y(n50846) );
  NAND2X1 U53196 ( .A(n58548), .B(n50846), .Y(n56831) );
  NAND2X1 U53197 ( .A(n40454), .B(n56831), .Y(n50847) );
  NAND2X1 U53198 ( .A(n50848), .B(n50847), .Y(n15742) );
  NAND2X1 U53199 ( .A(n17937), .B(n58540), .Y(n50849) );
  NAND2X1 U53200 ( .A(n57094), .B(n50849), .Y(n50853) );
  NOR2X1 U53201 ( .A(opcode_instr_w[11]), .B(n50859), .Y(n50851) );
  NAND2X1 U53202 ( .A(n50851), .B(n50850), .Y(n50852) );
  AND2X1 U53203 ( .A(n50853), .B(n50852), .Y(n50855) );
  NAND2X1 U53204 ( .A(n57094), .B(n50854), .Y(n57089) );
  NAND2X1 U53205 ( .A(n50855), .B(n57089), .Y(n57333) );
  NAND2X1 U53206 ( .A(n42939), .B(n50856), .Y(n50857) );
  NOR2X1 U53207 ( .A(opcode_instr_w_17), .B(n50857), .Y(n50865) );
  NAND2X1 U53208 ( .A(n42609), .B(n50859), .Y(n50861) );
  NAND2X1 U53209 ( .A(opcode_instr_w[12]), .B(n8955), .Y(n50860) );
  NOR2X1 U53210 ( .A(n50861), .B(n50860), .Y(n50863) );
  NOR2X1 U53211 ( .A(n42434), .B(n43410), .Y(n50862) );
  NOR2X1 U53212 ( .A(n50863), .B(n50862), .Y(n50864) );
  NAND2X1 U53213 ( .A(n50865), .B(n50864), .Y(n58543) );
  NOR2X1 U53214 ( .A(n57333), .B(n58543), .Y(n50866) );
  NAND2X1 U53215 ( .A(n42455), .B(n15742), .Y(n15594) );
  NOR2X1 U53216 ( .A(n44364), .B(n43451), .Y(n50868) );
  NOR2X1 U53217 ( .A(n44361), .B(n43335), .Y(n50867) );
  NOR2X1 U53218 ( .A(n50868), .B(n50867), .Y(n50870) );
  NOR2X1 U53219 ( .A(n22874), .B(n22873), .Y(n50869) );
  NAND2X1 U53220 ( .A(n50870), .B(n50869), .Y(u_decode_u_regfile_N1210) );
  NOR2X1 U53221 ( .A(n44442), .B(n43453), .Y(n50872) );
  NOR2X1 U53222 ( .A(n44439), .B(n37665), .Y(n50871) );
  NOR2X1 U53223 ( .A(n50872), .B(n50871), .Y(n50874) );
  NOR2X1 U53224 ( .A(n21634), .B(n21633), .Y(n50873) );
  NAND2X1 U53225 ( .A(n50874), .B(n50873), .Y(u_decode_u_regfile_N322) );
  NOR2X1 U53226 ( .A(n44382), .B(n43453), .Y(n50876) );
  NOR2X1 U53227 ( .A(n44379), .B(n37665), .Y(n50875) );
  NOR2X1 U53228 ( .A(n50876), .B(n50875), .Y(n50878) );
  NOR2X1 U53229 ( .A(n22614), .B(n22613), .Y(n50877) );
  NAND2X1 U53230 ( .A(n50878), .B(n50877), .Y(u_decode_u_regfile_N137) );
  NOR2X1 U53231 ( .A(n44304), .B(n43453), .Y(n50880) );
  NOR2X1 U53232 ( .A(n44301), .B(n37665), .Y(n50879) );
  NOR2X1 U53233 ( .A(n50880), .B(n50879), .Y(n50882) );
  NOR2X1 U53234 ( .A(n23968), .B(n23967), .Y(n50881) );
  NAND2X1 U53235 ( .A(n50882), .B(n50881), .Y(u_decode_u_regfile_N1025) );
  NOR2X1 U53236 ( .A(n44406), .B(n43453), .Y(n50884) );
  NOR2X1 U53237 ( .A(n44403), .B(n43336), .Y(n50883) );
  NOR2X1 U53238 ( .A(n50884), .B(n50883), .Y(n50886) );
  NOR2X1 U53239 ( .A(n22222), .B(n22221), .Y(n50885) );
  NAND2X1 U53240 ( .A(n50886), .B(n50885), .Y(u_decode_u_regfile_N211) );
  NOR2X1 U53241 ( .A(n44559), .B(n43452), .Y(n50888) );
  NOR2X1 U53242 ( .A(n44556), .B(n43336), .Y(n50887) );
  NOR2X1 U53243 ( .A(n50888), .B(n50887), .Y(n50890) );
  NOR2X1 U53244 ( .A(n19473), .B(n19471), .Y(n50889) );
  NAND2X1 U53245 ( .A(n50890), .B(n50889), .Y(u_decode_u_regfile_N729) );
  NOR2X1 U53246 ( .A(n44328), .B(n43452), .Y(n50892) );
  NOR2X1 U53247 ( .A(n44325), .B(n43336), .Y(n50891) );
  NOR2X1 U53248 ( .A(n50892), .B(n50891), .Y(n50894) );
  NOR2X1 U53249 ( .A(n23534), .B(n23533), .Y(n50893) );
  NAND2X1 U53250 ( .A(n50894), .B(n50893), .Y(u_decode_u_regfile_N1099) );
  NOR2X1 U53251 ( .A(n44430), .B(n43452), .Y(n50896) );
  NOR2X1 U53252 ( .A(n44427), .B(n43336), .Y(n50895) );
  NOR2X1 U53253 ( .A(n50896), .B(n50895), .Y(n50898) );
  NOR2X1 U53254 ( .A(n21830), .B(n21829), .Y(n50897) );
  NAND2X1 U53255 ( .A(n50898), .B(n50897), .Y(u_decode_u_regfile_N285) );
  NOR2X1 U53256 ( .A(n44418), .B(n43452), .Y(n50900) );
  NOR2X1 U53257 ( .A(n44415), .B(n43336), .Y(n50899) );
  NOR2X1 U53258 ( .A(n50900), .B(n50899), .Y(n50902) );
  NOR2X1 U53259 ( .A(n22026), .B(n22025), .Y(n50901) );
  NAND2X1 U53260 ( .A(n50902), .B(n50901), .Y(u_decode_u_regfile_N248) );
  NOR2X1 U53261 ( .A(n44472), .B(n43452), .Y(n50904) );
  NOR2X1 U53262 ( .A(n44469), .B(n43336), .Y(n50903) );
  NOR2X1 U53263 ( .A(n50904), .B(n50903), .Y(n50906) );
  NOR2X1 U53264 ( .A(n21044), .B(n21043), .Y(n50905) );
  NAND2X1 U53265 ( .A(n50906), .B(n50905), .Y(u_decode_u_regfile_N433) );
  NOR2X1 U53266 ( .A(n44583), .B(n43452), .Y(n50908) );
  NOR2X1 U53267 ( .A(n44580), .B(n43336), .Y(n50907) );
  NOR2X1 U53268 ( .A(n50908), .B(n50907), .Y(n50910) );
  NOR2X1 U53269 ( .A(n18689), .B(n18687), .Y(n50909) );
  NAND2X1 U53270 ( .A(n50910), .B(n50909), .Y(u_decode_u_regfile_N877) );
  NOR2X1 U53271 ( .A(n44571), .B(n43452), .Y(n50912) );
  NOR2X1 U53272 ( .A(n44568), .B(n43336), .Y(n50911) );
  NOR2X1 U53273 ( .A(n50912), .B(n50911), .Y(n50914) );
  NOR2X1 U53274 ( .A(n19081), .B(n19079), .Y(n50913) );
  NAND2X1 U53275 ( .A(n50914), .B(n50913), .Y(u_decode_u_regfile_N803) );
  NOR2X1 U53276 ( .A(n44592), .B(n43452), .Y(n50916) );
  NOR2X1 U53277 ( .A(n44589), .B(n43336), .Y(n50915) );
  NOR2X1 U53278 ( .A(n50916), .B(n50915), .Y(n50918) );
  NOR2X1 U53279 ( .A(n18494), .B(n18493), .Y(n50917) );
  NAND2X1 U53280 ( .A(n50918), .B(n50917), .Y(u_decode_u_regfile_N914) );
  NOR2X1 U53281 ( .A(n44502), .B(n43452), .Y(n50920) );
  NOR2X1 U53282 ( .A(n44499), .B(n43336), .Y(n50919) );
  NOR2X1 U53283 ( .A(n50920), .B(n50919), .Y(n50922) );
  NOR2X1 U53284 ( .A(n20456), .B(n20455), .Y(n50921) );
  NAND2X1 U53285 ( .A(n50922), .B(n50921), .Y(u_decode_u_regfile_N544) );
  NOR2X1 U53286 ( .A(n44340), .B(n43452), .Y(n50924) );
  NOR2X1 U53287 ( .A(n44337), .B(n43336), .Y(n50923) );
  NOR2X1 U53288 ( .A(n50924), .B(n50923), .Y(n50926) );
  NOR2X1 U53289 ( .A(n23314), .B(n23313), .Y(n50925) );
  NAND2X1 U53290 ( .A(n50926), .B(n50925), .Y(u_decode_u_regfile_N1136) );
  NOR2X1 U53291 ( .A(n44352), .B(n43452), .Y(n50928) );
  NOR2X1 U53292 ( .A(n44349), .B(n43336), .Y(n50927) );
  NOR2X1 U53293 ( .A(n50928), .B(n50927), .Y(n50930) );
  NOR2X1 U53294 ( .A(n23094), .B(n23093), .Y(n50929) );
  NAND2X1 U53295 ( .A(n50930), .B(n50929), .Y(u_decode_u_regfile_N1173) );
  NOR2X1 U53296 ( .A(n44577), .B(n43452), .Y(n50932) );
  NOR2X1 U53297 ( .A(n44574), .B(n43336), .Y(n50931) );
  NOR2X1 U53298 ( .A(n50932), .B(n50931), .Y(n50934) );
  NOR2X1 U53299 ( .A(n18885), .B(n18883), .Y(n50933) );
  NAND2X1 U53300 ( .A(n50934), .B(n50933), .Y(u_decode_u_regfile_N840) );
  NOR2X1 U53301 ( .A(n44526), .B(n43452), .Y(n50936) );
  NOR2X1 U53302 ( .A(n44523), .B(n43335), .Y(n50935) );
  NOR2X1 U53303 ( .A(n50936), .B(n50935), .Y(n50938) );
  NOR2X1 U53304 ( .A(n20064), .B(n20063), .Y(n50937) );
  NAND2X1 U53305 ( .A(n50938), .B(n50937), .Y(u_decode_u_regfile_N618) );
  NOR2X1 U53306 ( .A(n44514), .B(n43451), .Y(n50940) );
  NOR2X1 U53307 ( .A(n44511), .B(n43335), .Y(n50939) );
  NOR2X1 U53308 ( .A(n50940), .B(n50939), .Y(n50942) );
  NOR2X1 U53309 ( .A(n20260), .B(n20259), .Y(n50941) );
  NAND2X1 U53310 ( .A(n50942), .B(n50941), .Y(u_decode_u_regfile_N581) );
  NOR2X1 U53311 ( .A(n43451), .B(n43276), .Y(n50944) );
  NOR2X1 U53312 ( .A(n43335), .B(n43385), .Y(n50943) );
  NOR2X1 U53313 ( .A(n50944), .B(n50943), .Y(n50946) );
  NOR2X1 U53314 ( .A(n20652), .B(n20651), .Y(n50945) );
  NAND2X1 U53315 ( .A(n50946), .B(n50945), .Y(u_decode_u_regfile_N507) );
  NOR2X1 U53316 ( .A(n44460), .B(n43451), .Y(n50948) );
  NOR2X1 U53317 ( .A(n44457), .B(n43335), .Y(n50947) );
  NOR2X1 U53318 ( .A(n50948), .B(n50947), .Y(n50950) );
  NOR2X1 U53319 ( .A(n21241), .B(n21239), .Y(n50949) );
  NAND2X1 U53320 ( .A(n50950), .B(n50949), .Y(u_decode_u_regfile_N396) );
  NOR2X1 U53321 ( .A(n19678), .B(n43451), .Y(n50952) );
  NOR2X1 U53322 ( .A(n44535), .B(n43335), .Y(n50951) );
  NOR2X1 U53323 ( .A(n50952), .B(n50951), .Y(n50954) );
  NOR2X1 U53324 ( .A(n19868), .B(n19866), .Y(n50953) );
  NAND2X1 U53325 ( .A(n50954), .B(n50953), .Y(u_decode_u_regfile_N655) );
  NOR2X1 U53326 ( .A(n44550), .B(n43451), .Y(n50956) );
  NOR2X1 U53327 ( .A(n44547), .B(n43335), .Y(n50955) );
  NOR2X1 U53328 ( .A(n50956), .B(n50955), .Y(n50958) );
  NOR2X1 U53329 ( .A(n19671), .B(n19669), .Y(n50957) );
  NAND2X1 U53330 ( .A(n50958), .B(n50957), .Y(u_decode_u_regfile_N692) );
  NOR2X1 U53331 ( .A(n44565), .B(n43452), .Y(n50960) );
  NOR2X1 U53332 ( .A(n44562), .B(n43335), .Y(n50959) );
  NOR2X1 U53333 ( .A(n50960), .B(n50959), .Y(n50962) );
  NOR2X1 U53334 ( .A(n19277), .B(n19275), .Y(n50961) );
  NAND2X1 U53335 ( .A(n50962), .B(n50961), .Y(u_decode_u_regfile_N766) );
  NOR2X1 U53336 ( .A(n44394), .B(n43451), .Y(n50964) );
  NOR2X1 U53337 ( .A(n44391), .B(n43335), .Y(n50963) );
  NOR2X1 U53338 ( .A(n50964), .B(n50963), .Y(n50966) );
  NOR2X1 U53339 ( .A(n22418), .B(n22417), .Y(n50965) );
  NAND2X1 U53340 ( .A(n50966), .B(n50965), .Y(u_decode_u_regfile_N174) );
  NOR2X1 U53341 ( .A(n44316), .B(n43451), .Y(n50968) );
  NOR2X1 U53342 ( .A(n44313), .B(n43335), .Y(n50967) );
  NOR2X1 U53343 ( .A(n50968), .B(n50967), .Y(n50970) );
  NOR2X1 U53344 ( .A(n23748), .B(n23747), .Y(n50969) );
  NAND2X1 U53345 ( .A(n50970), .B(n50969), .Y(u_decode_u_regfile_N1062) );
  NOR2X1 U53346 ( .A(n44484), .B(n43451), .Y(n50972) );
  NOR2X1 U53347 ( .A(n44481), .B(n43335), .Y(n50971) );
  NOR2X1 U53348 ( .A(n50972), .B(n50971), .Y(n50974) );
  NOR2X1 U53349 ( .A(n20848), .B(n20847), .Y(n50973) );
  NAND2X1 U53350 ( .A(n50974), .B(n50973), .Y(u_decode_u_regfile_N470) );
  NOR2X1 U53351 ( .A(n44601), .B(n43451), .Y(n50976) );
  NOR2X1 U53352 ( .A(n44598), .B(n43335), .Y(n50975) );
  NOR2X1 U53353 ( .A(n50976), .B(n50975), .Y(n50978) );
  NOR2X1 U53354 ( .A(n18297), .B(n18294), .Y(n50977) );
  NAND2X1 U53355 ( .A(n50978), .B(n50977), .Y(u_decode_u_regfile_N951) );
  NOR2X1 U53356 ( .A(n43451), .B(n43273), .Y(n50980) );
  NOR2X1 U53357 ( .A(n43335), .B(n43391), .Y(n50979) );
  NOR2X1 U53358 ( .A(n50980), .B(n50979), .Y(n50982) );
  NOR2X1 U53359 ( .A(n24110), .B(n24108), .Y(n50981) );
  NAND2X1 U53360 ( .A(n50982), .B(n50981), .Y(u_decode_u_regfile_N100) );
  NOR2X1 U53361 ( .A(n43451), .B(n43270), .Y(n50984) );
  NOR2X1 U53362 ( .A(n43335), .B(n43388), .Y(n50983) );
  NOR2X1 U53363 ( .A(n50984), .B(n50983), .Y(n50986) );
  NOR2X1 U53364 ( .A(n21438), .B(n21436), .Y(n50985) );
  NAND2X1 U53365 ( .A(n50986), .B(n50985), .Y(u_decode_u_regfile_N359) );
  NOR2X1 U53366 ( .A(n16582), .B(n16583), .Y(n50988) );
  NOR2X1 U53367 ( .A(n16616), .B(n16617), .Y(n50987) );
  NAND2X1 U53368 ( .A(n50988), .B(n50987), .Y(u_exec_alu_p_w[1]) );
  NOR2X1 U53369 ( .A(n44364), .B(n43080), .Y(n50990) );
  NOR2X1 U53370 ( .A(n44361), .B(n43083), .Y(n50989) );
  NOR2X1 U53371 ( .A(n50990), .B(n50989), .Y(n50992) );
  NOR2X1 U53372 ( .A(n22868), .B(n22867), .Y(n50991) );
  NAND2X1 U53373 ( .A(n50992), .B(n50991), .Y(u_decode_u_regfile_N1211) );
  NOR2X1 U53374 ( .A(n44340), .B(n43082), .Y(n50994) );
  NOR2X1 U53375 ( .A(n44337), .B(n37666), .Y(n50993) );
  NOR2X1 U53376 ( .A(n50994), .B(n50993), .Y(n50996) );
  NOR2X1 U53377 ( .A(n23308), .B(n23307), .Y(n50995) );
  NAND2X1 U53378 ( .A(n50996), .B(n50995), .Y(u_decode_u_regfile_N1137) );
  NOR2X1 U53379 ( .A(n44352), .B(n43082), .Y(n50998) );
  NOR2X1 U53380 ( .A(n44349), .B(n37666), .Y(n50997) );
  NOR2X1 U53381 ( .A(n50998), .B(n50997), .Y(n51000) );
  NOR2X1 U53382 ( .A(n23088), .B(n23087), .Y(n50999) );
  NAND2X1 U53383 ( .A(n51000), .B(n50999), .Y(u_decode_u_regfile_N1174) );
  NOR2X1 U53384 ( .A(n44304), .B(n43082), .Y(n51002) );
  NOR2X1 U53385 ( .A(n44301), .B(n37666), .Y(n51001) );
  NOR2X1 U53386 ( .A(n51002), .B(n51001), .Y(n51004) );
  NOR2X1 U53387 ( .A(n23962), .B(n23961), .Y(n51003) );
  NAND2X1 U53388 ( .A(n51004), .B(n51003), .Y(u_decode_u_regfile_N1026) );
  NOR2X1 U53389 ( .A(n44328), .B(n43082), .Y(n51006) );
  NOR2X1 U53390 ( .A(n44325), .B(n43084), .Y(n51005) );
  NOR2X1 U53391 ( .A(n51006), .B(n51005), .Y(n51008) );
  NOR2X1 U53392 ( .A(n23522), .B(n23521), .Y(n51007) );
  NAND2X1 U53393 ( .A(n51008), .B(n51007), .Y(u_decode_u_regfile_N1100) );
  NOR2X1 U53394 ( .A(n44583), .B(n43081), .Y(n51010) );
  NOR2X1 U53395 ( .A(n44580), .B(n43084), .Y(n51009) );
  NOR2X1 U53396 ( .A(n51010), .B(n51009), .Y(n51012) );
  NOR2X1 U53397 ( .A(n18682), .B(n18681), .Y(n51011) );
  NAND2X1 U53398 ( .A(n51012), .B(n51011), .Y(u_decode_u_regfile_N878) );
  NOR2X1 U53399 ( .A(n44592), .B(n43081), .Y(n51014) );
  NOR2X1 U53400 ( .A(n44589), .B(n43084), .Y(n51013) );
  NOR2X1 U53401 ( .A(n51014), .B(n51013), .Y(n51016) );
  NOR2X1 U53402 ( .A(n18488), .B(n18487), .Y(n51015) );
  NAND2X1 U53403 ( .A(n51016), .B(n51015), .Y(u_decode_u_regfile_N915) );
  NOR2X1 U53404 ( .A(n44577), .B(n43081), .Y(n51018) );
  NOR2X1 U53405 ( .A(n44574), .B(n43084), .Y(n51017) );
  NOR2X1 U53406 ( .A(n51018), .B(n51017), .Y(n51020) );
  NOR2X1 U53407 ( .A(n18878), .B(n18877), .Y(n51019) );
  NAND2X1 U53408 ( .A(n51020), .B(n51019), .Y(u_decode_u_regfile_N841) );
  NOR2X1 U53409 ( .A(n44559), .B(n43081), .Y(n51022) );
  NOR2X1 U53410 ( .A(n44556), .B(n43084), .Y(n51021) );
  NOR2X1 U53411 ( .A(n51022), .B(n51021), .Y(n51024) );
  NOR2X1 U53412 ( .A(n19466), .B(n19465), .Y(n51023) );
  NAND2X1 U53413 ( .A(n51024), .B(n51023), .Y(u_decode_u_regfile_N730) );
  NOR2X1 U53414 ( .A(n44571), .B(n43081), .Y(n51026) );
  NOR2X1 U53415 ( .A(n44568), .B(n43084), .Y(n51025) );
  NOR2X1 U53416 ( .A(n51026), .B(n51025), .Y(n51028) );
  NOR2X1 U53417 ( .A(n19074), .B(n19073), .Y(n51027) );
  NAND2X1 U53418 ( .A(n51028), .B(n51027), .Y(u_decode_u_regfile_N804) );
  NOR2X1 U53419 ( .A(n44502), .B(n43081), .Y(n51030) );
  NOR2X1 U53420 ( .A(n44499), .B(n43084), .Y(n51029) );
  NOR2X1 U53421 ( .A(n51030), .B(n51029), .Y(n51032) );
  NOR2X1 U53422 ( .A(n20450), .B(n20449), .Y(n51031) );
  NAND2X1 U53423 ( .A(n51032), .B(n51031), .Y(u_decode_u_regfile_N545) );
  NOR2X1 U53424 ( .A(n44526), .B(n43081), .Y(n51034) );
  NOR2X1 U53425 ( .A(n44523), .B(n43084), .Y(n51033) );
  NOR2X1 U53426 ( .A(n51034), .B(n51033), .Y(n51036) );
  NOR2X1 U53427 ( .A(n20058), .B(n20057), .Y(n51035) );
  NAND2X1 U53428 ( .A(n51036), .B(n51035), .Y(u_decode_u_regfile_N619) );
  NOR2X1 U53429 ( .A(n44514), .B(n43081), .Y(n51038) );
  NOR2X1 U53430 ( .A(n44511), .B(n43084), .Y(n51037) );
  NOR2X1 U53431 ( .A(n51038), .B(n51037), .Y(n51040) );
  NOR2X1 U53432 ( .A(n20254), .B(n20253), .Y(n51039) );
  NAND2X1 U53433 ( .A(n51040), .B(n51039), .Y(u_decode_u_regfile_N582) );
  NOR2X1 U53434 ( .A(n44472), .B(n43081), .Y(n51042) );
  NOR2X1 U53435 ( .A(n44469), .B(n43084), .Y(n51041) );
  NOR2X1 U53436 ( .A(n51042), .B(n51041), .Y(n51044) );
  NOR2X1 U53437 ( .A(n21038), .B(n21037), .Y(n51043) );
  NAND2X1 U53438 ( .A(n51044), .B(n51043), .Y(u_decode_u_regfile_N434) );
  NOR2X1 U53439 ( .A(n43080), .B(n43276), .Y(n51046) );
  NOR2X1 U53440 ( .A(n43083), .B(n43385), .Y(n51045) );
  NOR2X1 U53441 ( .A(n51046), .B(n51045), .Y(n51048) );
  NOR2X1 U53442 ( .A(n20646), .B(n20645), .Y(n51047) );
  NAND2X1 U53443 ( .A(n51048), .B(n51047), .Y(u_decode_u_regfile_N508) );
  NOR2X1 U53444 ( .A(n44442), .B(n43081), .Y(n51050) );
  NOR2X1 U53445 ( .A(n44439), .B(n43084), .Y(n51049) );
  NOR2X1 U53446 ( .A(n51050), .B(n51049), .Y(n51052) );
  NOR2X1 U53447 ( .A(n21628), .B(n21627), .Y(n51051) );
  NAND2X1 U53448 ( .A(n51052), .B(n51051), .Y(u_decode_u_regfile_N323) );
  NOR2X1 U53449 ( .A(n44430), .B(n43081), .Y(n51054) );
  NOR2X1 U53450 ( .A(n44427), .B(n43084), .Y(n51053) );
  NOR2X1 U53451 ( .A(n51054), .B(n51053), .Y(n51056) );
  NOR2X1 U53452 ( .A(n21824), .B(n21823), .Y(n51055) );
  NAND2X1 U53453 ( .A(n51056), .B(n51055), .Y(u_decode_u_regfile_N286) );
  NOR2X1 U53454 ( .A(n44418), .B(n43081), .Y(n51058) );
  NOR2X1 U53455 ( .A(n44415), .B(n43084), .Y(n51057) );
  NOR2X1 U53456 ( .A(n51058), .B(n51057), .Y(n51060) );
  NOR2X1 U53457 ( .A(n22020), .B(n22019), .Y(n51059) );
  NAND2X1 U53458 ( .A(n51060), .B(n51059), .Y(u_decode_u_regfile_N249) );
  NOR2X1 U53459 ( .A(n44382), .B(n43081), .Y(n51062) );
  NOR2X1 U53460 ( .A(n44379), .B(n43083), .Y(n51061) );
  NOR2X1 U53461 ( .A(n51062), .B(n51061), .Y(n51064) );
  NOR2X1 U53462 ( .A(n22608), .B(n22607), .Y(n51063) );
  NAND2X1 U53463 ( .A(n51064), .B(n51063), .Y(u_decode_u_regfile_N138) );
  NOR2X1 U53464 ( .A(n44406), .B(n43080), .Y(n51066) );
  NOR2X1 U53465 ( .A(n44403), .B(n43083), .Y(n51065) );
  NOR2X1 U53466 ( .A(n51066), .B(n51065), .Y(n51068) );
  NOR2X1 U53467 ( .A(n22216), .B(n22215), .Y(n51067) );
  NAND2X1 U53468 ( .A(n51068), .B(n51067), .Y(u_decode_u_regfile_N212) );
  NOR2X1 U53469 ( .A(n44460), .B(n43080), .Y(n51070) );
  NOR2X1 U53470 ( .A(n44457), .B(n43083), .Y(n51069) );
  NOR2X1 U53471 ( .A(n51070), .B(n51069), .Y(n51072) );
  NOR2X1 U53472 ( .A(n21234), .B(n21233), .Y(n51071) );
  NAND2X1 U53473 ( .A(n51072), .B(n51071), .Y(u_decode_u_regfile_N397) );
  NOR2X1 U53474 ( .A(n44539), .B(n43080), .Y(n51074) );
  NOR2X1 U53475 ( .A(n44535), .B(n43083), .Y(n51073) );
  NOR2X1 U53476 ( .A(n51074), .B(n51073), .Y(n51076) );
  NOR2X1 U53477 ( .A(n19861), .B(n19860), .Y(n51075) );
  NAND2X1 U53478 ( .A(n51076), .B(n51075), .Y(u_decode_u_regfile_N656) );
  NOR2X1 U53479 ( .A(n44550), .B(n43081), .Y(n51078) );
  NOR2X1 U53480 ( .A(n44547), .B(n43083), .Y(n51077) );
  NOR2X1 U53481 ( .A(n51078), .B(n51077), .Y(n51080) );
  NOR2X1 U53482 ( .A(n19664), .B(n19663), .Y(n51079) );
  NAND2X1 U53483 ( .A(n51080), .B(n51079), .Y(u_decode_u_regfile_N693) );
  NOR2X1 U53484 ( .A(n44565), .B(n43080), .Y(n51082) );
  NOR2X1 U53485 ( .A(n44562), .B(n43083), .Y(n51081) );
  NOR2X1 U53486 ( .A(n51082), .B(n51081), .Y(n51084) );
  NOR2X1 U53487 ( .A(n19270), .B(n19269), .Y(n51083) );
  NAND2X1 U53488 ( .A(n51084), .B(n51083), .Y(u_decode_u_regfile_N767) );
  NOR2X1 U53489 ( .A(n44394), .B(n43080), .Y(n51086) );
  NOR2X1 U53490 ( .A(n44391), .B(n43084), .Y(n51085) );
  NOR2X1 U53491 ( .A(n51086), .B(n51085), .Y(n51088) );
  NOR2X1 U53492 ( .A(n22412), .B(n22411), .Y(n51087) );
  NAND2X1 U53493 ( .A(n51088), .B(n51087), .Y(u_decode_u_regfile_N175) );
  NOR2X1 U53494 ( .A(n44316), .B(n43080), .Y(n51090) );
  NOR2X1 U53495 ( .A(n44313), .B(n43083), .Y(n51089) );
  NOR2X1 U53496 ( .A(n51090), .B(n51089), .Y(n51092) );
  NOR2X1 U53497 ( .A(n23742), .B(n23741), .Y(n51091) );
  NAND2X1 U53498 ( .A(n51092), .B(n51091), .Y(u_decode_u_regfile_N1063) );
  NOR2X1 U53499 ( .A(n44484), .B(n43080), .Y(n51094) );
  NOR2X1 U53500 ( .A(n44481), .B(n43083), .Y(n51093) );
  NOR2X1 U53501 ( .A(n51094), .B(n51093), .Y(n51096) );
  NOR2X1 U53502 ( .A(n20842), .B(n20841), .Y(n51095) );
  NAND2X1 U53503 ( .A(n51096), .B(n51095), .Y(u_decode_u_regfile_N471) );
  NOR2X1 U53504 ( .A(n44601), .B(n43080), .Y(n51098) );
  NOR2X1 U53505 ( .A(n44598), .B(n43083), .Y(n51097) );
  NOR2X1 U53506 ( .A(n51098), .B(n51097), .Y(n51100) );
  NOR2X1 U53507 ( .A(n18289), .B(n18288), .Y(n51099) );
  NAND2X1 U53508 ( .A(n51100), .B(n51099), .Y(u_decode_u_regfile_N952) );
  NOR2X1 U53509 ( .A(n44607), .B(n43080), .Y(n51102) );
  NOR2X1 U53510 ( .A(n44604), .B(n43083), .Y(n51101) );
  NOR2X1 U53511 ( .A(n51102), .B(n51101), .Y(n51104) );
  NOR2X1 U53512 ( .A(n18074), .B(n18072), .Y(n51103) );
  NAND2X1 U53513 ( .A(n51104), .B(n51103), .Y(u_decode_u_regfile_N989) );
  NOR2X1 U53514 ( .A(n43080), .B(n43273), .Y(n51106) );
  NOR2X1 U53515 ( .A(n43083), .B(n43391), .Y(n51105) );
  NOR2X1 U53516 ( .A(n51106), .B(n51105), .Y(n51108) );
  NOR2X1 U53517 ( .A(n24040), .B(n24039), .Y(n51107) );
  NAND2X1 U53518 ( .A(n51108), .B(n51107), .Y(u_decode_u_regfile_N101) );
  NOR2X1 U53519 ( .A(n43080), .B(n43270), .Y(n51110) );
  NOR2X1 U53520 ( .A(n43083), .B(n43388), .Y(n51109) );
  NOR2X1 U53521 ( .A(n51110), .B(n51109), .Y(n51112) );
  NOR2X1 U53522 ( .A(n21431), .B(n21430), .Y(n51111) );
  NAND2X1 U53523 ( .A(n51112), .B(n51111), .Y(u_decode_u_regfile_N360) );
  NAND2X1 U53524 ( .A(n43410), .B(n43753), .Y(n51114) );
  NAND2X1 U53525 ( .A(n40453), .B(n56831), .Y(n51113) );
  NAND2X1 U53526 ( .A(n51114), .B(n51113), .Y(n16593) );
  OR2X1 U53527 ( .A(n57333), .B(n58544), .Y(n51115) );
  NOR2X1 U53528 ( .A(n58543), .B(n51115), .Y(n51411) );
  INVX1 U53529 ( .A(n15742), .Y(n73525) );
  INVX1 U53530 ( .A(n16635), .Y(n73571) );
  NAND2X1 U53531 ( .A(n42310), .B(n73571), .Y(n15465) );
  NAND2X1 U53532 ( .A(n43410), .B(n43732), .Y(n51117) );
  NAND2X1 U53533 ( .A(n39115), .B(n56831), .Y(n51116) );
  NAND2X1 U53534 ( .A(n51117), .B(n51116), .Y(n57316) );
  INVX1 U53535 ( .A(n57316), .Y(n57331) );
  INVX1 U53536 ( .A(n15465), .Y(n58576) );
  NAND2X1 U53537 ( .A(n43415), .B(n58576), .Y(n362) );
  NOR2X1 U53538 ( .A(n24422), .B(n57406), .Y(u_decode_N782) );
  NOR2X1 U53539 ( .A(n24422), .B(n57404), .Y(u_decode_N781) );
  NOR2X1 U53540 ( .A(n24422), .B(n57407), .Y(u_decode_N780) );
  NOR2X1 U53541 ( .A(opcode_instr_w_45), .B(opcode_instr_w_46), .Y(n51118) );
  NAND2X1 U53542 ( .A(n51118), .B(n55033), .Y(n58230) );
  INVX1 U53543 ( .A(n58230), .Y(n73522) );
  MX2X1 U53544 ( .A(n42731), .B(n36719), .S0(n73522), .Y(n26127) );
  NAND2X1 U53545 ( .A(n44281), .B(n26127), .Y(n26906) );
  INVX1 U53546 ( .A(n24469), .Y(n57592) );
  INVX1 U53547 ( .A(n24455), .Y(n57400) );
  NAND2X1 U53548 ( .A(n51119), .B(n57400), .Y(n51120) );
  NOR2X1 U53549 ( .A(n51121), .B(n51120), .Y(n51123) );
  NOR2X1 U53550 ( .A(n24474), .B(n51408), .Y(n51122) );
  NAND2X1 U53551 ( .A(n51123), .B(n51122), .Y(n57595) );
  OR2X1 U53552 ( .A(n42933), .B(n57595), .Y(n51124) );
  NOR2X1 U53553 ( .A(n57592), .B(n51124), .Y(u_decode_N792) );
  NAND2X1 U53554 ( .A(challenge[32]), .B(n44855), .Y(n51125) );
  NAND2X1 U53555 ( .A(n54381), .B(n51125), .Y(n17240) );
  NAND2X1 U53556 ( .A(opcode_instr_w_56), .B(n73544), .Y(n26138) );
  NAND2X1 U53557 ( .A(n29597), .B(n29598), .Y(n28520) );
  NAND2X1 U53558 ( .A(opcode_instr_w_55), .B(n73544), .Y(n28181) );
  INVX1 U53559 ( .A(n28181), .Y(n73419) );
  NAND2X1 U53560 ( .A(opcode_instr_w_57), .B(n73544), .Y(n51126) );
  NAND2X1 U53561 ( .A(n29627), .B(n51126), .Y(n28227) );
  INVX1 U53562 ( .A(n28227), .Y(n73420) );
  NAND2X1 U53563 ( .A(n72840), .B(n73420), .Y(n51127) );
  NOR2X1 U53564 ( .A(n73419), .B(n51127), .Y(n51130) );
  NOR2X1 U53565 ( .A(n28544), .B(n575), .Y(n51128) );
  NOR2X1 U53566 ( .A(n29620), .B(n51128), .Y(n51129) );
  NAND2X1 U53567 ( .A(n51130), .B(n51129), .Y(n28235) );
  NOR2X1 U53568 ( .A(n57414), .B(n58517), .Y(u_decode_N772) );
  NOR2X1 U53569 ( .A(n55035), .B(n58517), .Y(u_decode_N773) );
  AND2X1 U53570 ( .A(n29571), .B(n57360), .Y(n51132) );
  NOR2X1 U53571 ( .A(opcode_instr_w_37), .B(opcode_instr_w_36), .Y(n51131) );
  NAND2X1 U53572 ( .A(n51132), .B(n51131), .Y(n28558) );
  INVX1 U53573 ( .A(n28235), .Y(n73418) );
  INVX1 U53574 ( .A(n28558), .Y(n51133) );
  NAND2X1 U53575 ( .A(n73418), .B(n51133), .Y(n474) );
  INVX1 U53576 ( .A(n28520), .Y(n73519) );
  INVX1 U53577 ( .A(n474), .Y(n51964) );
  NAND2X1 U53578 ( .A(n73519), .B(n51964), .Y(n28035) );
  NOR2X1 U53579 ( .A(n16966), .B(n16967), .Y(n51135) );
  NOR2X1 U53580 ( .A(n17019), .B(n17020), .Y(n51134) );
  NAND2X1 U53581 ( .A(n51135), .B(n51134), .Y(u_exec_alu_p_w[13]) );
  NOR2X1 U53582 ( .A(n44539), .B(n43087), .Y(n51137) );
  NOR2X1 U53583 ( .A(n44535), .B(n37670), .Y(n51136) );
  NOR2X1 U53584 ( .A(n51137), .B(n51136), .Y(n51139) );
  NOR2X1 U53585 ( .A(n19789), .B(n19788), .Y(n51138) );
  NAND2X1 U53586 ( .A(n51139), .B(n51138), .Y(u_decode_u_regfile_N668) );
  NOR2X1 U53587 ( .A(n44601), .B(n43088), .Y(n51141) );
  NOR2X1 U53588 ( .A(n44598), .B(n37670), .Y(n51140) );
  NOR2X1 U53589 ( .A(n51141), .B(n51140), .Y(n51143) );
  NOR2X1 U53590 ( .A(n18216), .B(n18214), .Y(n51142) );
  NAND2X1 U53591 ( .A(n51143), .B(n51142), .Y(u_decode_u_regfile_N964) );
  NOR2X1 U53592 ( .A(n43086), .B(n43270), .Y(n51145) );
  NOR2X1 U53593 ( .A(n43089), .B(n43388), .Y(n51144) );
  NOR2X1 U53594 ( .A(n51145), .B(n51144), .Y(n51147) );
  NOR2X1 U53595 ( .A(n21359), .B(n21358), .Y(n51146) );
  NAND2X1 U53596 ( .A(n51147), .B(n51146), .Y(u_decode_u_regfile_N372) );
  NOR2X1 U53597 ( .A(n44472), .B(n43088), .Y(n51149) );
  NOR2X1 U53598 ( .A(n44469), .B(n37670), .Y(n51148) );
  NOR2X1 U53599 ( .A(n51149), .B(n51148), .Y(n51151) );
  NOR2X1 U53600 ( .A(n20966), .B(n20965), .Y(n51150) );
  NAND2X1 U53601 ( .A(n51151), .B(n51150), .Y(u_decode_u_regfile_N446) );
  NOR2X1 U53602 ( .A(n44559), .B(n43088), .Y(n51153) );
  NOR2X1 U53603 ( .A(n44556), .B(n37670), .Y(n51152) );
  NOR2X1 U53604 ( .A(n51153), .B(n51152), .Y(n51155) );
  NOR2X1 U53605 ( .A(n19394), .B(n19393), .Y(n51154) );
  NAND2X1 U53606 ( .A(n51155), .B(n51154), .Y(u_decode_u_regfile_N742) );
  NOR2X1 U53607 ( .A(n44382), .B(n43088), .Y(n51157) );
  NOR2X1 U53608 ( .A(n44379), .B(n43090), .Y(n51156) );
  NOR2X1 U53609 ( .A(n51157), .B(n51156), .Y(n51159) );
  NOR2X1 U53610 ( .A(n22536), .B(n22535), .Y(n51158) );
  NAND2X1 U53611 ( .A(n51159), .B(n51158), .Y(u_decode_u_regfile_N150) );
  NOR2X1 U53612 ( .A(n44304), .B(n43088), .Y(n51161) );
  NOR2X1 U53613 ( .A(n44301), .B(n43090), .Y(n51160) );
  NOR2X1 U53614 ( .A(n51161), .B(n51160), .Y(n51163) );
  NOR2X1 U53615 ( .A(n23884), .B(n23883), .Y(n51162) );
  NAND2X1 U53616 ( .A(n51163), .B(n51162), .Y(u_decode_u_regfile_N1038) );
  NOR2X1 U53617 ( .A(n44571), .B(n43088), .Y(n51165) );
  NOR2X1 U53618 ( .A(n44568), .B(n43090), .Y(n51164) );
  NOR2X1 U53619 ( .A(n51165), .B(n51164), .Y(n51167) );
  NOR2X1 U53620 ( .A(n19002), .B(n19001), .Y(n51166) );
  NAND2X1 U53621 ( .A(n51167), .B(n51166), .Y(u_decode_u_regfile_N816) );
  NOR2X1 U53622 ( .A(n43086), .B(n43276), .Y(n51169) );
  NOR2X1 U53623 ( .A(n43089), .B(n43385), .Y(n51168) );
  NOR2X1 U53624 ( .A(n51169), .B(n51168), .Y(n51171) );
  NOR2X1 U53625 ( .A(n20574), .B(n20573), .Y(n51170) );
  NAND2X1 U53626 ( .A(n51171), .B(n51170), .Y(u_decode_u_regfile_N520) );
  NOR2X1 U53627 ( .A(n44406), .B(n43087), .Y(n51173) );
  NOR2X1 U53628 ( .A(n44403), .B(n43090), .Y(n51172) );
  NOR2X1 U53629 ( .A(n51173), .B(n51172), .Y(n51175) );
  NOR2X1 U53630 ( .A(n22144), .B(n22143), .Y(n51174) );
  NAND2X1 U53631 ( .A(n51175), .B(n51174), .Y(u_decode_u_regfile_N224) );
  NOR2X1 U53632 ( .A(n44328), .B(n43087), .Y(n51177) );
  NOR2X1 U53633 ( .A(n44325), .B(n43090), .Y(n51176) );
  NOR2X1 U53634 ( .A(n51177), .B(n51176), .Y(n51179) );
  NOR2X1 U53635 ( .A(n23444), .B(n23443), .Y(n51178) );
  NAND2X1 U53636 ( .A(n51179), .B(n51178), .Y(u_decode_u_regfile_N1112) );
  NOR2X1 U53637 ( .A(n44583), .B(n43087), .Y(n51181) );
  NOR2X1 U53638 ( .A(n44580), .B(n43090), .Y(n51180) );
  NOR2X1 U53639 ( .A(n51181), .B(n51180), .Y(n51183) );
  NOR2X1 U53640 ( .A(n18610), .B(n18609), .Y(n51182) );
  NAND2X1 U53641 ( .A(n51183), .B(n51182), .Y(u_decode_u_regfile_N890) );
  NOR2X1 U53642 ( .A(n44430), .B(n43087), .Y(n51185) );
  NOR2X1 U53643 ( .A(n44427), .B(n43090), .Y(n51184) );
  NOR2X1 U53644 ( .A(n51185), .B(n51184), .Y(n51187) );
  NOR2X1 U53645 ( .A(n21752), .B(n21751), .Y(n51186) );
  NAND2X1 U53646 ( .A(n51187), .B(n51186), .Y(u_decode_u_regfile_N298) );
  NOR2X1 U53647 ( .A(n44514), .B(n43087), .Y(n51189) );
  NOR2X1 U53648 ( .A(n44511), .B(n43090), .Y(n51188) );
  NOR2X1 U53649 ( .A(n51189), .B(n51188), .Y(n51191) );
  NOR2X1 U53650 ( .A(n20182), .B(n20181), .Y(n51190) );
  NAND2X1 U53651 ( .A(n51191), .B(n51190), .Y(u_decode_u_regfile_N594) );
  NOR2X1 U53652 ( .A(n44352), .B(n43087), .Y(n51193) );
  NOR2X1 U53653 ( .A(n44349), .B(n43090), .Y(n51192) );
  NOR2X1 U53654 ( .A(n51193), .B(n51192), .Y(n51195) );
  NOR2X1 U53655 ( .A(n23010), .B(n23009), .Y(n51194) );
  NAND2X1 U53656 ( .A(n51195), .B(n51194), .Y(u_decode_u_regfile_N1186) );
  NOR2X1 U53657 ( .A(n44607), .B(n43087), .Y(n51197) );
  NOR2X1 U53658 ( .A(n44604), .B(n43090), .Y(n51196) );
  NOR2X1 U53659 ( .A(n51197), .B(n51196), .Y(n51199) );
  NOR2X1 U53660 ( .A(n24094), .B(n24093), .Y(n51198) );
  NAND2X1 U53661 ( .A(n51199), .B(n51198), .Y(u_decode_u_regfile_N1001) );
  NOR2X1 U53662 ( .A(n43086), .B(n43273), .Y(n51201) );
  NOR2X1 U53663 ( .A(n43089), .B(n43391), .Y(n51200) );
  NOR2X1 U53664 ( .A(n51201), .B(n51200), .Y(n51203) );
  NOR2X1 U53665 ( .A(n23330), .B(n23329), .Y(n51202) );
  NAND2X1 U53666 ( .A(n51203), .B(n51202), .Y(u_decode_u_regfile_N113) );
  NOR2X1 U53667 ( .A(n44460), .B(n43087), .Y(n51205) );
  NOR2X1 U53668 ( .A(n44457), .B(n43090), .Y(n51204) );
  NOR2X1 U53669 ( .A(n51205), .B(n51204), .Y(n51207) );
  NOR2X1 U53670 ( .A(n21162), .B(n21161), .Y(n51206) );
  NAND2X1 U53671 ( .A(n51207), .B(n51206), .Y(u_decode_u_regfile_N409) );
  NOR2X1 U53672 ( .A(n44550), .B(n43087), .Y(n51209) );
  NOR2X1 U53673 ( .A(n44547), .B(n43090), .Y(n51208) );
  NOR2X1 U53674 ( .A(n51209), .B(n51208), .Y(n51211) );
  NOR2X1 U53675 ( .A(n19592), .B(n19591), .Y(n51210) );
  NAND2X1 U53676 ( .A(n51211), .B(n51210), .Y(u_decode_u_regfile_N705) );
  NOR2X1 U53677 ( .A(n44565), .B(n43087), .Y(n51213) );
  NOR2X1 U53678 ( .A(n44562), .B(n43089), .Y(n51212) );
  NOR2X1 U53679 ( .A(n51213), .B(n51212), .Y(n51215) );
  NOR2X1 U53680 ( .A(n19198), .B(n19197), .Y(n51214) );
  NAND2X1 U53681 ( .A(n51215), .B(n51214), .Y(u_decode_u_regfile_N779) );
  NOR2X1 U53682 ( .A(n44316), .B(n43087), .Y(n51217) );
  NOR2X1 U53683 ( .A(n44313), .B(n43089), .Y(n51216) );
  NOR2X1 U53684 ( .A(n51217), .B(n51216), .Y(n51219) );
  NOR2X1 U53685 ( .A(n23664), .B(n23663), .Y(n51218) );
  NAND2X1 U53686 ( .A(n51219), .B(n51218), .Y(u_decode_u_regfile_N1075) );
  NOR2X1 U53687 ( .A(n44394), .B(n43087), .Y(n51221) );
  NOR2X1 U53688 ( .A(n44391), .B(n43089), .Y(n51220) );
  NOR2X1 U53689 ( .A(n51221), .B(n51220), .Y(n51223) );
  NOR2X1 U53690 ( .A(n22340), .B(n22339), .Y(n51222) );
  NAND2X1 U53691 ( .A(n51223), .B(n51222), .Y(u_decode_u_regfile_N187) );
  NOR2X1 U53692 ( .A(n44484), .B(n43086), .Y(n51225) );
  NOR2X1 U53693 ( .A(n44481), .B(n43089), .Y(n51224) );
  NOR2X1 U53694 ( .A(n51225), .B(n51224), .Y(n51227) );
  NOR2X1 U53695 ( .A(n20770), .B(n20769), .Y(n51226) );
  NAND2X1 U53696 ( .A(n51227), .B(n51226), .Y(u_decode_u_regfile_N483) );
  NOR2X1 U53697 ( .A(n44418), .B(n43086), .Y(n51229) );
  NOR2X1 U53698 ( .A(n44415), .B(n43089), .Y(n51228) );
  NOR2X1 U53699 ( .A(n51229), .B(n51228), .Y(n51231) );
  NOR2X1 U53700 ( .A(n21948), .B(n21947), .Y(n51230) );
  NAND2X1 U53701 ( .A(n51231), .B(n51230), .Y(u_decode_u_regfile_N261) );
  NOR2X1 U53702 ( .A(n44340), .B(n43086), .Y(n51233) );
  NOR2X1 U53703 ( .A(n44337), .B(n43089), .Y(n51232) );
  NOR2X1 U53704 ( .A(n51233), .B(n51232), .Y(n51235) );
  NOR2X1 U53705 ( .A(n23230), .B(n23229), .Y(n51234) );
  NAND2X1 U53706 ( .A(n51235), .B(n51234), .Y(u_decode_u_regfile_N1149) );
  NOR2X1 U53707 ( .A(n44502), .B(n43086), .Y(n51237) );
  NOR2X1 U53708 ( .A(n44499), .B(n43089), .Y(n51236) );
  NOR2X1 U53709 ( .A(n51237), .B(n51236), .Y(n51239) );
  NOR2X1 U53710 ( .A(n20378), .B(n20377), .Y(n51238) );
  NAND2X1 U53711 ( .A(n51239), .B(n51238), .Y(u_decode_u_regfile_N557) );
  NOR2X1 U53712 ( .A(n44577), .B(n43086), .Y(n51241) );
  NOR2X1 U53713 ( .A(n44574), .B(n43089), .Y(n51240) );
  NOR2X1 U53714 ( .A(n51241), .B(n51240), .Y(n51243) );
  NOR2X1 U53715 ( .A(n18806), .B(n18805), .Y(n51242) );
  NAND2X1 U53716 ( .A(n51243), .B(n51242), .Y(u_decode_u_regfile_N853) );
  NOR2X1 U53717 ( .A(n44526), .B(n43086), .Y(n51245) );
  NOR2X1 U53718 ( .A(n44523), .B(n43089), .Y(n51244) );
  NOR2X1 U53719 ( .A(n51245), .B(n51244), .Y(n51247) );
  NOR2X1 U53720 ( .A(n19986), .B(n19985), .Y(n51246) );
  NAND2X1 U53721 ( .A(n51247), .B(n51246), .Y(u_decode_u_regfile_N631) );
  NOR2X1 U53722 ( .A(n44592), .B(n43086), .Y(n51249) );
  NOR2X1 U53723 ( .A(n44589), .B(n43090), .Y(n51248) );
  NOR2X1 U53724 ( .A(n51249), .B(n51248), .Y(n51251) );
  NOR2X1 U53725 ( .A(n18416), .B(n18415), .Y(n51250) );
  NAND2X1 U53726 ( .A(n51251), .B(n51250), .Y(u_decode_u_regfile_N927) );
  NOR2X1 U53727 ( .A(n44364), .B(n43086), .Y(n51253) );
  NOR2X1 U53728 ( .A(n44361), .B(n43089), .Y(n51252) );
  NOR2X1 U53729 ( .A(n51253), .B(n51252), .Y(n51255) );
  NOR2X1 U53730 ( .A(n22790), .B(n22789), .Y(n51254) );
  NAND2X1 U53731 ( .A(n51255), .B(n51254), .Y(u_decode_u_regfile_N1223) );
  NOR2X1 U53732 ( .A(n44442), .B(n43087), .Y(n51257) );
  NOR2X1 U53733 ( .A(n44439), .B(n43090), .Y(n51256) );
  NOR2X1 U53734 ( .A(n51257), .B(n51256), .Y(n51259) );
  NOR2X1 U53735 ( .A(n21556), .B(n21555), .Y(n51258) );
  NAND2X1 U53736 ( .A(n51259), .B(n51258), .Y(u_decode_u_regfile_N335) );
  NOR2X1 U53737 ( .A(n44835), .B(n58457), .Y(n51260) );
  NAND2X1 U53738 ( .A(n51260), .B(n57889), .Y(n51979) );
  NOR2X1 U53739 ( .A(n42747), .B(n51979), .Y(n51261) );
  NAND2X1 U53740 ( .A(n51261), .B(n73364), .Y(n58816) );
  NOR2X1 U53741 ( .A(n73367), .B(n58816), .Y(n51262) );
  NAND2X1 U53742 ( .A(n51262), .B(n58818), .Y(n24942) );
  NAND2X1 U53743 ( .A(n43002), .B(n43874), .Y(n73121) );
  NAND2X1 U53744 ( .A(n28045), .B(n73121), .Y(n51263) );
  NAND2X1 U53745 ( .A(u_csr_csr_medeleg_q[13]), .B(n51263), .Y(n51265) );
  INVX1 U53746 ( .A(n24942), .Y(n58233) );
  NAND2X1 U53747 ( .A(n38609), .B(n58233), .Y(n58205) );
  INVX1 U53748 ( .A(n58205), .Y(n58229) );
  NAND2X1 U53749 ( .A(n73522), .B(n42442), .Y(n58234) );
  INVX1 U53750 ( .A(n58234), .Y(n73173) );
  NAND2X1 U53751 ( .A(n42143), .B(n43871), .Y(n51264) );
  NAND2X1 U53752 ( .A(n51265), .B(n51264), .Y(u_csr_csr_medeleg_r[13]) );
  MX2X1 U53753 ( .A(n42441), .B(u_mmu_load_q), .S0(n8574), .Y(n8441) );
  NOR2X1 U53754 ( .A(n16860), .B(n16861), .Y(n51267) );
  NOR2X1 U53755 ( .A(n16900), .B(n16901), .Y(n51266) );
  NAND2X1 U53756 ( .A(n51267), .B(n51266), .Y(u_exec_alu_p_w[15]) );
  NOR2X1 U53757 ( .A(n44539), .B(n43093), .Y(n51269) );
  NOR2X1 U53758 ( .A(n44535), .B(n37671), .Y(n51268) );
  NOR2X1 U53759 ( .A(n51269), .B(n51268), .Y(n51271) );
  NOR2X1 U53760 ( .A(n19777), .B(n19776), .Y(n51270) );
  NAND2X1 U53761 ( .A(n51271), .B(n51270), .Y(u_decode_u_regfile_N670) );
  NOR2X1 U53762 ( .A(n44601), .B(n43094), .Y(n51273) );
  NOR2X1 U53763 ( .A(n44598), .B(n37671), .Y(n51272) );
  NOR2X1 U53764 ( .A(n51273), .B(n51272), .Y(n51275) );
  NOR2X1 U53765 ( .A(n18202), .B(n18200), .Y(n51274) );
  NAND2X1 U53766 ( .A(n51275), .B(n51274), .Y(u_decode_u_regfile_N966) );
  NOR2X1 U53767 ( .A(n43092), .B(n43270), .Y(n51277) );
  NOR2X1 U53768 ( .A(n43095), .B(n43388), .Y(n51276) );
  NOR2X1 U53769 ( .A(n51277), .B(n51276), .Y(n51279) );
  NOR2X1 U53770 ( .A(n21347), .B(n21346), .Y(n51278) );
  NAND2X1 U53771 ( .A(n51279), .B(n51278), .Y(u_decode_u_regfile_N374) );
  NOR2X1 U53772 ( .A(n44472), .B(n43094), .Y(n51281) );
  NOR2X1 U53773 ( .A(n44469), .B(n37671), .Y(n51280) );
  NOR2X1 U53774 ( .A(n51281), .B(n51280), .Y(n51283) );
  NOR2X1 U53775 ( .A(n20954), .B(n20953), .Y(n51282) );
  NAND2X1 U53776 ( .A(n51283), .B(n51282), .Y(u_decode_u_regfile_N448) );
  NOR2X1 U53777 ( .A(n44559), .B(n43094), .Y(n51285) );
  NOR2X1 U53778 ( .A(n44556), .B(n37671), .Y(n51284) );
  NOR2X1 U53779 ( .A(n51285), .B(n51284), .Y(n51287) );
  NOR2X1 U53780 ( .A(n19382), .B(n19381), .Y(n51286) );
  NAND2X1 U53781 ( .A(n51287), .B(n51286), .Y(u_decode_u_regfile_N744) );
  NOR2X1 U53782 ( .A(n44382), .B(n43094), .Y(n51289) );
  NOR2X1 U53783 ( .A(n44379), .B(n43096), .Y(n51288) );
  NOR2X1 U53784 ( .A(n51289), .B(n51288), .Y(n51291) );
  NOR2X1 U53785 ( .A(n22524), .B(n22523), .Y(n51290) );
  NAND2X1 U53786 ( .A(n51291), .B(n51290), .Y(u_decode_u_regfile_N152) );
  NOR2X1 U53787 ( .A(n44304), .B(n43094), .Y(n51293) );
  NOR2X1 U53788 ( .A(n44301), .B(n43096), .Y(n51292) );
  NOR2X1 U53789 ( .A(n51293), .B(n51292), .Y(n51295) );
  NOR2X1 U53790 ( .A(n23866), .B(n23865), .Y(n51294) );
  NAND2X1 U53791 ( .A(n51295), .B(n51294), .Y(u_decode_u_regfile_N1040) );
  NOR2X1 U53792 ( .A(n44571), .B(n43094), .Y(n51297) );
  NOR2X1 U53793 ( .A(n44568), .B(n43096), .Y(n51296) );
  NOR2X1 U53794 ( .A(n51297), .B(n51296), .Y(n51299) );
  NOR2X1 U53795 ( .A(n18990), .B(n18989), .Y(n51298) );
  NAND2X1 U53796 ( .A(n51299), .B(n51298), .Y(u_decode_u_regfile_N818) );
  NOR2X1 U53797 ( .A(n43092), .B(n43276), .Y(n51301) );
  NOR2X1 U53798 ( .A(n43095), .B(n43385), .Y(n51300) );
  NOR2X1 U53799 ( .A(n51301), .B(n51300), .Y(n51303) );
  NOR2X1 U53800 ( .A(n20562), .B(n20561), .Y(n51302) );
  NAND2X1 U53801 ( .A(n51303), .B(n51302), .Y(u_decode_u_regfile_N522) );
  NOR2X1 U53802 ( .A(n44406), .B(n43093), .Y(n51305) );
  NOR2X1 U53803 ( .A(n44403), .B(n43096), .Y(n51304) );
  NOR2X1 U53804 ( .A(n51305), .B(n51304), .Y(n51307) );
  NOR2X1 U53805 ( .A(n22132), .B(n22131), .Y(n51306) );
  NAND2X1 U53806 ( .A(n51307), .B(n51306), .Y(u_decode_u_regfile_N226) );
  NOR2X1 U53807 ( .A(n44328), .B(n43093), .Y(n51309) );
  NOR2X1 U53808 ( .A(n44325), .B(n43096), .Y(n51308) );
  NOR2X1 U53809 ( .A(n51309), .B(n51308), .Y(n51311) );
  NOR2X1 U53810 ( .A(n23432), .B(n23431), .Y(n51310) );
  NAND2X1 U53811 ( .A(n51311), .B(n51310), .Y(u_decode_u_regfile_N1114) );
  NOR2X1 U53812 ( .A(n44583), .B(n43093), .Y(n51313) );
  NOR2X1 U53813 ( .A(n44580), .B(n43096), .Y(n51312) );
  NOR2X1 U53814 ( .A(n51313), .B(n51312), .Y(n51315) );
  NOR2X1 U53815 ( .A(n18598), .B(n18597), .Y(n51314) );
  NAND2X1 U53816 ( .A(n51315), .B(n51314), .Y(u_decode_u_regfile_N892) );
  NOR2X1 U53817 ( .A(n44430), .B(n43093), .Y(n51317) );
  NOR2X1 U53818 ( .A(n44427), .B(n43096), .Y(n51316) );
  NOR2X1 U53819 ( .A(n51317), .B(n51316), .Y(n51319) );
  NOR2X1 U53820 ( .A(n21740), .B(n21739), .Y(n51318) );
  NAND2X1 U53821 ( .A(n51319), .B(n51318), .Y(u_decode_u_regfile_N300) );
  NOR2X1 U53822 ( .A(n44514), .B(n43093), .Y(n51321) );
  NOR2X1 U53823 ( .A(n44511), .B(n43096), .Y(n51320) );
  NOR2X1 U53824 ( .A(n51321), .B(n51320), .Y(n51323) );
  NOR2X1 U53825 ( .A(n20170), .B(n20169), .Y(n51322) );
  NAND2X1 U53826 ( .A(n51323), .B(n51322), .Y(u_decode_u_regfile_N596) );
  NOR2X1 U53827 ( .A(n44352), .B(n43093), .Y(n51325) );
  NOR2X1 U53828 ( .A(n44349), .B(n43096), .Y(n51324) );
  NOR2X1 U53829 ( .A(n51325), .B(n51324), .Y(n51327) );
  NOR2X1 U53830 ( .A(n22998), .B(n22997), .Y(n51326) );
  NAND2X1 U53831 ( .A(n51327), .B(n51326), .Y(u_decode_u_regfile_N1188) );
  NOR2X1 U53832 ( .A(n44607), .B(n43093), .Y(n51329) );
  NOR2X1 U53833 ( .A(n44604), .B(n43096), .Y(n51328) );
  NOR2X1 U53834 ( .A(n51329), .B(n51328), .Y(n51331) );
  NOR2X1 U53835 ( .A(n24082), .B(n24081), .Y(n51330) );
  NAND2X1 U53836 ( .A(n51331), .B(n51330), .Y(u_decode_u_regfile_N1003) );
  NOR2X1 U53837 ( .A(n43092), .B(n43273), .Y(n51333) );
  NOR2X1 U53838 ( .A(n43095), .B(n43391), .Y(n51332) );
  NOR2X1 U53839 ( .A(n51333), .B(n51332), .Y(n51335) );
  NOR2X1 U53840 ( .A(n23224), .B(n23223), .Y(n51334) );
  NAND2X1 U53841 ( .A(n51335), .B(n51334), .Y(u_decode_u_regfile_N115) );
  NOR2X1 U53842 ( .A(n44460), .B(n43093), .Y(n51337) );
  NOR2X1 U53843 ( .A(n44457), .B(n43096), .Y(n51336) );
  NOR2X1 U53844 ( .A(n51337), .B(n51336), .Y(n51339) );
  NOR2X1 U53845 ( .A(n21150), .B(n21149), .Y(n51338) );
  NAND2X1 U53846 ( .A(n51339), .B(n51338), .Y(u_decode_u_regfile_N411) );
  NOR2X1 U53847 ( .A(n44550), .B(n43093), .Y(n51341) );
  NOR2X1 U53848 ( .A(n44547), .B(n43096), .Y(n51340) );
  NOR2X1 U53849 ( .A(n51341), .B(n51340), .Y(n51343) );
  NOR2X1 U53850 ( .A(n19580), .B(n19579), .Y(n51342) );
  NAND2X1 U53851 ( .A(n51343), .B(n51342), .Y(u_decode_u_regfile_N707) );
  NOR2X1 U53852 ( .A(n44565), .B(n43093), .Y(n51345) );
  NOR2X1 U53853 ( .A(n44562), .B(n43095), .Y(n51344) );
  NOR2X1 U53854 ( .A(n51345), .B(n51344), .Y(n51347) );
  NOR2X1 U53855 ( .A(n19186), .B(n19185), .Y(n51346) );
  NAND2X1 U53856 ( .A(n51347), .B(n51346), .Y(u_decode_u_regfile_N781) );
  NOR2X1 U53857 ( .A(n44316), .B(n43093), .Y(n51349) );
  NOR2X1 U53858 ( .A(n44313), .B(n43095), .Y(n51348) );
  NOR2X1 U53859 ( .A(n51349), .B(n51348), .Y(n51351) );
  NOR2X1 U53860 ( .A(n23652), .B(n23651), .Y(n51350) );
  NAND2X1 U53861 ( .A(n51351), .B(n51350), .Y(u_decode_u_regfile_N1077) );
  NOR2X1 U53862 ( .A(n44394), .B(n43093), .Y(n51353) );
  NOR2X1 U53863 ( .A(n44391), .B(n43095), .Y(n51352) );
  NOR2X1 U53864 ( .A(n51353), .B(n51352), .Y(n51355) );
  NOR2X1 U53865 ( .A(n22328), .B(n22327), .Y(n51354) );
  NAND2X1 U53866 ( .A(n51355), .B(n51354), .Y(u_decode_u_regfile_N189) );
  NOR2X1 U53867 ( .A(n44484), .B(n43092), .Y(n51357) );
  NOR2X1 U53868 ( .A(n44481), .B(n43095), .Y(n51356) );
  NOR2X1 U53869 ( .A(n51357), .B(n51356), .Y(n51359) );
  NOR2X1 U53870 ( .A(n20758), .B(n20757), .Y(n51358) );
  NAND2X1 U53871 ( .A(n51359), .B(n51358), .Y(u_decode_u_regfile_N485) );
  NOR2X1 U53872 ( .A(n44418), .B(n43092), .Y(n51361) );
  NOR2X1 U53873 ( .A(n44415), .B(n43095), .Y(n51360) );
  NOR2X1 U53874 ( .A(n51361), .B(n51360), .Y(n51363) );
  NOR2X1 U53875 ( .A(n21936), .B(n21935), .Y(n51362) );
  NAND2X1 U53876 ( .A(n51363), .B(n51362), .Y(u_decode_u_regfile_N263) );
  NOR2X1 U53877 ( .A(n44340), .B(n43092), .Y(n51365) );
  NOR2X1 U53878 ( .A(n44337), .B(n43095), .Y(n51364) );
  NOR2X1 U53879 ( .A(n51365), .B(n51364), .Y(n51367) );
  NOR2X1 U53880 ( .A(n23212), .B(n23211), .Y(n51366) );
  NAND2X1 U53881 ( .A(n51367), .B(n51366), .Y(u_decode_u_regfile_N1151) );
  NOR2X1 U53882 ( .A(n44502), .B(n43092), .Y(n51369) );
  NOR2X1 U53883 ( .A(n44499), .B(n43095), .Y(n51368) );
  NOR2X1 U53884 ( .A(n51369), .B(n51368), .Y(n51371) );
  NOR2X1 U53885 ( .A(n20366), .B(n20365), .Y(n51370) );
  NAND2X1 U53886 ( .A(n51371), .B(n51370), .Y(u_decode_u_regfile_N559) );
  NOR2X1 U53887 ( .A(n44577), .B(n43092), .Y(n51373) );
  NOR2X1 U53888 ( .A(n44574), .B(n43095), .Y(n51372) );
  NOR2X1 U53889 ( .A(n51373), .B(n51372), .Y(n51375) );
  NOR2X1 U53890 ( .A(n18794), .B(n18793), .Y(n51374) );
  NAND2X1 U53891 ( .A(n51375), .B(n51374), .Y(u_decode_u_regfile_N855) );
  NOR2X1 U53892 ( .A(n44526), .B(n43092), .Y(n51377) );
  NOR2X1 U53893 ( .A(n44523), .B(n43095), .Y(n51376) );
  NOR2X1 U53894 ( .A(n51377), .B(n51376), .Y(n51379) );
  NOR2X1 U53895 ( .A(n19974), .B(n19973), .Y(n51378) );
  NAND2X1 U53896 ( .A(n51379), .B(n51378), .Y(u_decode_u_regfile_N633) );
  NOR2X1 U53897 ( .A(n44592), .B(n43092), .Y(n51381) );
  NOR2X1 U53898 ( .A(n44589), .B(n43096), .Y(n51380) );
  NOR2X1 U53899 ( .A(n51381), .B(n51380), .Y(n51383) );
  NOR2X1 U53900 ( .A(n18404), .B(n18403), .Y(n51382) );
  NAND2X1 U53901 ( .A(n51383), .B(n51382), .Y(u_decode_u_regfile_N929) );
  NOR2X1 U53902 ( .A(n44364), .B(n43092), .Y(n51385) );
  NOR2X1 U53903 ( .A(n44361), .B(n43095), .Y(n51384) );
  NOR2X1 U53904 ( .A(n51385), .B(n51384), .Y(n51387) );
  NOR2X1 U53905 ( .A(n22778), .B(n22777), .Y(n51386) );
  NAND2X1 U53906 ( .A(n51387), .B(n51386), .Y(u_decode_u_regfile_N1225) );
  NOR2X1 U53907 ( .A(n44442), .B(n43093), .Y(n51389) );
  NOR2X1 U53908 ( .A(n44439), .B(n43096), .Y(n51388) );
  NOR2X1 U53909 ( .A(n51389), .B(n51388), .Y(n51391) );
  NOR2X1 U53910 ( .A(n21544), .B(n21543), .Y(n51390) );
  NAND2X1 U53911 ( .A(n51391), .B(n51390), .Y(u_decode_u_regfile_N337) );
  NAND2X1 U53912 ( .A(n43003), .B(n43895), .Y(n73114) );
  NAND2X1 U53913 ( .A(n28045), .B(n73114), .Y(n51392) );
  NAND2X1 U53914 ( .A(u_csr_csr_medeleg_q[15]), .B(n51392), .Y(n51394) );
  NAND2X1 U53915 ( .A(n42143), .B(n43892), .Y(n51393) );
  NAND2X1 U53916 ( .A(n51394), .B(n51393), .Y(u_csr_csr_medeleg_r[15]) );
  INVX1 U53917 ( .A(n58218), .Y(n72839) );
  NAND2X1 U53918 ( .A(u_csr_csr_medeleg_q[13]), .B(n72839), .Y(n51395) );
  AND2X1 U53919 ( .A(n28549), .B(n51395), .Y(n51397) );
  INVX1 U53920 ( .A(n58216), .Y(n58191) );
  NAND2X1 U53921 ( .A(u_csr_csr_medeleg_q[15]), .B(n58191), .Y(n51396) );
  NAND2X1 U53922 ( .A(n51397), .B(n51396), .Y(n28536) );
  NOR2X1 U53923 ( .A(n28536), .B(n72840), .Y(n51398) );
  NAND2X1 U53924 ( .A(n26931), .B(n28235), .Y(n28179) );
  NAND2X1 U53925 ( .A(n28035), .B(n28179), .Y(n26976) );
  NAND2X1 U53926 ( .A(n24508), .B(n73533), .Y(n51399) );
  OR2X1 U53927 ( .A(n24511), .B(n51399), .Y(n24440) );
  NOR2X1 U53928 ( .A(n24440), .B(n58514), .Y(n51400) );
  NAND2X1 U53929 ( .A(n51400), .B(n57581), .Y(n51405) );
  INVX1 U53930 ( .A(n51405), .Y(n51404) );
  INVX1 U53931 ( .A(n51401), .Y(n51402) );
  OR2X1 U53932 ( .A(n24502), .B(n51402), .Y(n51403) );
  NAND2X1 U53933 ( .A(n51404), .B(n51403), .Y(n57585) );
  NOR2X1 U53934 ( .A(n42932), .B(n57585), .Y(u_decode_N775) );
  NOR2X1 U53935 ( .A(n24437), .B(n51405), .Y(n51406) );
  NAND2X1 U53936 ( .A(n51406), .B(n24435), .Y(n58515) );
  NOR2X1 U53937 ( .A(n42932), .B(n58515), .Y(u_decode_N774) );
  NAND2X1 U53938 ( .A(n58249), .B(n51407), .Y(n971) );
  NAND2X1 U53939 ( .A(n971), .B(n73544), .Y(n28031) );
  NOR2X1 U53940 ( .A(n24535), .B(n57401), .Y(n51410) );
  NOR2X1 U53941 ( .A(n24533), .B(n51408), .Y(n51409) );
  NAND2X1 U53942 ( .A(n51410), .B(n51409), .Y(n57563) );
  NOR2X1 U53943 ( .A(n57563), .B(n57415), .Y(u_decode_N759) );
  NOR2X1 U53944 ( .A(n57563), .B(n57406), .Y(u_decode_N764) );
  NOR2X1 U53945 ( .A(n57563), .B(n57407), .Y(u_decode_N762) );
  NOR2X1 U53946 ( .A(n57563), .B(n57404), .Y(u_decode_N763) );
  NAND2X1 U53947 ( .A(n42315), .B(n73571), .Y(n15453) );
  INVX1 U53948 ( .A(n16593), .Y(n73523) );
  NAND2X1 U53949 ( .A(n43269), .B(n44070), .Y(n51413) );
  NAND2X1 U53950 ( .A(u_csr_N184), .B(n40679), .Y(n51412) );
  NAND2X1 U53951 ( .A(n51413), .B(n51412), .Y(n58597) );
  NAND2X1 U53952 ( .A(n43424), .B(n58597), .Y(n58734) );
  INVX1 U53953 ( .A(n58734), .Y(n56797) );
  INVX1 U53954 ( .A(n15453), .Y(n73512) );
  NAND2X1 U53955 ( .A(n56797), .B(n73512), .Y(n51414) );
  NAND2X1 U53956 ( .A(n15458), .B(n51414), .Y(n51415) );
  NOR2X1 U53957 ( .A(n15487), .B(n51415), .Y(n51417) );
  NOR2X1 U53958 ( .A(n15456), .B(n15488), .Y(n51416) );
  NAND2X1 U53959 ( .A(n51417), .B(n51416), .Y(u_exec_alu_p_w[8]) );
  NOR2X1 U53960 ( .A(n44539), .B(n43099), .Y(n51419) );
  NOR2X1 U53961 ( .A(n44535), .B(n37672), .Y(n51418) );
  NOR2X1 U53962 ( .A(n51419), .B(n51418), .Y(n51421) );
  NOR2X1 U53963 ( .A(n19819), .B(n19818), .Y(n51420) );
  NAND2X1 U53964 ( .A(n51421), .B(n51420), .Y(u_decode_u_regfile_N663) );
  NOR2X1 U53965 ( .A(n44601), .B(n43100), .Y(n51423) );
  NOR2X1 U53966 ( .A(n44598), .B(n37672), .Y(n51422) );
  NOR2X1 U53967 ( .A(n51423), .B(n51422), .Y(n51425) );
  NOR2X1 U53968 ( .A(n18247), .B(n18246), .Y(n51424) );
  NAND2X1 U53969 ( .A(n51425), .B(n51424), .Y(u_decode_u_regfile_N959) );
  NOR2X1 U53970 ( .A(n43098), .B(n43270), .Y(n51427) );
  NOR2X1 U53971 ( .A(n43101), .B(n43388), .Y(n51426) );
  NOR2X1 U53972 ( .A(n51427), .B(n51426), .Y(n51429) );
  NOR2X1 U53973 ( .A(n21389), .B(n21388), .Y(n51428) );
  NAND2X1 U53974 ( .A(n51429), .B(n51428), .Y(u_decode_u_regfile_N367) );
  NOR2X1 U53975 ( .A(n44472), .B(n43100), .Y(n51431) );
  NOR2X1 U53976 ( .A(n44469), .B(n37672), .Y(n51430) );
  NOR2X1 U53977 ( .A(n51431), .B(n51430), .Y(n51433) );
  NOR2X1 U53978 ( .A(n20996), .B(n20995), .Y(n51432) );
  NAND2X1 U53979 ( .A(n51433), .B(n51432), .Y(u_decode_u_regfile_N441) );
  NOR2X1 U53980 ( .A(n44559), .B(n43100), .Y(n51435) );
  NOR2X1 U53981 ( .A(n44556), .B(n37672), .Y(n51434) );
  NOR2X1 U53982 ( .A(n51435), .B(n51434), .Y(n51437) );
  NOR2X1 U53983 ( .A(n19424), .B(n19423), .Y(n51436) );
  NAND2X1 U53984 ( .A(n51437), .B(n51436), .Y(u_decode_u_regfile_N737) );
  NOR2X1 U53985 ( .A(n44382), .B(n43100), .Y(n51439) );
  NOR2X1 U53986 ( .A(n44379), .B(n43102), .Y(n51438) );
  NOR2X1 U53987 ( .A(n51439), .B(n51438), .Y(n51441) );
  NOR2X1 U53988 ( .A(n22566), .B(n22565), .Y(n51440) );
  NAND2X1 U53989 ( .A(n51441), .B(n51440), .Y(u_decode_u_regfile_N145) );
  NOR2X1 U53990 ( .A(n44304), .B(n43100), .Y(n51443) );
  NOR2X1 U53991 ( .A(n44301), .B(n43102), .Y(n51442) );
  NOR2X1 U53992 ( .A(n51443), .B(n51442), .Y(n51445) );
  NOR2X1 U53993 ( .A(n23914), .B(n23913), .Y(n51444) );
  NAND2X1 U53994 ( .A(n51445), .B(n51444), .Y(u_decode_u_regfile_N1033) );
  NOR2X1 U53995 ( .A(n44571), .B(n43100), .Y(n51447) );
  NOR2X1 U53996 ( .A(n44568), .B(n43102), .Y(n51446) );
  NOR2X1 U53997 ( .A(n51447), .B(n51446), .Y(n51449) );
  NOR2X1 U53998 ( .A(n19032), .B(n19031), .Y(n51448) );
  NAND2X1 U53999 ( .A(n51449), .B(n51448), .Y(u_decode_u_regfile_N811) );
  NOR2X1 U54000 ( .A(n43098), .B(n43276), .Y(n51451) );
  NOR2X1 U54001 ( .A(n43101), .B(n43385), .Y(n51450) );
  NOR2X1 U54002 ( .A(n51451), .B(n51450), .Y(n51453) );
  NOR2X1 U54003 ( .A(n20604), .B(n20603), .Y(n51452) );
  NAND2X1 U54004 ( .A(n51453), .B(n51452), .Y(u_decode_u_regfile_N515) );
  NOR2X1 U54005 ( .A(n44406), .B(n43099), .Y(n51455) );
  NOR2X1 U54006 ( .A(n44403), .B(n43102), .Y(n51454) );
  NOR2X1 U54007 ( .A(n51455), .B(n51454), .Y(n51457) );
  NOR2X1 U54008 ( .A(n22174), .B(n22173), .Y(n51456) );
  NAND2X1 U54009 ( .A(n51457), .B(n51456), .Y(u_decode_u_regfile_N219) );
  NOR2X1 U54010 ( .A(n44328), .B(n43099), .Y(n51459) );
  NOR2X1 U54011 ( .A(n44325), .B(n43102), .Y(n51458) );
  NOR2X1 U54012 ( .A(n51459), .B(n51458), .Y(n51461) );
  NOR2X1 U54013 ( .A(n23480), .B(n23479), .Y(n51460) );
  NAND2X1 U54014 ( .A(n51461), .B(n51460), .Y(u_decode_u_regfile_N1107) );
  NOR2X1 U54015 ( .A(n44583), .B(n43099), .Y(n51463) );
  NOR2X1 U54016 ( .A(n44580), .B(n43102), .Y(n51462) );
  NOR2X1 U54017 ( .A(n51463), .B(n51462), .Y(n51465) );
  NOR2X1 U54018 ( .A(n18640), .B(n18639), .Y(n51464) );
  NAND2X1 U54019 ( .A(n51465), .B(n51464), .Y(u_decode_u_regfile_N885) );
  NOR2X1 U54020 ( .A(n44430), .B(n43099), .Y(n51467) );
  NOR2X1 U54021 ( .A(n44427), .B(n43102), .Y(n51466) );
  NOR2X1 U54022 ( .A(n51467), .B(n51466), .Y(n51469) );
  NOR2X1 U54023 ( .A(n21782), .B(n21781), .Y(n51468) );
  NAND2X1 U54024 ( .A(n51469), .B(n51468), .Y(u_decode_u_regfile_N293) );
  NOR2X1 U54025 ( .A(n44514), .B(n43099), .Y(n51471) );
  NOR2X1 U54026 ( .A(n44511), .B(n43102), .Y(n51470) );
  NOR2X1 U54027 ( .A(n51471), .B(n51470), .Y(n51473) );
  NOR2X1 U54028 ( .A(n20212), .B(n20211), .Y(n51472) );
  NAND2X1 U54029 ( .A(n51473), .B(n51472), .Y(u_decode_u_regfile_N589) );
  NOR2X1 U54030 ( .A(n44352), .B(n43099), .Y(n51475) );
  NOR2X1 U54031 ( .A(n44349), .B(n43102), .Y(n51474) );
  NOR2X1 U54032 ( .A(n51475), .B(n51474), .Y(n51477) );
  NOR2X1 U54033 ( .A(n23040), .B(n23039), .Y(n51476) );
  NAND2X1 U54034 ( .A(n51477), .B(n51476), .Y(u_decode_u_regfile_N1181) );
  NOR2X1 U54035 ( .A(n44607), .B(n43099), .Y(n51479) );
  NOR2X1 U54036 ( .A(n44604), .B(n43102), .Y(n51478) );
  NOR2X1 U54037 ( .A(n51479), .B(n51478), .Y(n51481) );
  NOR2X1 U54038 ( .A(n18025), .B(n18023), .Y(n51480) );
  NAND2X1 U54039 ( .A(n51481), .B(n51480), .Y(u_decode_u_regfile_N996) );
  NOR2X1 U54040 ( .A(n43098), .B(n43273), .Y(n51483) );
  NOR2X1 U54041 ( .A(n43101), .B(n43391), .Y(n51482) );
  NOR2X1 U54042 ( .A(n51483), .B(n51482), .Y(n51485) );
  NOR2X1 U54043 ( .A(n23634), .B(n23633), .Y(n51484) );
  NAND2X1 U54044 ( .A(n51485), .B(n51484), .Y(u_decode_u_regfile_N108) );
  NOR2X1 U54045 ( .A(n44460), .B(n43099), .Y(n51487) );
  NOR2X1 U54046 ( .A(n44457), .B(n43102), .Y(n51486) );
  NOR2X1 U54047 ( .A(n51487), .B(n51486), .Y(n51489) );
  NOR2X1 U54048 ( .A(n21192), .B(n21191), .Y(n51488) );
  NAND2X1 U54049 ( .A(n51489), .B(n51488), .Y(u_decode_u_regfile_N404) );
  NOR2X1 U54050 ( .A(n44550), .B(n43099), .Y(n51491) );
  NOR2X1 U54051 ( .A(n44547), .B(n43102), .Y(n51490) );
  NOR2X1 U54052 ( .A(n51491), .B(n51490), .Y(n51493) );
  NOR2X1 U54053 ( .A(n19622), .B(n19621), .Y(n51492) );
  NAND2X1 U54054 ( .A(n51493), .B(n51492), .Y(u_decode_u_regfile_N700) );
  NOR2X1 U54055 ( .A(n44565), .B(n43099), .Y(n51495) );
  NOR2X1 U54056 ( .A(n44562), .B(n43101), .Y(n51494) );
  NOR2X1 U54057 ( .A(n51495), .B(n51494), .Y(n51497) );
  NOR2X1 U54058 ( .A(n19228), .B(n19227), .Y(n51496) );
  NAND2X1 U54059 ( .A(n51497), .B(n51496), .Y(u_decode_u_regfile_N774) );
  NOR2X1 U54060 ( .A(n44316), .B(n43099), .Y(n51499) );
  NOR2X1 U54061 ( .A(n44313), .B(n43101), .Y(n51498) );
  NOR2X1 U54062 ( .A(n51499), .B(n51498), .Y(n51501) );
  NOR2X1 U54063 ( .A(n23694), .B(n23693), .Y(n51500) );
  NAND2X1 U54064 ( .A(n51501), .B(n51500), .Y(u_decode_u_regfile_N1070) );
  NOR2X1 U54065 ( .A(n44394), .B(n43099), .Y(n51503) );
  NOR2X1 U54066 ( .A(n44391), .B(n43101), .Y(n51502) );
  NOR2X1 U54067 ( .A(n51503), .B(n51502), .Y(n51505) );
  NOR2X1 U54068 ( .A(n22370), .B(n22369), .Y(n51504) );
  NAND2X1 U54069 ( .A(n51505), .B(n51504), .Y(u_decode_u_regfile_N182) );
  NOR2X1 U54070 ( .A(n44484), .B(n43098), .Y(n51507) );
  NOR2X1 U54071 ( .A(n44481), .B(n43101), .Y(n51506) );
  NOR2X1 U54072 ( .A(n51507), .B(n51506), .Y(n51509) );
  NOR2X1 U54073 ( .A(n20800), .B(n20799), .Y(n51508) );
  NAND2X1 U54074 ( .A(n51509), .B(n51508), .Y(u_decode_u_regfile_N478) );
  NOR2X1 U54075 ( .A(n44418), .B(n43098), .Y(n51511) );
  NOR2X1 U54076 ( .A(n44415), .B(n43101), .Y(n51510) );
  NOR2X1 U54077 ( .A(n51511), .B(n51510), .Y(n51513) );
  NOR2X1 U54078 ( .A(n21978), .B(n21977), .Y(n51512) );
  NAND2X1 U54079 ( .A(n51513), .B(n51512), .Y(u_decode_u_regfile_N256) );
  NOR2X1 U54080 ( .A(n44340), .B(n43098), .Y(n51515) );
  NOR2X1 U54081 ( .A(n44337), .B(n43101), .Y(n51514) );
  NOR2X1 U54082 ( .A(n51515), .B(n51514), .Y(n51517) );
  NOR2X1 U54083 ( .A(n23260), .B(n23259), .Y(n51516) );
  NAND2X1 U54084 ( .A(n51517), .B(n51516), .Y(u_decode_u_regfile_N1144) );
  NOR2X1 U54085 ( .A(n44502), .B(n43098), .Y(n51519) );
  NOR2X1 U54086 ( .A(n44499), .B(n43101), .Y(n51518) );
  NOR2X1 U54087 ( .A(n51519), .B(n51518), .Y(n51521) );
  NOR2X1 U54088 ( .A(n20408), .B(n20407), .Y(n51520) );
  NAND2X1 U54089 ( .A(n51521), .B(n51520), .Y(u_decode_u_regfile_N552) );
  NOR2X1 U54090 ( .A(n44577), .B(n43098), .Y(n51523) );
  NOR2X1 U54091 ( .A(n44574), .B(n43101), .Y(n51522) );
  NOR2X1 U54092 ( .A(n51523), .B(n51522), .Y(n51525) );
  NOR2X1 U54093 ( .A(n18836), .B(n18835), .Y(n51524) );
  NAND2X1 U54094 ( .A(n51525), .B(n51524), .Y(u_decode_u_regfile_N848) );
  NOR2X1 U54095 ( .A(n44526), .B(n43098), .Y(n51527) );
  NOR2X1 U54096 ( .A(n44523), .B(n43101), .Y(n51526) );
  NOR2X1 U54097 ( .A(n51527), .B(n51526), .Y(n51529) );
  NOR2X1 U54098 ( .A(n20016), .B(n20015), .Y(n51528) );
  NAND2X1 U54099 ( .A(n51529), .B(n51528), .Y(u_decode_u_regfile_N626) );
  NOR2X1 U54100 ( .A(n44592), .B(n43098), .Y(n51531) );
  NOR2X1 U54101 ( .A(n44589), .B(n43102), .Y(n51530) );
  NOR2X1 U54102 ( .A(n51531), .B(n51530), .Y(n51533) );
  NOR2X1 U54103 ( .A(n18446), .B(n18445), .Y(n51532) );
  NAND2X1 U54104 ( .A(n51533), .B(n51532), .Y(u_decode_u_regfile_N922) );
  NOR2X1 U54105 ( .A(n44364), .B(n43098), .Y(n51535) );
  NOR2X1 U54106 ( .A(n44361), .B(n43101), .Y(n51534) );
  NOR2X1 U54107 ( .A(n51535), .B(n51534), .Y(n51537) );
  NOR2X1 U54108 ( .A(n22826), .B(n22825), .Y(n51536) );
  NAND2X1 U54109 ( .A(n51537), .B(n51536), .Y(u_decode_u_regfile_N1218) );
  NOR2X1 U54110 ( .A(n44442), .B(n43099), .Y(n51539) );
  NOR2X1 U54111 ( .A(n44439), .B(n43102), .Y(n51538) );
  NOR2X1 U54112 ( .A(n51539), .B(n51538), .Y(n51541) );
  NOR2X1 U54113 ( .A(n21586), .B(n21585), .Y(n51540) );
  NAND2X1 U54114 ( .A(n51541), .B(n51540), .Y(u_decode_u_regfile_N330) );
  NOR2X1 U54115 ( .A(n15508), .B(n15509), .Y(n51543) );
  NOR2X1 U54116 ( .A(n15544), .B(n15545), .Y(n51542) );
  NAND2X1 U54117 ( .A(n51543), .B(n51542), .Y(u_exec_alu_p_w[7]) );
  NOR2X1 U54118 ( .A(n44364), .B(n43103), .Y(n51545) );
  NOR2X1 U54119 ( .A(n44361), .B(n37673), .Y(n51544) );
  NOR2X1 U54120 ( .A(n51545), .B(n51544), .Y(n51547) );
  NOR2X1 U54121 ( .A(n22832), .B(n22831), .Y(n51546) );
  NAND2X1 U54122 ( .A(n51547), .B(n51546), .Y(u_decode_u_regfile_N1217) );
  NOR2X1 U54123 ( .A(n44442), .B(n43105), .Y(n51549) );
  NOR2X1 U54124 ( .A(n44439), .B(n37673), .Y(n51548) );
  NOR2X1 U54125 ( .A(n51549), .B(n51548), .Y(n51551) );
  NOR2X1 U54126 ( .A(n21592), .B(n21591), .Y(n51550) );
  NAND2X1 U54127 ( .A(n51551), .B(n51550), .Y(u_decode_u_regfile_N329) );
  NOR2X1 U54128 ( .A(n44382), .B(n43105), .Y(n51553) );
  NOR2X1 U54129 ( .A(n44379), .B(n37673), .Y(n51552) );
  NOR2X1 U54130 ( .A(n51553), .B(n51552), .Y(n51555) );
  NOR2X1 U54131 ( .A(n22572), .B(n22571), .Y(n51554) );
  NAND2X1 U54132 ( .A(n51555), .B(n51554), .Y(u_decode_u_regfile_N144) );
  NOR2X1 U54133 ( .A(n44304), .B(n43105), .Y(n51557) );
  NOR2X1 U54134 ( .A(n44301), .B(n37673), .Y(n51556) );
  NOR2X1 U54135 ( .A(n51557), .B(n51556), .Y(n51559) );
  NOR2X1 U54136 ( .A(n23920), .B(n23919), .Y(n51558) );
  NAND2X1 U54137 ( .A(n51559), .B(n51558), .Y(u_decode_u_regfile_N1032) );
  NOR2X1 U54138 ( .A(n44406), .B(n43105), .Y(n51561) );
  NOR2X1 U54139 ( .A(n44403), .B(n43107), .Y(n51560) );
  NOR2X1 U54140 ( .A(n51561), .B(n51560), .Y(n51563) );
  NOR2X1 U54141 ( .A(n22180), .B(n22179), .Y(n51562) );
  NAND2X1 U54142 ( .A(n51563), .B(n51562), .Y(u_decode_u_regfile_N218) );
  NOR2X1 U54143 ( .A(n44559), .B(n43105), .Y(n51565) );
  NOR2X1 U54144 ( .A(n44556), .B(n43107), .Y(n51564) );
  NOR2X1 U54145 ( .A(n51565), .B(n51564), .Y(n51567) );
  NOR2X1 U54146 ( .A(n19430), .B(n19429), .Y(n51566) );
  NAND2X1 U54147 ( .A(n51567), .B(n51566), .Y(u_decode_u_regfile_N736) );
  NOR2X1 U54148 ( .A(n44328), .B(n43105), .Y(n51569) );
  NOR2X1 U54149 ( .A(n44325), .B(n43107), .Y(n51568) );
  NOR2X1 U54150 ( .A(n51569), .B(n51568), .Y(n51571) );
  NOR2X1 U54151 ( .A(n23486), .B(n23485), .Y(n51570) );
  NAND2X1 U54152 ( .A(n51571), .B(n51570), .Y(u_decode_u_regfile_N1106) );
  NOR2X1 U54153 ( .A(n44430), .B(n43104), .Y(n51573) );
  NOR2X1 U54154 ( .A(n44427), .B(n43107), .Y(n51572) );
  NOR2X1 U54155 ( .A(n51573), .B(n51572), .Y(n51575) );
  NOR2X1 U54156 ( .A(n21788), .B(n21787), .Y(n51574) );
  NAND2X1 U54157 ( .A(n51575), .B(n51574), .Y(u_decode_u_regfile_N292) );
  NOR2X1 U54158 ( .A(n44418), .B(n43104), .Y(n51577) );
  NOR2X1 U54159 ( .A(n44415), .B(n43107), .Y(n51576) );
  NOR2X1 U54160 ( .A(n51577), .B(n51576), .Y(n51579) );
  NOR2X1 U54161 ( .A(n21984), .B(n21983), .Y(n51578) );
  NAND2X1 U54162 ( .A(n51579), .B(n51578), .Y(u_decode_u_regfile_N255) );
  NOR2X1 U54163 ( .A(n44472), .B(n43104), .Y(n51581) );
  NOR2X1 U54164 ( .A(n44469), .B(n43107), .Y(n51580) );
  NOR2X1 U54165 ( .A(n51581), .B(n51580), .Y(n51583) );
  NOR2X1 U54166 ( .A(n21002), .B(n21001), .Y(n51582) );
  NAND2X1 U54167 ( .A(n51583), .B(n51582), .Y(u_decode_u_regfile_N440) );
  NOR2X1 U54168 ( .A(n44583), .B(n43104), .Y(n51585) );
  NOR2X1 U54169 ( .A(n44580), .B(n43107), .Y(n51584) );
  NOR2X1 U54170 ( .A(n51585), .B(n51584), .Y(n51587) );
  NOR2X1 U54171 ( .A(n18646), .B(n18645), .Y(n51586) );
  NAND2X1 U54172 ( .A(n51587), .B(n51586), .Y(u_decode_u_regfile_N884) );
  NOR2X1 U54173 ( .A(n44571), .B(n43104), .Y(n51589) );
  NOR2X1 U54174 ( .A(n44568), .B(n43107), .Y(n51588) );
  NOR2X1 U54175 ( .A(n51589), .B(n51588), .Y(n51591) );
  NOR2X1 U54176 ( .A(n19038), .B(n19037), .Y(n51590) );
  NAND2X1 U54177 ( .A(n51591), .B(n51590), .Y(u_decode_u_regfile_N810) );
  NOR2X1 U54178 ( .A(n44592), .B(n43104), .Y(n51593) );
  NOR2X1 U54179 ( .A(n44589), .B(n43107), .Y(n51592) );
  NOR2X1 U54180 ( .A(n51593), .B(n51592), .Y(n51595) );
  NOR2X1 U54181 ( .A(n18452), .B(n18451), .Y(n51594) );
  NAND2X1 U54182 ( .A(n51595), .B(n51594), .Y(u_decode_u_regfile_N921) );
  NOR2X1 U54183 ( .A(n44502), .B(n43104), .Y(n51597) );
  NOR2X1 U54184 ( .A(n44499), .B(n43107), .Y(n51596) );
  NOR2X1 U54185 ( .A(n51597), .B(n51596), .Y(n51599) );
  NOR2X1 U54186 ( .A(n20414), .B(n20413), .Y(n51598) );
  NAND2X1 U54187 ( .A(n51599), .B(n51598), .Y(u_decode_u_regfile_N551) );
  NOR2X1 U54188 ( .A(n44340), .B(n43104), .Y(n51601) );
  NOR2X1 U54189 ( .A(n44337), .B(n43107), .Y(n51600) );
  NOR2X1 U54190 ( .A(n51601), .B(n51600), .Y(n51603) );
  NOR2X1 U54191 ( .A(n23266), .B(n23265), .Y(n51602) );
  NAND2X1 U54192 ( .A(n51603), .B(n51602), .Y(u_decode_u_regfile_N1143) );
  NOR2X1 U54193 ( .A(n44352), .B(n43104), .Y(n51605) );
  NOR2X1 U54194 ( .A(n44349), .B(n43107), .Y(n51604) );
  NOR2X1 U54195 ( .A(n51605), .B(n51604), .Y(n51607) );
  NOR2X1 U54196 ( .A(n23046), .B(n23045), .Y(n51606) );
  NAND2X1 U54197 ( .A(n51607), .B(n51606), .Y(u_decode_u_regfile_N1180) );
  NOR2X1 U54198 ( .A(n44577), .B(n43104), .Y(n51609) );
  NOR2X1 U54199 ( .A(n44574), .B(n43107), .Y(n51608) );
  NOR2X1 U54200 ( .A(n51609), .B(n51608), .Y(n51611) );
  NOR2X1 U54201 ( .A(n18842), .B(n18841), .Y(n51610) );
  NAND2X1 U54202 ( .A(n51611), .B(n51610), .Y(u_decode_u_regfile_N847) );
  NOR2X1 U54203 ( .A(n44526), .B(n43104), .Y(n51613) );
  NOR2X1 U54204 ( .A(n44523), .B(n43106), .Y(n51612) );
  NOR2X1 U54205 ( .A(n51613), .B(n51612), .Y(n51615) );
  NOR2X1 U54206 ( .A(n20022), .B(n20021), .Y(n51614) );
  NAND2X1 U54207 ( .A(n51615), .B(n51614), .Y(u_decode_u_regfile_N625) );
  NOR2X1 U54208 ( .A(n44514), .B(n43104), .Y(n51617) );
  NOR2X1 U54209 ( .A(n44511), .B(n43106), .Y(n51616) );
  NOR2X1 U54210 ( .A(n51617), .B(n51616), .Y(n51619) );
  NOR2X1 U54211 ( .A(n20218), .B(n20217), .Y(n51618) );
  NAND2X1 U54212 ( .A(n51619), .B(n51618), .Y(u_decode_u_regfile_N588) );
  NOR2X1 U54213 ( .A(n43103), .B(n43276), .Y(n51621) );
  NOR2X1 U54214 ( .A(n43106), .B(n43385), .Y(n51620) );
  NOR2X1 U54215 ( .A(n51621), .B(n51620), .Y(n51623) );
  NOR2X1 U54216 ( .A(n20610), .B(n20609), .Y(n51622) );
  NAND2X1 U54217 ( .A(n51623), .B(n51622), .Y(u_decode_u_regfile_N514) );
  NOR2X1 U54218 ( .A(n44460), .B(n43103), .Y(n51625) );
  NOR2X1 U54219 ( .A(n44457), .B(n43106), .Y(n51624) );
  NOR2X1 U54220 ( .A(n51625), .B(n51624), .Y(n51627) );
  NOR2X1 U54221 ( .A(n21198), .B(n21197), .Y(n51626) );
  NAND2X1 U54222 ( .A(n51627), .B(n51626), .Y(u_decode_u_regfile_N403) );
  NOR2X1 U54223 ( .A(n19678), .B(n43103), .Y(n51629) );
  NOR2X1 U54224 ( .A(n44535), .B(n43106), .Y(n51628) );
  NOR2X1 U54225 ( .A(n51629), .B(n51628), .Y(n51631) );
  NOR2X1 U54226 ( .A(n19825), .B(n19824), .Y(n51630) );
  NAND2X1 U54227 ( .A(n51631), .B(n51630), .Y(u_decode_u_regfile_N662) );
  NOR2X1 U54228 ( .A(n44550), .B(n43104), .Y(n51633) );
  NOR2X1 U54229 ( .A(n44547), .B(n43107), .Y(n51632) );
  NOR2X1 U54230 ( .A(n51633), .B(n51632), .Y(n51635) );
  NOR2X1 U54231 ( .A(n19628), .B(n19627), .Y(n51634) );
  NAND2X1 U54232 ( .A(n51635), .B(n51634), .Y(u_decode_u_regfile_N699) );
  NOR2X1 U54233 ( .A(n44565), .B(n43103), .Y(n51637) );
  NOR2X1 U54234 ( .A(n44562), .B(n43106), .Y(n51636) );
  NOR2X1 U54235 ( .A(n51637), .B(n51636), .Y(n51639) );
  NOR2X1 U54236 ( .A(n19234), .B(n19233), .Y(n51638) );
  NAND2X1 U54237 ( .A(n51639), .B(n51638), .Y(u_decode_u_regfile_N773) );
  NOR2X1 U54238 ( .A(n44394), .B(n43103), .Y(n51641) );
  NOR2X1 U54239 ( .A(n44391), .B(n43106), .Y(n51640) );
  NOR2X1 U54240 ( .A(n51641), .B(n51640), .Y(n51643) );
  NOR2X1 U54241 ( .A(n22376), .B(n22375), .Y(n51642) );
  NAND2X1 U54242 ( .A(n51643), .B(n51642), .Y(u_decode_u_regfile_N181) );
  NOR2X1 U54243 ( .A(n44316), .B(n43104), .Y(n51645) );
  NOR2X1 U54244 ( .A(n44313), .B(n43106), .Y(n51644) );
  NOR2X1 U54245 ( .A(n51645), .B(n51644), .Y(n51647) );
  NOR2X1 U54246 ( .A(n23706), .B(n23705), .Y(n51646) );
  NAND2X1 U54247 ( .A(n51647), .B(n51646), .Y(u_decode_u_regfile_N1069) );
  NOR2X1 U54248 ( .A(n44484), .B(n43103), .Y(n51649) );
  NOR2X1 U54249 ( .A(n44481), .B(n43106), .Y(n51648) );
  NOR2X1 U54250 ( .A(n51649), .B(n51648), .Y(n51651) );
  NOR2X1 U54251 ( .A(n20806), .B(n20805), .Y(n51650) );
  NAND2X1 U54252 ( .A(n51651), .B(n51650), .Y(u_decode_u_regfile_N477) );
  NOR2X1 U54253 ( .A(n44601), .B(n43103), .Y(n51653) );
  NOR2X1 U54254 ( .A(n44598), .B(n43106), .Y(n51652) );
  NOR2X1 U54255 ( .A(n51653), .B(n51652), .Y(n51655) );
  NOR2X1 U54256 ( .A(n18253), .B(n18252), .Y(n51654) );
  NAND2X1 U54257 ( .A(n51655), .B(n51654), .Y(u_decode_u_regfile_N958) );
  NOR2X1 U54258 ( .A(n44607), .B(n43103), .Y(n51657) );
  NOR2X1 U54259 ( .A(n44604), .B(n43106), .Y(n51656) );
  NOR2X1 U54260 ( .A(n51657), .B(n51656), .Y(n51659) );
  NOR2X1 U54261 ( .A(n18032), .B(n18030), .Y(n51658) );
  NAND2X1 U54262 ( .A(n51659), .B(n51658), .Y(u_decode_u_regfile_N995) );
  NOR2X1 U54263 ( .A(n43103), .B(n43273), .Y(n51661) );
  NOR2X1 U54264 ( .A(n43106), .B(n43391), .Y(n51660) );
  NOR2X1 U54265 ( .A(n51661), .B(n51660), .Y(n51663) );
  NOR2X1 U54266 ( .A(n23700), .B(n23699), .Y(n51662) );
  NAND2X1 U54267 ( .A(n51663), .B(n51662), .Y(u_decode_u_regfile_N107) );
  NOR2X1 U54268 ( .A(n43103), .B(n43270), .Y(n51665) );
  NOR2X1 U54269 ( .A(n43106), .B(n43388), .Y(n51664) );
  NOR2X1 U54270 ( .A(n51665), .B(n51664), .Y(n51667) );
  NOR2X1 U54271 ( .A(n21395), .B(n21394), .Y(n51666) );
  NAND2X1 U54272 ( .A(n51667), .B(n51666), .Y(u_decode_u_regfile_N366) );
  NOR2X1 U54273 ( .A(n15561), .B(n15562), .Y(n51669) );
  NOR2X1 U54274 ( .A(n15596), .B(n15597), .Y(n51668) );
  NAND2X1 U54275 ( .A(n51669), .B(n51668), .Y(u_exec_alu_p_w[6]) );
  NOR2X1 U54276 ( .A(n44364), .B(n43108), .Y(n51671) );
  NOR2X1 U54277 ( .A(n44361), .B(n43111), .Y(n51670) );
  NOR2X1 U54278 ( .A(n51671), .B(n51670), .Y(n51673) );
  NOR2X1 U54279 ( .A(n22838), .B(n22837), .Y(n51672) );
  NAND2X1 U54280 ( .A(n51673), .B(n51672), .Y(u_decode_u_regfile_N1216) );
  NOR2X1 U54281 ( .A(n44442), .B(n43110), .Y(n51675) );
  NOR2X1 U54282 ( .A(n44439), .B(n37667), .Y(n51674) );
  NOR2X1 U54283 ( .A(n51675), .B(n51674), .Y(n51677) );
  NOR2X1 U54284 ( .A(n21598), .B(n21597), .Y(n51676) );
  NAND2X1 U54285 ( .A(n51677), .B(n51676), .Y(u_decode_u_regfile_N328) );
  NOR2X1 U54286 ( .A(n44382), .B(n43110), .Y(n51679) );
  NOR2X1 U54287 ( .A(n44379), .B(n37667), .Y(n51678) );
  NOR2X1 U54288 ( .A(n51679), .B(n51678), .Y(n51681) );
  NOR2X1 U54289 ( .A(n22578), .B(n22577), .Y(n51680) );
  NAND2X1 U54290 ( .A(n51681), .B(n51680), .Y(u_decode_u_regfile_N143) );
  NOR2X1 U54291 ( .A(n44304), .B(n43110), .Y(n51683) );
  NOR2X1 U54292 ( .A(n44301), .B(n37667), .Y(n51682) );
  NOR2X1 U54293 ( .A(n51683), .B(n51682), .Y(n51685) );
  NOR2X1 U54294 ( .A(n23926), .B(n23925), .Y(n51684) );
  NAND2X1 U54295 ( .A(n51685), .B(n51684), .Y(u_decode_u_regfile_N1031) );
  NOR2X1 U54296 ( .A(n44406), .B(n43110), .Y(n51687) );
  NOR2X1 U54297 ( .A(n44403), .B(n43112), .Y(n51686) );
  NOR2X1 U54298 ( .A(n51687), .B(n51686), .Y(n51689) );
  NOR2X1 U54299 ( .A(n22186), .B(n22185), .Y(n51688) );
  NAND2X1 U54300 ( .A(n51689), .B(n51688), .Y(u_decode_u_regfile_N217) );
  NOR2X1 U54301 ( .A(n44559), .B(n43109), .Y(n51691) );
  NOR2X1 U54302 ( .A(n44556), .B(n43112), .Y(n51690) );
  NOR2X1 U54303 ( .A(n51691), .B(n51690), .Y(n51693) );
  NOR2X1 U54304 ( .A(n19436), .B(n19435), .Y(n51692) );
  NAND2X1 U54305 ( .A(n51693), .B(n51692), .Y(u_decode_u_regfile_N735) );
  NOR2X1 U54306 ( .A(n44328), .B(n43109), .Y(n51695) );
  NOR2X1 U54307 ( .A(n44325), .B(n43112), .Y(n51694) );
  NOR2X1 U54308 ( .A(n51695), .B(n51694), .Y(n51697) );
  NOR2X1 U54309 ( .A(n23492), .B(n23491), .Y(n51696) );
  NAND2X1 U54310 ( .A(n51697), .B(n51696), .Y(u_decode_u_regfile_N1105) );
  NOR2X1 U54311 ( .A(n44430), .B(n43109), .Y(n51699) );
  NOR2X1 U54312 ( .A(n44427), .B(n43112), .Y(n51698) );
  NOR2X1 U54313 ( .A(n51699), .B(n51698), .Y(n51701) );
  NOR2X1 U54314 ( .A(n21794), .B(n21793), .Y(n51700) );
  NAND2X1 U54315 ( .A(n51701), .B(n51700), .Y(u_decode_u_regfile_N291) );
  NOR2X1 U54316 ( .A(n44418), .B(n43109), .Y(n51703) );
  NOR2X1 U54317 ( .A(n44415), .B(n43112), .Y(n51702) );
  NOR2X1 U54318 ( .A(n51703), .B(n51702), .Y(n51705) );
  NOR2X1 U54319 ( .A(n21990), .B(n21989), .Y(n51704) );
  NAND2X1 U54320 ( .A(n51705), .B(n51704), .Y(u_decode_u_regfile_N254) );
  NOR2X1 U54321 ( .A(n44472), .B(n43109), .Y(n51707) );
  NOR2X1 U54322 ( .A(n44469), .B(n43112), .Y(n51706) );
  NOR2X1 U54323 ( .A(n51707), .B(n51706), .Y(n51709) );
  NOR2X1 U54324 ( .A(n21008), .B(n21007), .Y(n51708) );
  NAND2X1 U54325 ( .A(n51709), .B(n51708), .Y(u_decode_u_regfile_N439) );
  NOR2X1 U54326 ( .A(n44583), .B(n43109), .Y(n51711) );
  NOR2X1 U54327 ( .A(n44580), .B(n43112), .Y(n51710) );
  NOR2X1 U54328 ( .A(n51711), .B(n51710), .Y(n51713) );
  NOR2X1 U54329 ( .A(n18652), .B(n18651), .Y(n51712) );
  NAND2X1 U54330 ( .A(n51713), .B(n51712), .Y(u_decode_u_regfile_N883) );
  NOR2X1 U54331 ( .A(n44571), .B(n43109), .Y(n51715) );
  NOR2X1 U54332 ( .A(n44568), .B(n43112), .Y(n51714) );
  NOR2X1 U54333 ( .A(n51715), .B(n51714), .Y(n51717) );
  NOR2X1 U54334 ( .A(n19044), .B(n19043), .Y(n51716) );
  NAND2X1 U54335 ( .A(n51717), .B(n51716), .Y(u_decode_u_regfile_N809) );
  NOR2X1 U54336 ( .A(n44592), .B(n43109), .Y(n51719) );
  NOR2X1 U54337 ( .A(n44589), .B(n43112), .Y(n51718) );
  NOR2X1 U54338 ( .A(n51719), .B(n51718), .Y(n51721) );
  NOR2X1 U54339 ( .A(n18458), .B(n18457), .Y(n51720) );
  NAND2X1 U54340 ( .A(n51721), .B(n51720), .Y(u_decode_u_regfile_N920) );
  NOR2X1 U54341 ( .A(n44502), .B(n43109), .Y(n51723) );
  NOR2X1 U54342 ( .A(n44499), .B(n43112), .Y(n51722) );
  NOR2X1 U54343 ( .A(n51723), .B(n51722), .Y(n51725) );
  NOR2X1 U54344 ( .A(n20420), .B(n20419), .Y(n51724) );
  NAND2X1 U54345 ( .A(n51725), .B(n51724), .Y(u_decode_u_regfile_N550) );
  NOR2X1 U54346 ( .A(n44340), .B(n43109), .Y(n51727) );
  NOR2X1 U54347 ( .A(n44337), .B(n43112), .Y(n51726) );
  NOR2X1 U54348 ( .A(n51727), .B(n51726), .Y(n51729) );
  NOR2X1 U54349 ( .A(n23272), .B(n23271), .Y(n51728) );
  NAND2X1 U54350 ( .A(n51729), .B(n51728), .Y(u_decode_u_regfile_N1142) );
  NOR2X1 U54351 ( .A(n44352), .B(n43109), .Y(n51731) );
  NOR2X1 U54352 ( .A(n44349), .B(n43112), .Y(n51730) );
  NOR2X1 U54353 ( .A(n51731), .B(n51730), .Y(n51733) );
  NOR2X1 U54354 ( .A(n23058), .B(n23057), .Y(n51732) );
  NAND2X1 U54355 ( .A(n51733), .B(n51732), .Y(u_decode_u_regfile_N1179) );
  NOR2X1 U54356 ( .A(n44577), .B(n43109), .Y(n51735) );
  NOR2X1 U54357 ( .A(n44574), .B(n43112), .Y(n51734) );
  NOR2X1 U54358 ( .A(n51735), .B(n51734), .Y(n51737) );
  NOR2X1 U54359 ( .A(n18848), .B(n18847), .Y(n51736) );
  NAND2X1 U54360 ( .A(n51737), .B(n51736), .Y(u_decode_u_regfile_N846) );
  NOR2X1 U54361 ( .A(n44526), .B(n43109), .Y(n51739) );
  NOR2X1 U54362 ( .A(n44523), .B(n43111), .Y(n51738) );
  NOR2X1 U54363 ( .A(n51739), .B(n51738), .Y(n51741) );
  NOR2X1 U54364 ( .A(n20028), .B(n20027), .Y(n51740) );
  NAND2X1 U54365 ( .A(n51741), .B(n51740), .Y(u_decode_u_regfile_N624) );
  NOR2X1 U54366 ( .A(n44514), .B(n43108), .Y(n51743) );
  NOR2X1 U54367 ( .A(n44511), .B(n43111), .Y(n51742) );
  NOR2X1 U54368 ( .A(n51743), .B(n51742), .Y(n51745) );
  NOR2X1 U54369 ( .A(n20224), .B(n20223), .Y(n51744) );
  NAND2X1 U54370 ( .A(n51745), .B(n51744), .Y(u_decode_u_regfile_N587) );
  NOR2X1 U54371 ( .A(n43108), .B(n43276), .Y(n51747) );
  NOR2X1 U54372 ( .A(n43111), .B(n43384), .Y(n51746) );
  NOR2X1 U54373 ( .A(n51747), .B(n51746), .Y(n51749) );
  NOR2X1 U54374 ( .A(n20616), .B(n20615), .Y(n51748) );
  NAND2X1 U54375 ( .A(n51749), .B(n51748), .Y(u_decode_u_regfile_N513) );
  NOR2X1 U54376 ( .A(n44460), .B(n43108), .Y(n51751) );
  NOR2X1 U54377 ( .A(n44457), .B(n43111), .Y(n51750) );
  NOR2X1 U54378 ( .A(n51751), .B(n51750), .Y(n51753) );
  NOR2X1 U54379 ( .A(n21204), .B(n21203), .Y(n51752) );
  NAND2X1 U54380 ( .A(n51753), .B(n51752), .Y(u_decode_u_regfile_N402) );
  NOR2X1 U54381 ( .A(n19678), .B(n43108), .Y(n51755) );
  NOR2X1 U54382 ( .A(n44535), .B(n43111), .Y(n51754) );
  NOR2X1 U54383 ( .A(n51755), .B(n51754), .Y(n51757) );
  NOR2X1 U54384 ( .A(n19831), .B(n19830), .Y(n51756) );
  NAND2X1 U54385 ( .A(n51757), .B(n51756), .Y(u_decode_u_regfile_N661) );
  NOR2X1 U54386 ( .A(n44550), .B(n43109), .Y(n51759) );
  NOR2X1 U54387 ( .A(n44547), .B(n43111), .Y(n51758) );
  NOR2X1 U54388 ( .A(n51759), .B(n51758), .Y(n51761) );
  NOR2X1 U54389 ( .A(n19634), .B(n19633), .Y(n51760) );
  NAND2X1 U54390 ( .A(n51761), .B(n51760), .Y(u_decode_u_regfile_N698) );
  NOR2X1 U54391 ( .A(n44565), .B(n43108), .Y(n51763) );
  NOR2X1 U54392 ( .A(n44562), .B(n43111), .Y(n51762) );
  NOR2X1 U54393 ( .A(n51763), .B(n51762), .Y(n51765) );
  NOR2X1 U54394 ( .A(n19240), .B(n19239), .Y(n51764) );
  NAND2X1 U54395 ( .A(n51765), .B(n51764), .Y(u_decode_u_regfile_N772) );
  NOR2X1 U54396 ( .A(n44394), .B(n43108), .Y(n51767) );
  NOR2X1 U54397 ( .A(n44391), .B(n43112), .Y(n51766) );
  NOR2X1 U54398 ( .A(n51767), .B(n51766), .Y(n51769) );
  NOR2X1 U54399 ( .A(n22382), .B(n22381), .Y(n51768) );
  NAND2X1 U54400 ( .A(n51769), .B(n51768), .Y(u_decode_u_regfile_N180) );
  NOR2X1 U54401 ( .A(n44316), .B(n43108), .Y(n51771) );
  NOR2X1 U54402 ( .A(n44313), .B(n43111), .Y(n51770) );
  NOR2X1 U54403 ( .A(n51771), .B(n51770), .Y(n51773) );
  NOR2X1 U54404 ( .A(n23712), .B(n23711), .Y(n51772) );
  NAND2X1 U54405 ( .A(n51773), .B(n51772), .Y(u_decode_u_regfile_N1068) );
  NOR2X1 U54406 ( .A(n44484), .B(n43108), .Y(n51775) );
  NOR2X1 U54407 ( .A(n44481), .B(n43111), .Y(n51774) );
  NOR2X1 U54408 ( .A(n51775), .B(n51774), .Y(n51777) );
  NOR2X1 U54409 ( .A(n20812), .B(n20811), .Y(n51776) );
  NAND2X1 U54410 ( .A(n51777), .B(n51776), .Y(u_decode_u_regfile_N476) );
  NOR2X1 U54411 ( .A(n44601), .B(n43108), .Y(n51779) );
  NOR2X1 U54412 ( .A(n44598), .B(n43111), .Y(n51778) );
  NOR2X1 U54413 ( .A(n51779), .B(n51778), .Y(n51781) );
  NOR2X1 U54414 ( .A(n18259), .B(n18258), .Y(n51780) );
  NAND2X1 U54415 ( .A(n51781), .B(n51780), .Y(u_decode_u_regfile_N957) );
  NOR2X1 U54416 ( .A(n44607), .B(n43108), .Y(n51783) );
  NOR2X1 U54417 ( .A(n44604), .B(n43111), .Y(n51782) );
  NOR2X1 U54418 ( .A(n51783), .B(n51782), .Y(n51785) );
  NOR2X1 U54419 ( .A(n18039), .B(n18037), .Y(n51784) );
  NAND2X1 U54420 ( .A(n51785), .B(n51784), .Y(u_decode_u_regfile_N994) );
  NOR2X1 U54421 ( .A(n43108), .B(n43273), .Y(n51787) );
  NOR2X1 U54422 ( .A(n43111), .B(n43390), .Y(n51786) );
  NOR2X1 U54423 ( .A(n51787), .B(n51786), .Y(n51789) );
  NOR2X1 U54424 ( .A(n23754), .B(n23753), .Y(n51788) );
  NAND2X1 U54425 ( .A(n51789), .B(n51788), .Y(u_decode_u_regfile_N106) );
  NOR2X1 U54426 ( .A(n43108), .B(n43270), .Y(n51791) );
  NOR2X1 U54427 ( .A(n43111), .B(n43387), .Y(n51790) );
  NOR2X1 U54428 ( .A(n51791), .B(n51790), .Y(n51793) );
  NOR2X1 U54429 ( .A(n21401), .B(n21400), .Y(n51792) );
  NAND2X1 U54430 ( .A(n51793), .B(n51792), .Y(u_decode_u_regfile_N365) );
  NOR2X1 U54431 ( .A(n15613), .B(n15614), .Y(n51795) );
  NOR2X1 U54432 ( .A(n15650), .B(n15651), .Y(n51794) );
  NAND2X1 U54433 ( .A(n51795), .B(n51794), .Y(u_exec_alu_p_w[5]) );
  NOR2X1 U54434 ( .A(n44364), .B(n43114), .Y(n51797) );
  NOR2X1 U54435 ( .A(n44361), .B(n43117), .Y(n51796) );
  NOR2X1 U54436 ( .A(n51797), .B(n51796), .Y(n51799) );
  NOR2X1 U54437 ( .A(n22844), .B(n22843), .Y(n51798) );
  NAND2X1 U54438 ( .A(n51799), .B(n51798), .Y(u_decode_u_regfile_N1215) );
  NOR2X1 U54439 ( .A(n44442), .B(n43116), .Y(n51801) );
  NOR2X1 U54440 ( .A(n44439), .B(n37668), .Y(n51800) );
  NOR2X1 U54441 ( .A(n51801), .B(n51800), .Y(n51803) );
  NOR2X1 U54442 ( .A(n21604), .B(n21603), .Y(n51802) );
  NAND2X1 U54443 ( .A(n51803), .B(n51802), .Y(u_decode_u_regfile_N327) );
  NOR2X1 U54444 ( .A(n44382), .B(n43116), .Y(n51805) );
  NOR2X1 U54445 ( .A(n44379), .B(n37668), .Y(n51804) );
  NOR2X1 U54446 ( .A(n51805), .B(n51804), .Y(n51807) );
  NOR2X1 U54447 ( .A(n22584), .B(n22583), .Y(n51806) );
  NAND2X1 U54448 ( .A(n51807), .B(n51806), .Y(u_decode_u_regfile_N142) );
  NOR2X1 U54449 ( .A(n44304), .B(n43116), .Y(n51809) );
  NOR2X1 U54450 ( .A(n44301), .B(n37668), .Y(n51808) );
  NOR2X1 U54451 ( .A(n51809), .B(n51808), .Y(n51811) );
  NOR2X1 U54452 ( .A(n23932), .B(n23931), .Y(n51810) );
  NAND2X1 U54453 ( .A(n51811), .B(n51810), .Y(u_decode_u_regfile_N1030) );
  NOR2X1 U54454 ( .A(n44406), .B(n43116), .Y(n51813) );
  NOR2X1 U54455 ( .A(n44403), .B(n43118), .Y(n51812) );
  NOR2X1 U54456 ( .A(n51813), .B(n51812), .Y(n51815) );
  NOR2X1 U54457 ( .A(n22192), .B(n22191), .Y(n51814) );
  NAND2X1 U54458 ( .A(n51815), .B(n51814), .Y(u_decode_u_regfile_N216) );
  NOR2X1 U54459 ( .A(n44559), .B(n43115), .Y(n51817) );
  NOR2X1 U54460 ( .A(n44556), .B(n43118), .Y(n51816) );
  NOR2X1 U54461 ( .A(n51817), .B(n51816), .Y(n51819) );
  NOR2X1 U54462 ( .A(n19442), .B(n19441), .Y(n51818) );
  NAND2X1 U54463 ( .A(n51819), .B(n51818), .Y(u_decode_u_regfile_N734) );
  NOR2X1 U54464 ( .A(n44328), .B(n43115), .Y(n51821) );
  NOR2X1 U54465 ( .A(n44325), .B(n43118), .Y(n51820) );
  NOR2X1 U54466 ( .A(n51821), .B(n51820), .Y(n51823) );
  NOR2X1 U54467 ( .A(n23498), .B(n23497), .Y(n51822) );
  NAND2X1 U54468 ( .A(n51823), .B(n51822), .Y(u_decode_u_regfile_N1104) );
  NOR2X1 U54469 ( .A(n44430), .B(n43115), .Y(n51825) );
  NOR2X1 U54470 ( .A(n44427), .B(n43118), .Y(n51824) );
  NOR2X1 U54471 ( .A(n51825), .B(n51824), .Y(n51827) );
  NOR2X1 U54472 ( .A(n21800), .B(n21799), .Y(n51826) );
  NAND2X1 U54473 ( .A(n51827), .B(n51826), .Y(u_decode_u_regfile_N290) );
  NOR2X1 U54474 ( .A(n44418), .B(n43115), .Y(n51829) );
  NOR2X1 U54475 ( .A(n44415), .B(n43118), .Y(n51828) );
  NOR2X1 U54476 ( .A(n51829), .B(n51828), .Y(n51831) );
  NOR2X1 U54477 ( .A(n21996), .B(n21995), .Y(n51830) );
  NAND2X1 U54478 ( .A(n51831), .B(n51830), .Y(u_decode_u_regfile_N253) );
  NOR2X1 U54479 ( .A(n44472), .B(n43115), .Y(n51833) );
  NOR2X1 U54480 ( .A(n44469), .B(n43118), .Y(n51832) );
  NOR2X1 U54481 ( .A(n51833), .B(n51832), .Y(n51835) );
  NOR2X1 U54482 ( .A(n21014), .B(n21013), .Y(n51834) );
  NAND2X1 U54483 ( .A(n51835), .B(n51834), .Y(u_decode_u_regfile_N438) );
  NOR2X1 U54484 ( .A(n44583), .B(n43115), .Y(n51837) );
  NOR2X1 U54485 ( .A(n44580), .B(n43118), .Y(n51836) );
  NOR2X1 U54486 ( .A(n51837), .B(n51836), .Y(n51839) );
  NOR2X1 U54487 ( .A(n18658), .B(n18657), .Y(n51838) );
  NAND2X1 U54488 ( .A(n51839), .B(n51838), .Y(u_decode_u_regfile_N882) );
  NOR2X1 U54489 ( .A(n44571), .B(n43115), .Y(n51841) );
  NOR2X1 U54490 ( .A(n44568), .B(n43118), .Y(n51840) );
  NOR2X1 U54491 ( .A(n51841), .B(n51840), .Y(n51843) );
  NOR2X1 U54492 ( .A(n19050), .B(n19049), .Y(n51842) );
  NAND2X1 U54493 ( .A(n51843), .B(n51842), .Y(u_decode_u_regfile_N808) );
  NOR2X1 U54494 ( .A(n44592), .B(n43115), .Y(n51845) );
  NOR2X1 U54495 ( .A(n44589), .B(n43118), .Y(n51844) );
  NOR2X1 U54496 ( .A(n51845), .B(n51844), .Y(n51847) );
  NOR2X1 U54497 ( .A(n18464), .B(n18463), .Y(n51846) );
  NAND2X1 U54498 ( .A(n51847), .B(n51846), .Y(u_decode_u_regfile_N919) );
  NOR2X1 U54499 ( .A(n44502), .B(n43115), .Y(n51849) );
  NOR2X1 U54500 ( .A(n44499), .B(n43118), .Y(n51848) );
  NOR2X1 U54501 ( .A(n51849), .B(n51848), .Y(n51851) );
  NOR2X1 U54502 ( .A(n20426), .B(n20425), .Y(n51850) );
  NAND2X1 U54503 ( .A(n51851), .B(n51850), .Y(u_decode_u_regfile_N549) );
  NOR2X1 U54504 ( .A(n44340), .B(n43115), .Y(n51853) );
  NOR2X1 U54505 ( .A(n44337), .B(n43118), .Y(n51852) );
  NOR2X1 U54506 ( .A(n51853), .B(n51852), .Y(n51855) );
  NOR2X1 U54507 ( .A(n23278), .B(n23277), .Y(n51854) );
  NAND2X1 U54508 ( .A(n51855), .B(n51854), .Y(u_decode_u_regfile_N1141) );
  NOR2X1 U54509 ( .A(n44352), .B(n43115), .Y(n51857) );
  NOR2X1 U54510 ( .A(n44349), .B(n43118), .Y(n51856) );
  NOR2X1 U54511 ( .A(n51857), .B(n51856), .Y(n51859) );
  NOR2X1 U54512 ( .A(n23064), .B(n23063), .Y(n51858) );
  NAND2X1 U54513 ( .A(n51859), .B(n51858), .Y(u_decode_u_regfile_N1178) );
  NOR2X1 U54514 ( .A(n44577), .B(n43115), .Y(n51861) );
  NOR2X1 U54515 ( .A(n44574), .B(n43118), .Y(n51860) );
  NOR2X1 U54516 ( .A(n51861), .B(n51860), .Y(n51863) );
  NOR2X1 U54517 ( .A(n18854), .B(n18853), .Y(n51862) );
  NAND2X1 U54518 ( .A(n51863), .B(n51862), .Y(u_decode_u_regfile_N845) );
  NOR2X1 U54519 ( .A(n44526), .B(n43115), .Y(n51865) );
  NOR2X1 U54520 ( .A(n44523), .B(n43117), .Y(n51864) );
  NOR2X1 U54521 ( .A(n51865), .B(n51864), .Y(n51867) );
  NOR2X1 U54522 ( .A(n20034), .B(n20033), .Y(n51866) );
  NAND2X1 U54523 ( .A(n51867), .B(n51866), .Y(u_decode_u_regfile_N623) );
  NOR2X1 U54524 ( .A(n44514), .B(n43114), .Y(n51869) );
  NOR2X1 U54525 ( .A(n44511), .B(n43117), .Y(n51868) );
  NOR2X1 U54526 ( .A(n51869), .B(n51868), .Y(n51871) );
  NOR2X1 U54527 ( .A(n20230), .B(n20229), .Y(n51870) );
  NAND2X1 U54528 ( .A(n51871), .B(n51870), .Y(u_decode_u_regfile_N586) );
  NOR2X1 U54529 ( .A(n43114), .B(n43276), .Y(n51873) );
  NOR2X1 U54530 ( .A(n43117), .B(n43384), .Y(n51872) );
  NOR2X1 U54531 ( .A(n51873), .B(n51872), .Y(n51875) );
  NOR2X1 U54532 ( .A(n20622), .B(n20621), .Y(n51874) );
  NAND2X1 U54533 ( .A(n51875), .B(n51874), .Y(u_decode_u_regfile_N512) );
  NOR2X1 U54534 ( .A(n44460), .B(n43114), .Y(n51877) );
  NOR2X1 U54535 ( .A(n44457), .B(n43117), .Y(n51876) );
  NOR2X1 U54536 ( .A(n51877), .B(n51876), .Y(n51879) );
  NOR2X1 U54537 ( .A(n21210), .B(n21209), .Y(n51878) );
  NAND2X1 U54538 ( .A(n51879), .B(n51878), .Y(u_decode_u_regfile_N401) );
  NOR2X1 U54539 ( .A(n19678), .B(n43114), .Y(n51881) );
  NOR2X1 U54540 ( .A(n44535), .B(n43117), .Y(n51880) );
  NOR2X1 U54541 ( .A(n51881), .B(n51880), .Y(n51883) );
  NOR2X1 U54542 ( .A(n19837), .B(n19836), .Y(n51882) );
  NAND2X1 U54543 ( .A(n51883), .B(n51882), .Y(u_decode_u_regfile_N660) );
  NOR2X1 U54544 ( .A(n44550), .B(n43115), .Y(n51885) );
  NOR2X1 U54545 ( .A(n44547), .B(n43117), .Y(n51884) );
  NOR2X1 U54546 ( .A(n51885), .B(n51884), .Y(n51887) );
  NOR2X1 U54547 ( .A(n19640), .B(n19639), .Y(n51886) );
  NAND2X1 U54548 ( .A(n51887), .B(n51886), .Y(u_decode_u_regfile_N697) );
  NOR2X1 U54549 ( .A(n44565), .B(n43114), .Y(n51889) );
  NOR2X1 U54550 ( .A(n44562), .B(n43117), .Y(n51888) );
  NOR2X1 U54551 ( .A(n51889), .B(n51888), .Y(n51891) );
  NOR2X1 U54552 ( .A(n19246), .B(n19245), .Y(n51890) );
  NAND2X1 U54553 ( .A(n51891), .B(n51890), .Y(u_decode_u_regfile_N771) );
  NOR2X1 U54554 ( .A(n44394), .B(n43114), .Y(n51893) );
  NOR2X1 U54555 ( .A(n44391), .B(n43118), .Y(n51892) );
  NOR2X1 U54556 ( .A(n51893), .B(n51892), .Y(n51895) );
  NOR2X1 U54557 ( .A(n22388), .B(n22387), .Y(n51894) );
  NAND2X1 U54558 ( .A(n51895), .B(n51894), .Y(u_decode_u_regfile_N179) );
  NOR2X1 U54559 ( .A(n44316), .B(n43114), .Y(n51897) );
  NOR2X1 U54560 ( .A(n44313), .B(n43117), .Y(n51896) );
  NOR2X1 U54561 ( .A(n51897), .B(n51896), .Y(n51899) );
  NOR2X1 U54562 ( .A(n23718), .B(n23717), .Y(n51898) );
  NAND2X1 U54563 ( .A(n51899), .B(n51898), .Y(u_decode_u_regfile_N1067) );
  NOR2X1 U54564 ( .A(n44484), .B(n43114), .Y(n51901) );
  NOR2X1 U54565 ( .A(n44481), .B(n43117), .Y(n51900) );
  NOR2X1 U54566 ( .A(n51901), .B(n51900), .Y(n51903) );
  NOR2X1 U54567 ( .A(n20818), .B(n20817), .Y(n51902) );
  NAND2X1 U54568 ( .A(n51903), .B(n51902), .Y(u_decode_u_regfile_N475) );
  NOR2X1 U54569 ( .A(n44601), .B(n43114), .Y(n51905) );
  NOR2X1 U54570 ( .A(n44598), .B(n43117), .Y(n51904) );
  NOR2X1 U54571 ( .A(n51905), .B(n51904), .Y(n51907) );
  NOR2X1 U54572 ( .A(n18265), .B(n18264), .Y(n51906) );
  NAND2X1 U54573 ( .A(n51907), .B(n51906), .Y(u_decode_u_regfile_N956) );
  NOR2X1 U54574 ( .A(n44607), .B(n43114), .Y(n51909) );
  NOR2X1 U54575 ( .A(n44604), .B(n43117), .Y(n51908) );
  NOR2X1 U54576 ( .A(n51909), .B(n51908), .Y(n51911) );
  NOR2X1 U54577 ( .A(n18046), .B(n18044), .Y(n51910) );
  NAND2X1 U54578 ( .A(n51911), .B(n51910), .Y(u_decode_u_regfile_N993) );
  NOR2X1 U54579 ( .A(n43114), .B(n43273), .Y(n51913) );
  NOR2X1 U54580 ( .A(n43117), .B(n43390), .Y(n51912) );
  NOR2X1 U54581 ( .A(n51913), .B(n51912), .Y(n51915) );
  NOR2X1 U54582 ( .A(n23806), .B(n23805), .Y(n51914) );
  NAND2X1 U54583 ( .A(n51915), .B(n51914), .Y(u_decode_u_regfile_N105) );
  NOR2X1 U54584 ( .A(n43114), .B(n43270), .Y(n51917) );
  NOR2X1 U54585 ( .A(n43117), .B(n43387), .Y(n51916) );
  NOR2X1 U54586 ( .A(n51917), .B(n51916), .Y(n51919) );
  NOR2X1 U54587 ( .A(n21407), .B(n21406), .Y(n51918) );
  NAND2X1 U54588 ( .A(n51919), .B(n51918), .Y(u_decode_u_regfile_N364) );
  INVX1 U54589 ( .A(n16631), .Y(n73573) );
  NAND2X1 U54590 ( .A(n42310), .B(n73573), .Y(n15463) );
  NAND2X1 U54591 ( .A(n42947), .B(n58576), .Y(n364) );
  MX2X1 U54592 ( .A(n42727), .B(n43461), .S0(n73522), .Y(n26014) );
  NAND2X1 U54593 ( .A(n44281), .B(n26014), .Y(n26331) );
  NAND2X1 U54594 ( .A(opcode_opcode_w[26]), .B(opcode_opcode_w[29]), .Y(n51920) );
  NOR2X1 U54595 ( .A(n51979), .B(n51920), .Y(n51922) );
  NOR2X1 U54596 ( .A(n42747), .B(opcode_opcode_w[27]), .Y(n51921) );
  NAND2X1 U54597 ( .A(n51922), .B(n51921), .Y(n24943) );
  XNOR2X1 U54598 ( .A(n51924), .B(n51923), .Y(n51925) );
  XOR2X1 U54599 ( .A(n51926), .B(n51925), .Y(n51927) );
  NOR2X1 U54600 ( .A(n51927), .B(n42930), .Y(n51931) );
  NOR2X1 U54601 ( .A(opcode_pc_w[1]), .B(opcode_opcode_w[8]), .Y(n51929) );
  NAND2X1 U54602 ( .A(opcode_opcode_w[8]), .B(opcode_pc_w[1]), .Y(n54448) );
  NAND2X1 U54603 ( .A(n54897), .B(n54448), .Y(n51928) );
  NOR2X1 U54604 ( .A(n51929), .B(n51928), .Y(n51930) );
  NOR2X1 U54605 ( .A(n51931), .B(n51930), .Y(n51935) );
  NAND2X1 U54606 ( .A(opcode_pc_w[1]), .B(n40453), .Y(n54387) );
  INVX1 U54607 ( .A(n54387), .Y(n54465) );
  NOR2X1 U54608 ( .A(n37342), .B(n54465), .Y(n51933) );
  NAND2X1 U54609 ( .A(n42468), .B(n56782), .Y(n51932) );
  NAND2X1 U54610 ( .A(n51933), .B(n51932), .Y(n51934) );
  NAND2X1 U54611 ( .A(n51935), .B(n51934), .Y(n56773) );
  INVX1 U54612 ( .A(n56773), .Y(n51938) );
  INVX1 U54613 ( .A(n26976), .Y(n51936) );
  NAND2X1 U54614 ( .A(n28560), .B(n73544), .Y(n51937) );
  NAND2X1 U54615 ( .A(n51937), .B(n26138), .Y(n72842) );
  INVX1 U54616 ( .A(n72842), .Y(n51941) );
  NAND2X1 U54617 ( .A(n51941), .B(n42439), .Y(n51967) );
  NOR2X1 U54618 ( .A(n51938), .B(n57240), .Y(n51948) );
  NAND2X1 U54619 ( .A(n72840), .B(n73544), .Y(n51971) );
  NAND2X1 U54620 ( .A(n51941), .B(n38001), .Y(n51970) );
  NOR2X1 U54621 ( .A(n51971), .B(n51970), .Y(n51939) );
  INVX1 U54622 ( .A(n28179), .Y(n73516) );
  NAND2X1 U54623 ( .A(n51939), .B(n73516), .Y(n54831) );
  INVX1 U54624 ( .A(n51970), .Y(n51969) );
  INVX1 U54625 ( .A(n28035), .Y(n73518) );
  NAND2X1 U54626 ( .A(n51969), .B(n73518), .Y(n55039) );
  NAND2X1 U54627 ( .A(n54831), .B(n55039), .Y(n56578) );
  NAND2X1 U54628 ( .A(n38001), .B(n28034), .Y(n51940) );
  NAND2X1 U54629 ( .A(n51941), .B(n51940), .Y(n51973) );
  NOR2X1 U54630 ( .A(n28032), .B(n28031), .Y(n51942) );
  OR2X1 U54631 ( .A(n26976), .B(n51942), .Y(n58246) );
  NAND2X1 U54632 ( .A(n51943), .B(n58246), .Y(n54405) );
  NAND2X1 U54633 ( .A(n43242), .B(n54405), .Y(n57241) );
  NAND2X1 U54634 ( .A(opcode_pc_w[1]), .B(n57241), .Y(n51946) );
  NAND2X1 U54635 ( .A(n27560), .B(n26331), .Y(n51944) );
  NAND2X1 U54636 ( .A(u_csr_csr_mepc_q[1]), .B(n51944), .Y(n51945) );
  NAND2X1 U54637 ( .A(n51946), .B(n51945), .Y(n51947) );
  NOR2X1 U54638 ( .A(n51948), .B(n51947), .Y(n51955) );
  NAND2X1 U54639 ( .A(n57427), .B(n73516), .Y(n58222) );
  NOR2X1 U54640 ( .A(n42952), .B(n37746), .Y(n51953) );
  INVX1 U54641 ( .A(n26014), .Y(n51949) );
  NAND2X1 U54642 ( .A(n51949), .B(n42442), .Y(n58343) );
  INVX1 U54643 ( .A(n58343), .Y(n73509) );
  INVX1 U54644 ( .A(n24943), .Y(n58243) );
  NAND2X1 U54645 ( .A(n38537), .B(n58243), .Y(n58202) );
  INVX1 U54646 ( .A(n58202), .Y(n57247) );
  NAND2X1 U54647 ( .A(n73509), .B(n57247), .Y(n51951) );
  NAND2X1 U54648 ( .A(n43286), .B(n56772), .Y(n51950) );
  NAND2X1 U54649 ( .A(n51951), .B(n51950), .Y(n51952) );
  NOR2X1 U54650 ( .A(n51953), .B(n51952), .Y(n51954) );
  NAND2X1 U54651 ( .A(n51955), .B(n51954), .Y(u_csr_csr_mepc_r[1]) );
  INVX1 U54652 ( .A(n24435), .Y(n51956) );
  NOR2X1 U54653 ( .A(n24440), .B(n51956), .Y(n51957) );
  NAND2X1 U54654 ( .A(n51957), .B(n24436), .Y(n51963) );
  NOR2X1 U54655 ( .A(n51959), .B(n51958), .Y(n51961) );
  NAND2X1 U54656 ( .A(n51961), .B(n51960), .Y(n51962) );
  NOR2X1 U54657 ( .A(n51963), .B(n51962), .Y(u_decode_N776) );
  NAND2X1 U54658 ( .A(n28520), .B(n51964), .Y(n26928) );
  NAND2X1 U54659 ( .A(n26928), .B(n26931), .Y(n26920) );
  INVX1 U54660 ( .A(n27325), .Y(n73576) );
  INVX1 U54661 ( .A(n28249), .Y(n73574) );
  NAND2X1 U54662 ( .A(n42215), .B(n73574), .Y(n26951) );
  INVX1 U54663 ( .A(n26920), .Y(n51966) );
  NAND2X1 U54664 ( .A(n26951), .B(n51966), .Y(n26252) );
  INVX1 U54665 ( .A(n26931), .Y(n73517) );
  NAND2X1 U54666 ( .A(n42308), .B(n43309), .Y(n57254) );
  NOR2X1 U54667 ( .A(n8836), .B(n57254), .Y(n51978) );
  OR2X1 U54668 ( .A(n51966), .B(n51965), .Y(n51968) );
  NAND2X1 U54669 ( .A(n43289), .B(n56773), .Y(n51976) );
  INVX1 U54670 ( .A(n26928), .Y(n73508) );
  NAND2X1 U54671 ( .A(n51969), .B(n73508), .Y(n55058) );
  NOR2X1 U54672 ( .A(n26931), .B(n51970), .Y(n51972) );
  INVX1 U54673 ( .A(n51971), .Y(n58128) );
  NAND2X1 U54674 ( .A(n51972), .B(n58128), .Y(n54850) );
  NAND2X1 U54675 ( .A(n55058), .B(n54850), .Y(n56590) );
  INVX1 U54676 ( .A(n26252), .Y(n73507) );
  NOR2X1 U54677 ( .A(n73507), .B(n57427), .Y(n51974) );
  NAND2X1 U54678 ( .A(n51974), .B(n51973), .Y(n54418) );
  NAND2X1 U54679 ( .A(n43252), .B(n54418), .Y(n57256) );
  NAND2X1 U54680 ( .A(opcode_pc_w[1]), .B(n57256), .Y(n51975) );
  NAND2X1 U54681 ( .A(n51976), .B(n51975), .Y(n51977) );
  NOR2X1 U54682 ( .A(n51978), .B(n51977), .Y(n51989) );
  INVX1 U54683 ( .A(n51979), .Y(n73365) );
  NAND2X1 U54684 ( .A(n73365), .B(opcode_opcode_w[26]), .Y(n51980) );
  NOR2X1 U54685 ( .A(n42748), .B(n51980), .Y(n51982) );
  NOR2X1 U54686 ( .A(opcode_opcode_w[29]), .B(opcode_opcode_w[27]), .Y(n51981)
         );
  NAND2X1 U54687 ( .A(n51982), .B(n51981), .Y(n58200) );
  INVX1 U54688 ( .A(n58200), .Y(n73506) );
  NAND2X1 U54689 ( .A(n73506), .B(n38537), .Y(n58274) );
  NOR2X1 U54690 ( .A(n58274), .B(n58343), .Y(n51985) );
  NAND2X1 U54691 ( .A(n57427), .B(n73517), .Y(n58251) );
  NOR2X1 U54692 ( .A(n42956), .B(n37746), .Y(n51984) );
  NOR2X1 U54693 ( .A(n51985), .B(n51984), .Y(n51987) );
  NAND2X1 U54694 ( .A(n26714), .B(u_csr_csr_sepc_q[1]), .Y(n51986) );
  AND2X1 U54695 ( .A(n51987), .B(n51986), .Y(n51988) );
  NAND2X1 U54696 ( .A(n51989), .B(n51988), .Y(u_csr_csr_sepc_r[1]) );
  AND2X1 U54697 ( .A(n28502), .B(n28500), .Y(n51995) );
  NOR2X1 U54698 ( .A(n73367), .B(n58211), .Y(n51990) );
  NOR2X1 U54699 ( .A(n58476), .B(n43292), .Y(n51993) );
  NAND2X1 U54700 ( .A(n28510), .B(opcode_instr_w_40), .Y(n51991) );
  NOR2X1 U54701 ( .A(n58475), .B(n43295), .Y(n51992) );
  NOR2X1 U54702 ( .A(n51993), .B(n51992), .Y(n51994) );
  NAND2X1 U54703 ( .A(n51995), .B(n51994), .Y(u_csr_N3666) );
  NAND2X1 U54704 ( .A(n43298), .B(n56773), .Y(n51997) );
  NAND2X1 U54705 ( .A(n43301), .B(n56772), .Y(n51996) );
  NAND2X1 U54706 ( .A(n51997), .B(n51996), .Y(net2282) );
  NAND2X1 U54707 ( .A(n43305), .B(n44863), .Y(n51999) );
  INVX1 U54708 ( .A(n51998), .Y(n57558) );
  NAND2X1 U54709 ( .A(n57558), .B(n44863), .Y(n54435) );
  NAND2X1 U54710 ( .A(challenge[100]), .B(n44855), .Y(n52000) );
  NAND2X1 U54711 ( .A(n42254), .B(n52000), .Y(n17308) );
  INVX1 U54712 ( .A(n52001), .Y(n58188) );
  NAND2X1 U54713 ( .A(n58188), .B(n57895), .Y(n55818) );
  INVX1 U54714 ( .A(n55818), .Y(n52007) );
  NAND2X1 U54715 ( .A(n57380), .B(n37550), .Y(n55816) );
  NOR2X1 U54716 ( .A(n58179), .B(n55816), .Y(n52006) );
  NAND2X1 U54717 ( .A(n52002), .B(n55307), .Y(n52004) );
  NAND2X1 U54718 ( .A(n58166), .B(n57895), .Y(n52003) );
  NAND2X1 U54719 ( .A(n52004), .B(n52003), .Y(n52005) );
  NAND2X1 U54720 ( .A(n52006), .B(n52005), .Y(n57397) );
  MX2X1 U54721 ( .A(u_mmu_dtlb_req_q), .B(n52007), .S0(n43380), .Y(n8554) );
  NAND2X1 U54722 ( .A(n42760), .B(n58817), .Y(n58213) );
  NOR2X1 U54723 ( .A(n58818), .B(n58816), .Y(n52009) );
  NOR2X1 U54724 ( .A(opcode_opcode_w[29]), .B(n38802), .Y(n52008) );
  NAND2X1 U54725 ( .A(n52009), .B(n52008), .Y(n57553) );
  OR2X1 U54726 ( .A(n27326), .B(n57553), .Y(n52010) );
  NOR2X1 U54727 ( .A(n58213), .B(n52010), .Y(n57385) );
  NOR2X1 U54728 ( .A(u_mmu_itlb_valid_q), .B(n37548), .Y(n52011) );
  NOR2X1 U54729 ( .A(n57385), .B(n52011), .Y(n8505) );
  NOR2X1 U54730 ( .A(n19678), .B(n43261), .Y(n52013) );
  NOR2X1 U54731 ( .A(n44535), .B(n43264), .Y(n52012) );
  NOR2X1 U54732 ( .A(n52013), .B(n52012), .Y(n52015) );
  NOR2X1 U54733 ( .A(n19843), .B(n19842), .Y(n52014) );
  NAND2X1 U54734 ( .A(n52015), .B(n52014), .Y(u_decode_u_regfile_N659) );
  NOR2X1 U54735 ( .A(n44601), .B(n43263), .Y(n52017) );
  NOR2X1 U54736 ( .A(n44598), .B(n37669), .Y(n52016) );
  NOR2X1 U54737 ( .A(n52017), .B(n52016), .Y(n52019) );
  NOR2X1 U54738 ( .A(n18271), .B(n18270), .Y(n52018) );
  NAND2X1 U54739 ( .A(n52019), .B(n52018), .Y(u_decode_u_regfile_N955) );
  NOR2X1 U54740 ( .A(n43261), .B(n43270), .Y(n52021) );
  NOR2X1 U54741 ( .A(n43264), .B(n43387), .Y(n52020) );
  NOR2X1 U54742 ( .A(n52021), .B(n52020), .Y(n52023) );
  NOR2X1 U54743 ( .A(n21413), .B(n21412), .Y(n52022) );
  NAND2X1 U54744 ( .A(n52023), .B(n52022), .Y(u_decode_u_regfile_N363) );
  NOR2X1 U54745 ( .A(n44472), .B(n43263), .Y(n52025) );
  NOR2X1 U54746 ( .A(n44469), .B(n37669), .Y(n52024) );
  NOR2X1 U54747 ( .A(n52025), .B(n52024), .Y(n52027) );
  NOR2X1 U54748 ( .A(n21020), .B(n21019), .Y(n52026) );
  NAND2X1 U54749 ( .A(n52027), .B(n52026), .Y(u_decode_u_regfile_N437) );
  NOR2X1 U54750 ( .A(n44559), .B(n43263), .Y(n52029) );
  NOR2X1 U54751 ( .A(n44556), .B(n37669), .Y(n52028) );
  NOR2X1 U54752 ( .A(n52029), .B(n52028), .Y(n52031) );
  NOR2X1 U54753 ( .A(n19448), .B(n19447), .Y(n52030) );
  NAND2X1 U54754 ( .A(n52031), .B(n52030), .Y(u_decode_u_regfile_N733) );
  NOR2X1 U54755 ( .A(n44382), .B(n43263), .Y(n52033) );
  NOR2X1 U54756 ( .A(n44379), .B(n43265), .Y(n52032) );
  NOR2X1 U54757 ( .A(n52033), .B(n52032), .Y(n52035) );
  NOR2X1 U54758 ( .A(n22590), .B(n22589), .Y(n52034) );
  NAND2X1 U54759 ( .A(n52035), .B(n52034), .Y(u_decode_u_regfile_N141) );
  NOR2X1 U54760 ( .A(n44304), .B(n43262), .Y(n52037) );
  NOR2X1 U54761 ( .A(n44301), .B(n43265), .Y(n52036) );
  NOR2X1 U54762 ( .A(n52037), .B(n52036), .Y(n52039) );
  NOR2X1 U54763 ( .A(n23944), .B(n23943), .Y(n52038) );
  NAND2X1 U54764 ( .A(n52039), .B(n52038), .Y(u_decode_u_regfile_N1029) );
  NOR2X1 U54765 ( .A(n44571), .B(n43262), .Y(n52041) );
  NOR2X1 U54766 ( .A(n44568), .B(n43265), .Y(n52040) );
  NOR2X1 U54767 ( .A(n52041), .B(n52040), .Y(n52043) );
  NOR2X1 U54768 ( .A(n19056), .B(n19055), .Y(n52042) );
  NAND2X1 U54769 ( .A(n52043), .B(n52042), .Y(u_decode_u_regfile_N807) );
  NOR2X1 U54770 ( .A(n43261), .B(n43276), .Y(n52045) );
  NOR2X1 U54771 ( .A(n43264), .B(n43384), .Y(n52044) );
  NOR2X1 U54772 ( .A(n52045), .B(n52044), .Y(n52047) );
  NOR2X1 U54773 ( .A(n20628), .B(n20627), .Y(n52046) );
  NAND2X1 U54774 ( .A(n52047), .B(n52046), .Y(u_decode_u_regfile_N511) );
  NOR2X1 U54775 ( .A(n44406), .B(n43262), .Y(n52049) );
  NOR2X1 U54776 ( .A(n44403), .B(n43265), .Y(n52048) );
  NOR2X1 U54777 ( .A(n52049), .B(n52048), .Y(n52051) );
  NOR2X1 U54778 ( .A(n22198), .B(n22197), .Y(n52050) );
  NAND2X1 U54779 ( .A(n52051), .B(n52050), .Y(u_decode_u_regfile_N215) );
  NOR2X1 U54780 ( .A(n44328), .B(n43262), .Y(n52053) );
  NOR2X1 U54781 ( .A(n44325), .B(n43265), .Y(n52052) );
  NOR2X1 U54782 ( .A(n52053), .B(n52052), .Y(n52055) );
  NOR2X1 U54783 ( .A(n23504), .B(n23503), .Y(n52054) );
  NAND2X1 U54784 ( .A(n52055), .B(n52054), .Y(u_decode_u_regfile_N1103) );
  NOR2X1 U54785 ( .A(n44583), .B(n43262), .Y(n52057) );
  NOR2X1 U54786 ( .A(n44580), .B(n43265), .Y(n52056) );
  NOR2X1 U54787 ( .A(n52057), .B(n52056), .Y(n52059) );
  NOR2X1 U54788 ( .A(n18664), .B(n18663), .Y(n52058) );
  NAND2X1 U54789 ( .A(n52059), .B(n52058), .Y(u_decode_u_regfile_N881) );
  NOR2X1 U54790 ( .A(n44430), .B(n43262), .Y(n52061) );
  NOR2X1 U54791 ( .A(n44427), .B(n43265), .Y(n52060) );
  NOR2X1 U54792 ( .A(n52061), .B(n52060), .Y(n52063) );
  NOR2X1 U54793 ( .A(n21806), .B(n21805), .Y(n52062) );
  NAND2X1 U54794 ( .A(n52063), .B(n52062), .Y(u_decode_u_regfile_N289) );
  NOR2X1 U54795 ( .A(n44514), .B(n43262), .Y(n52065) );
  NOR2X1 U54796 ( .A(n44511), .B(n43265), .Y(n52064) );
  NOR2X1 U54797 ( .A(n52065), .B(n52064), .Y(n52067) );
  NOR2X1 U54798 ( .A(n20236), .B(n20235), .Y(n52066) );
  NAND2X1 U54799 ( .A(n52067), .B(n52066), .Y(u_decode_u_regfile_N585) );
  NOR2X1 U54800 ( .A(n44352), .B(n43262), .Y(n52069) );
  NOR2X1 U54801 ( .A(n44349), .B(n43265), .Y(n52068) );
  NOR2X1 U54802 ( .A(n52069), .B(n52068), .Y(n52071) );
  NOR2X1 U54803 ( .A(n23070), .B(n23069), .Y(n52070) );
  NAND2X1 U54804 ( .A(n52071), .B(n52070), .Y(u_decode_u_regfile_N1177) );
  NOR2X1 U54805 ( .A(n44607), .B(n43262), .Y(n52073) );
  NOR2X1 U54806 ( .A(n44604), .B(n43265), .Y(n52072) );
  NOR2X1 U54807 ( .A(n52073), .B(n52072), .Y(n52075) );
  NOR2X1 U54808 ( .A(n18053), .B(n18051), .Y(n52074) );
  NAND2X1 U54809 ( .A(n52075), .B(n52074), .Y(u_decode_u_regfile_N992) );
  NOR2X1 U54810 ( .A(n43261), .B(n43273), .Y(n52077) );
  NOR2X1 U54811 ( .A(n43264), .B(n43390), .Y(n52076) );
  NOR2X1 U54812 ( .A(n52077), .B(n52076), .Y(n52079) );
  NOR2X1 U54813 ( .A(n23872), .B(n23871), .Y(n52078) );
  NAND2X1 U54814 ( .A(n52079), .B(n52078), .Y(u_decode_u_regfile_N104) );
  NOR2X1 U54815 ( .A(n44460), .B(n43262), .Y(n52081) );
  NOR2X1 U54816 ( .A(n44457), .B(n43265), .Y(n52080) );
  NOR2X1 U54817 ( .A(n52081), .B(n52080), .Y(n52083) );
  NOR2X1 U54818 ( .A(n21216), .B(n21215), .Y(n52082) );
  NAND2X1 U54819 ( .A(n52083), .B(n52082), .Y(u_decode_u_regfile_N400) );
  NOR2X1 U54820 ( .A(n44550), .B(n43262), .Y(n52085) );
  NOR2X1 U54821 ( .A(n44547), .B(n43265), .Y(n52084) );
  NOR2X1 U54822 ( .A(n52085), .B(n52084), .Y(n52087) );
  NOR2X1 U54823 ( .A(n19646), .B(n19645), .Y(n52086) );
  NAND2X1 U54824 ( .A(n52087), .B(n52086), .Y(u_decode_u_regfile_N696) );
  NOR2X1 U54825 ( .A(n44565), .B(n43262), .Y(n52089) );
  NOR2X1 U54826 ( .A(n44562), .B(n43264), .Y(n52088) );
  NOR2X1 U54827 ( .A(n52089), .B(n52088), .Y(n52091) );
  NOR2X1 U54828 ( .A(n19252), .B(n19251), .Y(n52090) );
  NAND2X1 U54829 ( .A(n52091), .B(n52090), .Y(u_decode_u_regfile_N770) );
  NOR2X1 U54830 ( .A(n44316), .B(n43261), .Y(n52093) );
  NOR2X1 U54831 ( .A(n44313), .B(n43264), .Y(n52092) );
  NOR2X1 U54832 ( .A(n52093), .B(n52092), .Y(n52095) );
  NOR2X1 U54833 ( .A(n23724), .B(n23723), .Y(n52094) );
  NAND2X1 U54834 ( .A(n52095), .B(n52094), .Y(u_decode_u_regfile_N1066) );
  NOR2X1 U54835 ( .A(n44394), .B(n43261), .Y(n52097) );
  NOR2X1 U54836 ( .A(n44391), .B(n43264), .Y(n52096) );
  NOR2X1 U54837 ( .A(n52097), .B(n52096), .Y(n52099) );
  NOR2X1 U54838 ( .A(n22394), .B(n22393), .Y(n52098) );
  NAND2X1 U54839 ( .A(n52099), .B(n52098), .Y(u_decode_u_regfile_N178) );
  NOR2X1 U54840 ( .A(n44484), .B(n43261), .Y(n52101) );
  NOR2X1 U54841 ( .A(n44481), .B(n43264), .Y(n52100) );
  NOR2X1 U54842 ( .A(n52101), .B(n52100), .Y(n52103) );
  NOR2X1 U54843 ( .A(n20824), .B(n20823), .Y(n52102) );
  NAND2X1 U54844 ( .A(n52103), .B(n52102), .Y(u_decode_u_regfile_N474) );
  NOR2X1 U54845 ( .A(n44418), .B(n43262), .Y(n52105) );
  NOR2X1 U54846 ( .A(n44415), .B(n43265), .Y(n52104) );
  NOR2X1 U54847 ( .A(n52105), .B(n52104), .Y(n52107) );
  NOR2X1 U54848 ( .A(n22002), .B(n22001), .Y(n52106) );
  NAND2X1 U54849 ( .A(n52107), .B(n52106), .Y(u_decode_u_regfile_N252) );
  NOR2X1 U54850 ( .A(n44340), .B(n43261), .Y(n52109) );
  NOR2X1 U54851 ( .A(n44337), .B(n43264), .Y(n52108) );
  NOR2X1 U54852 ( .A(n52109), .B(n52108), .Y(n52111) );
  NOR2X1 U54853 ( .A(n23284), .B(n23283), .Y(n52110) );
  NAND2X1 U54854 ( .A(n52111), .B(n52110), .Y(u_decode_u_regfile_N1140) );
  NOR2X1 U54855 ( .A(n44502), .B(n43261), .Y(n52113) );
  NOR2X1 U54856 ( .A(n44499), .B(n43264), .Y(n52112) );
  NOR2X1 U54857 ( .A(n52113), .B(n52112), .Y(n52115) );
  NOR2X1 U54858 ( .A(n20432), .B(n20431), .Y(n52114) );
  NAND2X1 U54859 ( .A(n52115), .B(n52114), .Y(u_decode_u_regfile_N548) );
  NOR2X1 U54860 ( .A(n44577), .B(n43261), .Y(n52117) );
  NOR2X1 U54861 ( .A(n44574), .B(n43264), .Y(n52116) );
  NOR2X1 U54862 ( .A(n52117), .B(n52116), .Y(n52119) );
  NOR2X1 U54863 ( .A(n18860), .B(n18859), .Y(n52118) );
  NAND2X1 U54864 ( .A(n52119), .B(n52118), .Y(u_decode_u_regfile_N844) );
  NOR2X1 U54865 ( .A(n44526), .B(n43261), .Y(n52121) );
  NOR2X1 U54866 ( .A(n44523), .B(n43264), .Y(n52120) );
  NOR2X1 U54867 ( .A(n52121), .B(n52120), .Y(n52123) );
  NOR2X1 U54868 ( .A(n20040), .B(n20039), .Y(n52122) );
  NAND2X1 U54869 ( .A(n52123), .B(n52122), .Y(u_decode_u_regfile_N622) );
  NOR2X1 U54870 ( .A(n44592), .B(n43261), .Y(n52125) );
  NOR2X1 U54871 ( .A(n44589), .B(n43264), .Y(n52124) );
  NOR2X1 U54872 ( .A(n52125), .B(n52124), .Y(n52127) );
  NOR2X1 U54873 ( .A(n18470), .B(n18469), .Y(n52126) );
  NAND2X1 U54874 ( .A(n52127), .B(n52126), .Y(u_decode_u_regfile_N918) );
  NOR2X1 U54875 ( .A(n44442), .B(n43261), .Y(n52129) );
  NOR2X1 U54876 ( .A(n44439), .B(n43264), .Y(n52128) );
  NOR2X1 U54877 ( .A(n52129), .B(n52128), .Y(n52131) );
  NOR2X1 U54878 ( .A(n21610), .B(n21609), .Y(n52130) );
  NAND2X1 U54879 ( .A(n52131), .B(n52130), .Y(u_decode_u_regfile_N326) );
  NOR2X1 U54880 ( .A(n44460), .B(n43329), .Y(n52133) );
  NOR2X1 U54881 ( .A(n44457), .B(n43332), .Y(n52132) );
  NOR2X1 U54882 ( .A(n52133), .B(n52132), .Y(n52135) );
  NOR2X1 U54883 ( .A(n21228), .B(n21227), .Y(n52134) );
  NAND2X1 U54884 ( .A(n52135), .B(n52134), .Y(u_decode_u_regfile_N398) );
  NOR2X1 U54885 ( .A(n44352), .B(n43331), .Y(n52137) );
  NOR2X1 U54886 ( .A(n44349), .B(n37687), .Y(n52136) );
  NOR2X1 U54887 ( .A(n52137), .B(n52136), .Y(n52139) );
  NOR2X1 U54888 ( .A(n23082), .B(n23081), .Y(n52138) );
  NAND2X1 U54889 ( .A(n52139), .B(n52138), .Y(u_decode_u_regfile_N1175) );
  NOR2X1 U54890 ( .A(n44340), .B(n43331), .Y(n52141) );
  NOR2X1 U54891 ( .A(n44337), .B(n37687), .Y(n52140) );
  NOR2X1 U54892 ( .A(n52141), .B(n52140), .Y(n52143) );
  NOR2X1 U54893 ( .A(n23302), .B(n23301), .Y(n52142) );
  NAND2X1 U54894 ( .A(n52143), .B(n52142), .Y(u_decode_u_regfile_N1138) );
  NOR2X1 U54895 ( .A(n44592), .B(n43331), .Y(n52145) );
  NOR2X1 U54896 ( .A(n44589), .B(n37687), .Y(n52144) );
  NOR2X1 U54897 ( .A(n52145), .B(n52144), .Y(n52147) );
  NOR2X1 U54898 ( .A(n18482), .B(n18481), .Y(n52146) );
  NAND2X1 U54899 ( .A(n52147), .B(n52146), .Y(u_decode_u_regfile_N916) );
  NOR2X1 U54900 ( .A(n44577), .B(n43331), .Y(n52149) );
  NOR2X1 U54901 ( .A(n44574), .B(n43333), .Y(n52148) );
  NOR2X1 U54902 ( .A(n52149), .B(n52148), .Y(n52151) );
  NOR2X1 U54903 ( .A(n18872), .B(n18871), .Y(n52150) );
  NAND2X1 U54904 ( .A(n52151), .B(n52150), .Y(u_decode_u_regfile_N842) );
  NOR2X1 U54905 ( .A(n44565), .B(n43331), .Y(n52153) );
  NOR2X1 U54906 ( .A(n44562), .B(n43333), .Y(n52152) );
  NOR2X1 U54907 ( .A(n52153), .B(n52152), .Y(n52155) );
  NOR2X1 U54908 ( .A(n19264), .B(n19263), .Y(n52154) );
  NAND2X1 U54909 ( .A(n52155), .B(n52154), .Y(u_decode_u_regfile_N768) );
  NOR2X1 U54910 ( .A(n44559), .B(n43331), .Y(n52157) );
  NOR2X1 U54911 ( .A(n44556), .B(n43333), .Y(n52156) );
  NOR2X1 U54912 ( .A(n52157), .B(n52156), .Y(n52159) );
  NOR2X1 U54913 ( .A(n19460), .B(n19459), .Y(n52158) );
  NAND2X1 U54914 ( .A(n52159), .B(n52158), .Y(u_decode_u_regfile_N731) );
  NOR2X1 U54915 ( .A(n44571), .B(n43330), .Y(n52161) );
  NOR2X1 U54916 ( .A(n44568), .B(n43333), .Y(n52160) );
  NOR2X1 U54917 ( .A(n52161), .B(n52160), .Y(n52163) );
  NOR2X1 U54918 ( .A(n19068), .B(n19067), .Y(n52162) );
  NAND2X1 U54919 ( .A(n52163), .B(n52162), .Y(u_decode_u_regfile_N805) );
  NOR2X1 U54920 ( .A(n44442), .B(n43330), .Y(n52165) );
  NOR2X1 U54921 ( .A(n44439), .B(n43333), .Y(n52164) );
  NOR2X1 U54922 ( .A(n52165), .B(n52164), .Y(n52167) );
  NOR2X1 U54923 ( .A(n21622), .B(n21621), .Y(n52166) );
  NAND2X1 U54924 ( .A(n52167), .B(n52166), .Y(u_decode_u_regfile_N324) );
  NOR2X1 U54925 ( .A(n44406), .B(n43330), .Y(n52169) );
  NOR2X1 U54926 ( .A(n44403), .B(n43333), .Y(n52168) );
  NOR2X1 U54927 ( .A(n52169), .B(n52168), .Y(n52171) );
  NOR2X1 U54928 ( .A(n22210), .B(n22209), .Y(n52170) );
  NAND2X1 U54929 ( .A(n52171), .B(n52170), .Y(u_decode_u_regfile_N213) );
  NOR2X1 U54930 ( .A(n44382), .B(n43330), .Y(n52173) );
  NOR2X1 U54931 ( .A(n44379), .B(n43333), .Y(n52172) );
  NOR2X1 U54932 ( .A(n52173), .B(n52172), .Y(n52175) );
  NOR2X1 U54933 ( .A(n22602), .B(n22601), .Y(n52174) );
  NAND2X1 U54934 ( .A(n52175), .B(n52174), .Y(u_decode_u_regfile_N139) );
  NOR2X1 U54935 ( .A(n44418), .B(n43330), .Y(n52177) );
  NOR2X1 U54936 ( .A(n44415), .B(n43333), .Y(n52176) );
  NOR2X1 U54937 ( .A(n52177), .B(n52176), .Y(n52179) );
  NOR2X1 U54938 ( .A(n22014), .B(n22013), .Y(n52178) );
  NAND2X1 U54939 ( .A(n52179), .B(n52178), .Y(u_decode_u_regfile_N250) );
  NOR2X1 U54940 ( .A(n44394), .B(n43330), .Y(n52181) );
  NOR2X1 U54941 ( .A(n44391), .B(n43333), .Y(n52180) );
  NOR2X1 U54942 ( .A(n52181), .B(n52180), .Y(n52183) );
  NOR2X1 U54943 ( .A(n22406), .B(n22405), .Y(n52182) );
  NAND2X1 U54944 ( .A(n52183), .B(n52182), .Y(u_decode_u_regfile_N176) );
  NOR2X1 U54945 ( .A(n44583), .B(n43330), .Y(n52185) );
  NOR2X1 U54946 ( .A(n44580), .B(n43333), .Y(n52184) );
  NOR2X1 U54947 ( .A(n52185), .B(n52184), .Y(n52187) );
  NOR2X1 U54948 ( .A(n18676), .B(n18675), .Y(n52186) );
  NAND2X1 U54949 ( .A(n52187), .B(n52186), .Y(u_decode_u_regfile_N879) );
  NOR2X1 U54950 ( .A(n44430), .B(n43330), .Y(n52189) );
  NOR2X1 U54951 ( .A(n44427), .B(n43333), .Y(n52188) );
  NOR2X1 U54952 ( .A(n52189), .B(n52188), .Y(n52191) );
  NOR2X1 U54953 ( .A(n21818), .B(n21817), .Y(n52190) );
  NAND2X1 U54954 ( .A(n52191), .B(n52190), .Y(u_decode_u_regfile_N287) );
  NOR2X1 U54955 ( .A(n43329), .B(n43273), .Y(n52193) );
  NOR2X1 U54956 ( .A(n43332), .B(n43390), .Y(n52192) );
  NOR2X1 U54957 ( .A(n52193), .B(n52192), .Y(n52195) );
  NOR2X1 U54958 ( .A(n23974), .B(n23973), .Y(n52194) );
  NAND2X1 U54959 ( .A(n52195), .B(n52194), .Y(u_decode_u_regfile_N102) );
  NOR2X1 U54960 ( .A(n44550), .B(n43330), .Y(n52197) );
  NOR2X1 U54961 ( .A(n44547), .B(n43333), .Y(n52196) );
  NOR2X1 U54962 ( .A(n52197), .B(n52196), .Y(n52199) );
  NOR2X1 U54963 ( .A(n19658), .B(n19657), .Y(n52198) );
  NAND2X1 U54964 ( .A(n52199), .B(n52198), .Y(u_decode_u_regfile_N694) );
  NOR2X1 U54965 ( .A(n43329), .B(n43270), .Y(n52201) );
  NOR2X1 U54966 ( .A(n43332), .B(n43387), .Y(n52200) );
  NOR2X1 U54967 ( .A(n52201), .B(n52200), .Y(n52203) );
  NOR2X1 U54968 ( .A(n21425), .B(n21424), .Y(n52202) );
  NAND2X1 U54969 ( .A(n52203), .B(n52202), .Y(u_decode_u_regfile_N361) );
  NOR2X1 U54970 ( .A(n44502), .B(n43330), .Y(n52205) );
  NOR2X1 U54971 ( .A(n44499), .B(n43332), .Y(n52204) );
  NOR2X1 U54972 ( .A(n52205), .B(n52204), .Y(n52207) );
  NOR2X1 U54973 ( .A(n20444), .B(n20443), .Y(n52206) );
  NAND2X1 U54974 ( .A(n52207), .B(n52206), .Y(u_decode_u_regfile_N546) );
  NOR2X1 U54975 ( .A(n43329), .B(n43276), .Y(n52209) );
  NOR2X1 U54976 ( .A(n43332), .B(n43384), .Y(n52208) );
  NOR2X1 U54977 ( .A(n52209), .B(n52208), .Y(n52211) );
  NOR2X1 U54978 ( .A(n20640), .B(n20639), .Y(n52210) );
  NAND2X1 U54979 ( .A(n52211), .B(n52210), .Y(u_decode_u_regfile_N509) );
  NOR2X1 U54980 ( .A(n44472), .B(n43330), .Y(n52213) );
  NOR2X1 U54981 ( .A(n44469), .B(n43332), .Y(n52212) );
  NOR2X1 U54982 ( .A(n52213), .B(n52212), .Y(n52215) );
  NOR2X1 U54983 ( .A(n21032), .B(n21031), .Y(n52214) );
  NAND2X1 U54984 ( .A(n52215), .B(n52214), .Y(u_decode_u_regfile_N435) );
  NOR2X1 U54985 ( .A(n44514), .B(n43330), .Y(n52217) );
  NOR2X1 U54986 ( .A(n44511), .B(n43333), .Y(n52216) );
  NOR2X1 U54987 ( .A(n52217), .B(n52216), .Y(n52219) );
  NOR2X1 U54988 ( .A(n20248), .B(n20247), .Y(n52218) );
  NAND2X1 U54989 ( .A(n52219), .B(n52218), .Y(u_decode_u_regfile_N583) );
  NOR2X1 U54990 ( .A(n44526), .B(n43330), .Y(n52221) );
  NOR2X1 U54991 ( .A(n44523), .B(n43332), .Y(n52220) );
  NOR2X1 U54992 ( .A(n52221), .B(n52220), .Y(n52223) );
  NOR2X1 U54993 ( .A(n20052), .B(n20051), .Y(n52222) );
  NAND2X1 U54994 ( .A(n52223), .B(n52222), .Y(u_decode_u_regfile_N620) );
  NOR2X1 U54995 ( .A(n44484), .B(n43329), .Y(n52225) );
  NOR2X1 U54996 ( .A(n44481), .B(n43332), .Y(n52224) );
  NOR2X1 U54997 ( .A(n52225), .B(n52224), .Y(n52227) );
  NOR2X1 U54998 ( .A(n20836), .B(n20835), .Y(n52226) );
  NAND2X1 U54999 ( .A(n52227), .B(n52226), .Y(u_decode_u_regfile_N472) );
  NOR2X1 U55000 ( .A(n44601), .B(n43329), .Y(n52229) );
  NOR2X1 U55001 ( .A(n44598), .B(n43332), .Y(n52228) );
  NOR2X1 U55002 ( .A(n52229), .B(n52228), .Y(n52231) );
  NOR2X1 U55003 ( .A(n18283), .B(n18282), .Y(n52230) );
  NAND2X1 U55004 ( .A(n52231), .B(n52230), .Y(u_decode_u_regfile_N953) );
  NOR2X1 U55005 ( .A(n44316), .B(n43329), .Y(n52233) );
  NOR2X1 U55006 ( .A(n44313), .B(n43332), .Y(n52232) );
  NOR2X1 U55007 ( .A(n52233), .B(n52232), .Y(n52235) );
  NOR2X1 U55008 ( .A(n23736), .B(n23735), .Y(n52234) );
  NAND2X1 U55009 ( .A(n52235), .B(n52234), .Y(u_decode_u_regfile_N1064) );
  NOR2X1 U55010 ( .A(n44328), .B(n43329), .Y(n52237) );
  NOR2X1 U55011 ( .A(n44325), .B(n43332), .Y(n52236) );
  NOR2X1 U55012 ( .A(n52237), .B(n52236), .Y(n52239) );
  NOR2X1 U55013 ( .A(n23516), .B(n23515), .Y(n52238) );
  NAND2X1 U55014 ( .A(n52239), .B(n52238), .Y(u_decode_u_regfile_N1101) );
  NOR2X1 U55015 ( .A(n44304), .B(n43329), .Y(n52241) );
  NOR2X1 U55016 ( .A(n44301), .B(n43332), .Y(n52240) );
  NOR2X1 U55017 ( .A(n52241), .B(n52240), .Y(n52243) );
  NOR2X1 U55018 ( .A(n23956), .B(n23955), .Y(n52242) );
  NAND2X1 U55019 ( .A(n52243), .B(n52242), .Y(u_decode_u_regfile_N1027) );
  NOR2X1 U55020 ( .A(n44607), .B(n43329), .Y(n52245) );
  NOR2X1 U55021 ( .A(n44604), .B(n43332), .Y(n52244) );
  NOR2X1 U55022 ( .A(n52245), .B(n52244), .Y(n52247) );
  NOR2X1 U55023 ( .A(n18067), .B(n18065), .Y(n52246) );
  NAND2X1 U55024 ( .A(n52247), .B(n52246), .Y(u_decode_u_regfile_N990) );
  NOR2X1 U55025 ( .A(n19678), .B(n43329), .Y(n52249) );
  NOR2X1 U55026 ( .A(n44535), .B(n43332), .Y(n52248) );
  NOR2X1 U55027 ( .A(n52249), .B(n52248), .Y(n52251) );
  NOR2X1 U55028 ( .A(n19855), .B(n19854), .Y(n52250) );
  NAND2X1 U55029 ( .A(n52251), .B(n52250), .Y(u_decode_u_regfile_N657) );
  NOR2X1 U55030 ( .A(n15400), .B(n15401), .Y(n52253) );
  NOR2X1 U55031 ( .A(n15436), .B(n15437), .Y(n52252) );
  NAND2X1 U55032 ( .A(n52253), .B(n52252), .Y(u_exec_alu_p_w[9]) );
  NOR2X1 U55033 ( .A(n44539), .B(n43121), .Y(n52255) );
  NOR2X1 U55034 ( .A(n44535), .B(n37674), .Y(n52254) );
  NOR2X1 U55035 ( .A(n52255), .B(n52254), .Y(n52257) );
  NOR2X1 U55036 ( .A(n19813), .B(n19812), .Y(n52256) );
  NAND2X1 U55037 ( .A(n52257), .B(n52256), .Y(u_decode_u_regfile_N664) );
  NOR2X1 U55038 ( .A(n44601), .B(n43122), .Y(n52259) );
  NOR2X1 U55039 ( .A(n44598), .B(n37674), .Y(n52258) );
  NOR2X1 U55040 ( .A(n52259), .B(n52258), .Y(n52261) );
  NOR2X1 U55041 ( .A(n18241), .B(n18240), .Y(n52260) );
  NAND2X1 U55042 ( .A(n52261), .B(n52260), .Y(u_decode_u_regfile_N960) );
  NOR2X1 U55043 ( .A(n43120), .B(n43270), .Y(n52263) );
  NOR2X1 U55044 ( .A(n43123), .B(n43387), .Y(n52262) );
  NOR2X1 U55045 ( .A(n52263), .B(n52262), .Y(n52265) );
  NOR2X1 U55046 ( .A(n21383), .B(n21382), .Y(n52264) );
  NAND2X1 U55047 ( .A(n52265), .B(n52264), .Y(u_decode_u_regfile_N368) );
  NOR2X1 U55048 ( .A(n44472), .B(n43122), .Y(n52267) );
  NOR2X1 U55049 ( .A(n44469), .B(n37674), .Y(n52266) );
  NOR2X1 U55050 ( .A(n52267), .B(n52266), .Y(n52269) );
  NOR2X1 U55051 ( .A(n20990), .B(n20989), .Y(n52268) );
  NAND2X1 U55052 ( .A(n52269), .B(n52268), .Y(u_decode_u_regfile_N442) );
  NOR2X1 U55053 ( .A(n44559), .B(n43122), .Y(n52271) );
  NOR2X1 U55054 ( .A(n44556), .B(n37674), .Y(n52270) );
  NOR2X1 U55055 ( .A(n52271), .B(n52270), .Y(n52273) );
  NOR2X1 U55056 ( .A(n19418), .B(n19417), .Y(n52272) );
  NAND2X1 U55057 ( .A(n52273), .B(n52272), .Y(u_decode_u_regfile_N738) );
  NOR2X1 U55058 ( .A(n44382), .B(n43122), .Y(n52275) );
  NOR2X1 U55059 ( .A(n44379), .B(n43124), .Y(n52274) );
  NOR2X1 U55060 ( .A(n52275), .B(n52274), .Y(n52277) );
  NOR2X1 U55061 ( .A(n22560), .B(n22559), .Y(n52276) );
  NAND2X1 U55062 ( .A(n52277), .B(n52276), .Y(u_decode_u_regfile_N146) );
  NOR2X1 U55063 ( .A(n44304), .B(n43122), .Y(n52279) );
  NOR2X1 U55064 ( .A(n44301), .B(n43124), .Y(n52278) );
  NOR2X1 U55065 ( .A(n52279), .B(n52278), .Y(n52281) );
  NOR2X1 U55066 ( .A(n23908), .B(n23907), .Y(n52280) );
  NAND2X1 U55067 ( .A(n52281), .B(n52280), .Y(u_decode_u_regfile_N1034) );
  NOR2X1 U55068 ( .A(n44571), .B(n43122), .Y(n52283) );
  NOR2X1 U55069 ( .A(n44568), .B(n43124), .Y(n52282) );
  NOR2X1 U55070 ( .A(n52283), .B(n52282), .Y(n52285) );
  NOR2X1 U55071 ( .A(n19026), .B(n19025), .Y(n52284) );
  NAND2X1 U55072 ( .A(n52285), .B(n52284), .Y(u_decode_u_regfile_N812) );
  NOR2X1 U55073 ( .A(n43120), .B(n43276), .Y(n52287) );
  NOR2X1 U55074 ( .A(n43123), .B(n43384), .Y(n52286) );
  NOR2X1 U55075 ( .A(n52287), .B(n52286), .Y(n52289) );
  NOR2X1 U55076 ( .A(n20598), .B(n20597), .Y(n52288) );
  NAND2X1 U55077 ( .A(n52289), .B(n52288), .Y(u_decode_u_regfile_N516) );
  NOR2X1 U55078 ( .A(n44406), .B(n43121), .Y(n52291) );
  NOR2X1 U55079 ( .A(n44403), .B(n43124), .Y(n52290) );
  NOR2X1 U55080 ( .A(n52291), .B(n52290), .Y(n52293) );
  NOR2X1 U55081 ( .A(n22168), .B(n22167), .Y(n52292) );
  NAND2X1 U55082 ( .A(n52293), .B(n52292), .Y(u_decode_u_regfile_N220) );
  NOR2X1 U55083 ( .A(n44328), .B(n43121), .Y(n52295) );
  NOR2X1 U55084 ( .A(n44325), .B(n43124), .Y(n52294) );
  NOR2X1 U55085 ( .A(n52295), .B(n52294), .Y(n52297) );
  NOR2X1 U55086 ( .A(n23474), .B(n23473), .Y(n52296) );
  NAND2X1 U55087 ( .A(n52297), .B(n52296), .Y(u_decode_u_regfile_N1108) );
  NOR2X1 U55088 ( .A(n44583), .B(n43121), .Y(n52299) );
  NOR2X1 U55089 ( .A(n44580), .B(n43124), .Y(n52298) );
  NOR2X1 U55090 ( .A(n52299), .B(n52298), .Y(n52301) );
  NOR2X1 U55091 ( .A(n18634), .B(n18633), .Y(n52300) );
  NAND2X1 U55092 ( .A(n52301), .B(n52300), .Y(u_decode_u_regfile_N886) );
  NOR2X1 U55093 ( .A(n44430), .B(n43121), .Y(n52303) );
  NOR2X1 U55094 ( .A(n44427), .B(n43124), .Y(n52302) );
  NOR2X1 U55095 ( .A(n52303), .B(n52302), .Y(n52305) );
  NOR2X1 U55096 ( .A(n21776), .B(n21775), .Y(n52304) );
  NAND2X1 U55097 ( .A(n52305), .B(n52304), .Y(u_decode_u_regfile_N294) );
  NOR2X1 U55098 ( .A(n44514), .B(n43121), .Y(n52307) );
  NOR2X1 U55099 ( .A(n44511), .B(n43124), .Y(n52306) );
  NOR2X1 U55100 ( .A(n52307), .B(n52306), .Y(n52309) );
  NOR2X1 U55101 ( .A(n20206), .B(n20205), .Y(n52308) );
  NAND2X1 U55102 ( .A(n52309), .B(n52308), .Y(u_decode_u_regfile_N590) );
  NOR2X1 U55103 ( .A(n44352), .B(n43121), .Y(n52311) );
  NOR2X1 U55104 ( .A(n44349), .B(n43124), .Y(n52310) );
  NOR2X1 U55105 ( .A(n52311), .B(n52310), .Y(n52313) );
  NOR2X1 U55106 ( .A(n23034), .B(n23033), .Y(n52312) );
  NAND2X1 U55107 ( .A(n52313), .B(n52312), .Y(u_decode_u_regfile_N1182) );
  NOR2X1 U55108 ( .A(n44607), .B(n43121), .Y(n52315) );
  NOR2X1 U55109 ( .A(n44604), .B(n43124), .Y(n52314) );
  NOR2X1 U55110 ( .A(n52315), .B(n52314), .Y(n52317) );
  NOR2X1 U55111 ( .A(n18018), .B(n18016), .Y(n52316) );
  NAND2X1 U55112 ( .A(n52317), .B(n52316), .Y(u_decode_u_regfile_N997) );
  NOR2X1 U55113 ( .A(n43120), .B(n43273), .Y(n52319) );
  NOR2X1 U55114 ( .A(n43123), .B(n43390), .Y(n52318) );
  NOR2X1 U55115 ( .A(n52319), .B(n52318), .Y(n52321) );
  NOR2X1 U55116 ( .A(n23568), .B(n23567), .Y(n52320) );
  NAND2X1 U55117 ( .A(n52321), .B(n52320), .Y(u_decode_u_regfile_N109) );
  NOR2X1 U55118 ( .A(n44460), .B(n43121), .Y(n52323) );
  NOR2X1 U55119 ( .A(n44457), .B(n43124), .Y(n52322) );
  NOR2X1 U55120 ( .A(n52323), .B(n52322), .Y(n52325) );
  NOR2X1 U55121 ( .A(n21186), .B(n21185), .Y(n52324) );
  NAND2X1 U55122 ( .A(n52325), .B(n52324), .Y(u_decode_u_regfile_N405) );
  NOR2X1 U55123 ( .A(n44550), .B(n43121), .Y(n52327) );
  NOR2X1 U55124 ( .A(n44547), .B(n43124), .Y(n52326) );
  NOR2X1 U55125 ( .A(n52327), .B(n52326), .Y(n52329) );
  NOR2X1 U55126 ( .A(n19616), .B(n19615), .Y(n52328) );
  NAND2X1 U55127 ( .A(n52329), .B(n52328), .Y(u_decode_u_regfile_N701) );
  NOR2X1 U55128 ( .A(n44565), .B(n43121), .Y(n52331) );
  NOR2X1 U55129 ( .A(n44562), .B(n43123), .Y(n52330) );
  NOR2X1 U55130 ( .A(n52331), .B(n52330), .Y(n52333) );
  NOR2X1 U55131 ( .A(n19222), .B(n19221), .Y(n52332) );
  NAND2X1 U55132 ( .A(n52333), .B(n52332), .Y(u_decode_u_regfile_N775) );
  NOR2X1 U55133 ( .A(n44316), .B(n43121), .Y(n52335) );
  NOR2X1 U55134 ( .A(n44313), .B(n43123), .Y(n52334) );
  NOR2X1 U55135 ( .A(n52335), .B(n52334), .Y(n52337) );
  NOR2X1 U55136 ( .A(n23688), .B(n23687), .Y(n52336) );
  NAND2X1 U55137 ( .A(n52337), .B(n52336), .Y(u_decode_u_regfile_N1071) );
  NOR2X1 U55138 ( .A(n44394), .B(n43121), .Y(n52339) );
  NOR2X1 U55139 ( .A(n44391), .B(n43123), .Y(n52338) );
  NOR2X1 U55140 ( .A(n52339), .B(n52338), .Y(n52341) );
  NOR2X1 U55141 ( .A(n22364), .B(n22363), .Y(n52340) );
  NAND2X1 U55142 ( .A(n52341), .B(n52340), .Y(u_decode_u_regfile_N183) );
  NOR2X1 U55143 ( .A(n44484), .B(n43120), .Y(n52343) );
  NOR2X1 U55144 ( .A(n44481), .B(n43123), .Y(n52342) );
  NOR2X1 U55145 ( .A(n52343), .B(n52342), .Y(n52345) );
  NOR2X1 U55146 ( .A(n20794), .B(n20793), .Y(n52344) );
  NAND2X1 U55147 ( .A(n52345), .B(n52344), .Y(u_decode_u_regfile_N479) );
  NOR2X1 U55148 ( .A(n44418), .B(n43120), .Y(n52347) );
  NOR2X1 U55149 ( .A(n44415), .B(n43123), .Y(n52346) );
  NOR2X1 U55150 ( .A(n52347), .B(n52346), .Y(n52349) );
  NOR2X1 U55151 ( .A(n21972), .B(n21971), .Y(n52348) );
  NAND2X1 U55152 ( .A(n52349), .B(n52348), .Y(u_decode_u_regfile_N257) );
  NOR2X1 U55153 ( .A(n44340), .B(n43120), .Y(n52351) );
  NOR2X1 U55154 ( .A(n44337), .B(n43123), .Y(n52350) );
  NOR2X1 U55155 ( .A(n52351), .B(n52350), .Y(n52353) );
  NOR2X1 U55156 ( .A(n23254), .B(n23253), .Y(n52352) );
  NAND2X1 U55157 ( .A(n52353), .B(n52352), .Y(u_decode_u_regfile_N1145) );
  NOR2X1 U55158 ( .A(n44502), .B(n43120), .Y(n52355) );
  NOR2X1 U55159 ( .A(n44499), .B(n43123), .Y(n52354) );
  NOR2X1 U55160 ( .A(n52355), .B(n52354), .Y(n52357) );
  NOR2X1 U55161 ( .A(n20402), .B(n20401), .Y(n52356) );
  NAND2X1 U55162 ( .A(n52357), .B(n52356), .Y(u_decode_u_regfile_N553) );
  NOR2X1 U55163 ( .A(n44577), .B(n43120), .Y(n52359) );
  NOR2X1 U55164 ( .A(n44574), .B(n43123), .Y(n52358) );
  NOR2X1 U55165 ( .A(n52359), .B(n52358), .Y(n52361) );
  NOR2X1 U55166 ( .A(n18830), .B(n18829), .Y(n52360) );
  NAND2X1 U55167 ( .A(n52361), .B(n52360), .Y(u_decode_u_regfile_N849) );
  NOR2X1 U55168 ( .A(n44526), .B(n43120), .Y(n52363) );
  NOR2X1 U55169 ( .A(n44523), .B(n43123), .Y(n52362) );
  NOR2X1 U55170 ( .A(n52363), .B(n52362), .Y(n52365) );
  NOR2X1 U55171 ( .A(n20010), .B(n20009), .Y(n52364) );
  NAND2X1 U55172 ( .A(n52365), .B(n52364), .Y(u_decode_u_regfile_N627) );
  NOR2X1 U55173 ( .A(n44592), .B(n43120), .Y(n52367) );
  NOR2X1 U55174 ( .A(n44589), .B(n43124), .Y(n52366) );
  NOR2X1 U55175 ( .A(n52367), .B(n52366), .Y(n52369) );
  NOR2X1 U55176 ( .A(n18440), .B(n18439), .Y(n52368) );
  NAND2X1 U55177 ( .A(n52369), .B(n52368), .Y(u_decode_u_regfile_N923) );
  NOR2X1 U55178 ( .A(n44364), .B(n43120), .Y(n52371) );
  NOR2X1 U55179 ( .A(n44361), .B(n43123), .Y(n52370) );
  NOR2X1 U55180 ( .A(n52371), .B(n52370), .Y(n52373) );
  NOR2X1 U55181 ( .A(n22820), .B(n22819), .Y(n52372) );
  NAND2X1 U55182 ( .A(n52373), .B(n52372), .Y(u_decode_u_regfile_N1219) );
  NOR2X1 U55183 ( .A(n44442), .B(n43121), .Y(n52375) );
  NOR2X1 U55184 ( .A(n44439), .B(n43124), .Y(n52374) );
  NOR2X1 U55185 ( .A(n52375), .B(n52374), .Y(n52377) );
  NOR2X1 U55186 ( .A(n21580), .B(n21579), .Y(n52376) );
  NAND2X1 U55187 ( .A(n52377), .B(n52376), .Y(u_decode_u_regfile_N331) );
  NOR2X1 U55188 ( .A(n17196), .B(n17197), .Y(n52379) );
  NOR2X1 U55189 ( .A(n17378), .B(n17379), .Y(n52378) );
  NAND2X1 U55190 ( .A(n52379), .B(n52378), .Y(u_exec_alu_p_w[10]) );
  NOR2X1 U55191 ( .A(n44538), .B(n43126), .Y(n52381) );
  NOR2X1 U55192 ( .A(n44536), .B(n37675), .Y(n52380) );
  NOR2X1 U55193 ( .A(n52381), .B(n52380), .Y(n52383) );
  NOR2X1 U55194 ( .A(n19807), .B(n19806), .Y(n52382) );
  NAND2X1 U55195 ( .A(n52383), .B(n52382), .Y(u_decode_u_regfile_N665) );
  NOR2X1 U55196 ( .A(n44602), .B(n43127), .Y(n52385) );
  NOR2X1 U55197 ( .A(n44599), .B(n37675), .Y(n52384) );
  NOR2X1 U55198 ( .A(n52385), .B(n52384), .Y(n52387) );
  NOR2X1 U55199 ( .A(n18235), .B(n18234), .Y(n52386) );
  NAND2X1 U55200 ( .A(n52387), .B(n52386), .Y(u_decode_u_regfile_N961) );
  NOR2X1 U55201 ( .A(n43125), .B(n43271), .Y(n52389) );
  NOR2X1 U55202 ( .A(n43128), .B(n43387), .Y(n52388) );
  NOR2X1 U55203 ( .A(n52389), .B(n52388), .Y(n52391) );
  NOR2X1 U55204 ( .A(n21377), .B(n21376), .Y(n52390) );
  NAND2X1 U55205 ( .A(n52391), .B(n52390), .Y(u_decode_u_regfile_N369) );
  NOR2X1 U55206 ( .A(n44473), .B(n43127), .Y(n52393) );
  NOR2X1 U55207 ( .A(n44470), .B(n37675), .Y(n52392) );
  NOR2X1 U55208 ( .A(n52393), .B(n52392), .Y(n52395) );
  NOR2X1 U55209 ( .A(n20984), .B(n20983), .Y(n52394) );
  NAND2X1 U55210 ( .A(n52395), .B(n52394), .Y(u_decode_u_regfile_N443) );
  NOR2X1 U55211 ( .A(n44560), .B(n43127), .Y(n52397) );
  NOR2X1 U55212 ( .A(n44557), .B(n37675), .Y(n52396) );
  NOR2X1 U55213 ( .A(n52397), .B(n52396), .Y(n52399) );
  NOR2X1 U55214 ( .A(n19412), .B(n19411), .Y(n52398) );
  NAND2X1 U55215 ( .A(n52399), .B(n52398), .Y(u_decode_u_regfile_N739) );
  NOR2X1 U55216 ( .A(n44383), .B(n43127), .Y(n52401) );
  NOR2X1 U55217 ( .A(n44380), .B(n43129), .Y(n52400) );
  NOR2X1 U55218 ( .A(n52401), .B(n52400), .Y(n52403) );
  NOR2X1 U55219 ( .A(n22554), .B(n22553), .Y(n52402) );
  NAND2X1 U55220 ( .A(n52403), .B(n52402), .Y(u_decode_u_regfile_N147) );
  NOR2X1 U55221 ( .A(n44305), .B(n43127), .Y(n52405) );
  NOR2X1 U55222 ( .A(n44302), .B(n43129), .Y(n52404) );
  NOR2X1 U55223 ( .A(n52405), .B(n52404), .Y(n52407) );
  NOR2X1 U55224 ( .A(n23902), .B(n23901), .Y(n52406) );
  NAND2X1 U55225 ( .A(n52407), .B(n52406), .Y(u_decode_u_regfile_N1035) );
  NOR2X1 U55226 ( .A(n44572), .B(n43127), .Y(n52409) );
  NOR2X1 U55227 ( .A(n44569), .B(n43129), .Y(n52408) );
  NOR2X1 U55228 ( .A(n52409), .B(n52408), .Y(n52411) );
  NOR2X1 U55229 ( .A(n19020), .B(n19019), .Y(n52410) );
  NAND2X1 U55230 ( .A(n52411), .B(n52410), .Y(u_decode_u_regfile_N813) );
  NOR2X1 U55231 ( .A(n43125), .B(n43277), .Y(n52413) );
  NOR2X1 U55232 ( .A(n43128), .B(n43384), .Y(n52412) );
  NOR2X1 U55233 ( .A(n52413), .B(n52412), .Y(n52415) );
  NOR2X1 U55234 ( .A(n20592), .B(n20591), .Y(n52414) );
  NAND2X1 U55235 ( .A(n52415), .B(n52414), .Y(u_decode_u_regfile_N517) );
  NOR2X1 U55236 ( .A(n44407), .B(n43126), .Y(n52417) );
  NOR2X1 U55237 ( .A(n44404), .B(n43129), .Y(n52416) );
  NOR2X1 U55238 ( .A(n52417), .B(n52416), .Y(n52419) );
  NOR2X1 U55239 ( .A(n22162), .B(n22161), .Y(n52418) );
  NAND2X1 U55240 ( .A(n52419), .B(n52418), .Y(u_decode_u_regfile_N221) );
  NOR2X1 U55241 ( .A(n44329), .B(n43126), .Y(n52421) );
  NOR2X1 U55242 ( .A(n44326), .B(n43129), .Y(n52420) );
  NOR2X1 U55243 ( .A(n52421), .B(n52420), .Y(n52423) );
  NOR2X1 U55244 ( .A(n23468), .B(n23467), .Y(n52422) );
  NAND2X1 U55245 ( .A(n52423), .B(n52422), .Y(u_decode_u_regfile_N1109) );
  NOR2X1 U55246 ( .A(n44584), .B(n43126), .Y(n52425) );
  NOR2X1 U55247 ( .A(n44581), .B(n43129), .Y(n52424) );
  NOR2X1 U55248 ( .A(n52425), .B(n52424), .Y(n52427) );
  NOR2X1 U55249 ( .A(n18628), .B(n18627), .Y(n52426) );
  NAND2X1 U55250 ( .A(n52427), .B(n52426), .Y(u_decode_u_regfile_N887) );
  NOR2X1 U55251 ( .A(n44431), .B(n43126), .Y(n52429) );
  NOR2X1 U55252 ( .A(n44428), .B(n43129), .Y(n52428) );
  NOR2X1 U55253 ( .A(n52429), .B(n52428), .Y(n52431) );
  NOR2X1 U55254 ( .A(n21770), .B(n21769), .Y(n52430) );
  NAND2X1 U55255 ( .A(n52431), .B(n52430), .Y(u_decode_u_regfile_N295) );
  NOR2X1 U55256 ( .A(n44515), .B(n43126), .Y(n52433) );
  NOR2X1 U55257 ( .A(n44512), .B(n43129), .Y(n52432) );
  NOR2X1 U55258 ( .A(n52433), .B(n52432), .Y(n52435) );
  NOR2X1 U55259 ( .A(n20200), .B(n20199), .Y(n52434) );
  NAND2X1 U55260 ( .A(n52435), .B(n52434), .Y(u_decode_u_regfile_N591) );
  NOR2X1 U55261 ( .A(n44353), .B(n43126), .Y(n52437) );
  NOR2X1 U55262 ( .A(n44350), .B(n43129), .Y(n52436) );
  NOR2X1 U55263 ( .A(n52437), .B(n52436), .Y(n52439) );
  NOR2X1 U55264 ( .A(n23028), .B(n23027), .Y(n52438) );
  NAND2X1 U55265 ( .A(n52439), .B(n52438), .Y(u_decode_u_regfile_N1183) );
  NOR2X1 U55266 ( .A(n44607), .B(n43126), .Y(n52441) );
  NOR2X1 U55267 ( .A(n44604), .B(n43129), .Y(n52440) );
  NOR2X1 U55268 ( .A(n52441), .B(n52440), .Y(n52443) );
  NOR2X1 U55269 ( .A(n18011), .B(n18009), .Y(n52442) );
  NAND2X1 U55270 ( .A(n52443), .B(n52442), .Y(u_decode_u_regfile_N998) );
  NOR2X1 U55271 ( .A(n43125), .B(n43274), .Y(n52445) );
  NOR2X1 U55272 ( .A(n43128), .B(n43390), .Y(n52444) );
  NOR2X1 U55273 ( .A(n52445), .B(n52444), .Y(n52447) );
  NOR2X1 U55274 ( .A(n23528), .B(n23527), .Y(n52446) );
  NAND2X1 U55275 ( .A(n52447), .B(n52446), .Y(u_decode_u_regfile_N110) );
  NOR2X1 U55276 ( .A(n44461), .B(n43126), .Y(n52449) );
  NOR2X1 U55277 ( .A(n44458), .B(n43129), .Y(n52448) );
  NOR2X1 U55278 ( .A(n52449), .B(n52448), .Y(n52451) );
  NOR2X1 U55279 ( .A(n21180), .B(n21179), .Y(n52450) );
  NAND2X1 U55280 ( .A(n52451), .B(n52450), .Y(u_decode_u_regfile_N406) );
  NOR2X1 U55281 ( .A(n44551), .B(n43126), .Y(n52453) );
  NOR2X1 U55282 ( .A(n44548), .B(n43129), .Y(n52452) );
  NOR2X1 U55283 ( .A(n52453), .B(n52452), .Y(n52455) );
  NOR2X1 U55284 ( .A(n19610), .B(n19609), .Y(n52454) );
  NAND2X1 U55285 ( .A(n52455), .B(n52454), .Y(u_decode_u_regfile_N702) );
  NOR2X1 U55286 ( .A(n44566), .B(n43126), .Y(n52457) );
  NOR2X1 U55287 ( .A(n44563), .B(n43128), .Y(n52456) );
  NOR2X1 U55288 ( .A(n52457), .B(n52456), .Y(n52459) );
  NOR2X1 U55289 ( .A(n19216), .B(n19215), .Y(n52458) );
  NAND2X1 U55290 ( .A(n52459), .B(n52458), .Y(u_decode_u_regfile_N776) );
  NOR2X1 U55291 ( .A(n44317), .B(n43126), .Y(n52461) );
  NOR2X1 U55292 ( .A(n44314), .B(n43128), .Y(n52460) );
  NOR2X1 U55293 ( .A(n52461), .B(n52460), .Y(n52463) );
  NOR2X1 U55294 ( .A(n23682), .B(n23681), .Y(n52462) );
  NAND2X1 U55295 ( .A(n52463), .B(n52462), .Y(u_decode_u_regfile_N1072) );
  NOR2X1 U55296 ( .A(n44395), .B(n43126), .Y(n52465) );
  NOR2X1 U55297 ( .A(n44392), .B(n43128), .Y(n52464) );
  NOR2X1 U55298 ( .A(n52465), .B(n52464), .Y(n52467) );
  NOR2X1 U55299 ( .A(n22358), .B(n22357), .Y(n52466) );
  NAND2X1 U55300 ( .A(n52467), .B(n52466), .Y(u_decode_u_regfile_N184) );
  NOR2X1 U55301 ( .A(n44485), .B(n43125), .Y(n52469) );
  NOR2X1 U55302 ( .A(n44482), .B(n43128), .Y(n52468) );
  NOR2X1 U55303 ( .A(n52469), .B(n52468), .Y(n52471) );
  NOR2X1 U55304 ( .A(n20788), .B(n20787), .Y(n52470) );
  NAND2X1 U55305 ( .A(n52471), .B(n52470), .Y(u_decode_u_regfile_N480) );
  NOR2X1 U55306 ( .A(n44419), .B(n43125), .Y(n52473) );
  NOR2X1 U55307 ( .A(n44416), .B(n43128), .Y(n52472) );
  NOR2X1 U55308 ( .A(n52473), .B(n52472), .Y(n52475) );
  NOR2X1 U55309 ( .A(n21966), .B(n21965), .Y(n52474) );
  NAND2X1 U55310 ( .A(n52475), .B(n52474), .Y(u_decode_u_regfile_N258) );
  NOR2X1 U55311 ( .A(n44341), .B(n43125), .Y(n52477) );
  NOR2X1 U55312 ( .A(n44338), .B(n43128), .Y(n52476) );
  NOR2X1 U55313 ( .A(n52477), .B(n52476), .Y(n52479) );
  NOR2X1 U55314 ( .A(n23248), .B(n23247), .Y(n52478) );
  NAND2X1 U55315 ( .A(n52479), .B(n52478), .Y(u_decode_u_regfile_N1146) );
  NOR2X1 U55316 ( .A(n44503), .B(n43125), .Y(n52481) );
  NOR2X1 U55317 ( .A(n44500), .B(n43128), .Y(n52480) );
  NOR2X1 U55318 ( .A(n52481), .B(n52480), .Y(n52483) );
  NOR2X1 U55319 ( .A(n20396), .B(n20395), .Y(n52482) );
  NAND2X1 U55320 ( .A(n52483), .B(n52482), .Y(u_decode_u_regfile_N554) );
  NOR2X1 U55321 ( .A(n44578), .B(n43125), .Y(n52485) );
  NOR2X1 U55322 ( .A(n44575), .B(n43128), .Y(n52484) );
  NOR2X1 U55323 ( .A(n52485), .B(n52484), .Y(n52487) );
  NOR2X1 U55324 ( .A(n18824), .B(n18823), .Y(n52486) );
  NAND2X1 U55325 ( .A(n52487), .B(n52486), .Y(u_decode_u_regfile_N850) );
  NOR2X1 U55326 ( .A(n44527), .B(n43125), .Y(n52489) );
  NOR2X1 U55327 ( .A(n44524), .B(n43128), .Y(n52488) );
  NOR2X1 U55328 ( .A(n52489), .B(n52488), .Y(n52491) );
  NOR2X1 U55329 ( .A(n20004), .B(n20003), .Y(n52490) );
  NAND2X1 U55330 ( .A(n52491), .B(n52490), .Y(u_decode_u_regfile_N628) );
  NOR2X1 U55331 ( .A(n44593), .B(n43125), .Y(n52493) );
  NOR2X1 U55332 ( .A(n44590), .B(n43129), .Y(n52492) );
  NOR2X1 U55333 ( .A(n52493), .B(n52492), .Y(n52495) );
  NOR2X1 U55334 ( .A(n18434), .B(n18433), .Y(n52494) );
  NAND2X1 U55335 ( .A(n52495), .B(n52494), .Y(u_decode_u_regfile_N924) );
  NOR2X1 U55336 ( .A(n44364), .B(n43125), .Y(n52497) );
  NOR2X1 U55337 ( .A(n44361), .B(n43128), .Y(n52496) );
  NOR2X1 U55338 ( .A(n52497), .B(n52496), .Y(n52499) );
  NOR2X1 U55339 ( .A(n22808), .B(n22807), .Y(n52498) );
  NAND2X1 U55340 ( .A(n52499), .B(n52498), .Y(u_decode_u_regfile_N1220) );
  NOR2X1 U55341 ( .A(n44443), .B(n43126), .Y(n52501) );
  NOR2X1 U55342 ( .A(n44440), .B(n43129), .Y(n52500) );
  NOR2X1 U55343 ( .A(n52501), .B(n52500), .Y(n52503) );
  NOR2X1 U55344 ( .A(n21574), .B(n21573), .Y(n52502) );
  NAND2X1 U55345 ( .A(n52503), .B(n52502), .Y(u_decode_u_regfile_N332) );
  NOR2X1 U55346 ( .A(n17112), .B(n17113), .Y(n52505) );
  NOR2X1 U55347 ( .A(n17164), .B(n17165), .Y(n52504) );
  NAND2X1 U55348 ( .A(n52505), .B(n52504), .Y(u_exec_alu_p_w[11]) );
  NOR2X1 U55349 ( .A(n44538), .B(n43131), .Y(n52507) );
  NOR2X1 U55350 ( .A(n44536), .B(n37676), .Y(n52506) );
  NOR2X1 U55351 ( .A(n52507), .B(n52506), .Y(n52509) );
  NOR2X1 U55352 ( .A(n19801), .B(n19800), .Y(n52508) );
  NAND2X1 U55353 ( .A(n52509), .B(n52508), .Y(u_decode_u_regfile_N666) );
  NOR2X1 U55354 ( .A(n44602), .B(n43132), .Y(n52511) );
  NOR2X1 U55355 ( .A(n44599), .B(n37676), .Y(n52510) );
  NOR2X1 U55356 ( .A(n52511), .B(n52510), .Y(n52513) );
  NOR2X1 U55357 ( .A(n18229), .B(n18228), .Y(n52512) );
  NAND2X1 U55358 ( .A(n52513), .B(n52512), .Y(u_decode_u_regfile_N962) );
  NOR2X1 U55359 ( .A(n43130), .B(n43271), .Y(n52515) );
  NOR2X1 U55360 ( .A(n43133), .B(n43387), .Y(n52514) );
  NOR2X1 U55361 ( .A(n52515), .B(n52514), .Y(n52517) );
  NOR2X1 U55362 ( .A(n21371), .B(n21370), .Y(n52516) );
  NAND2X1 U55363 ( .A(n52517), .B(n52516), .Y(u_decode_u_regfile_N370) );
  NOR2X1 U55364 ( .A(n44473), .B(n43132), .Y(n52519) );
  NOR2X1 U55365 ( .A(n44470), .B(n37676), .Y(n52518) );
  NOR2X1 U55366 ( .A(n52519), .B(n52518), .Y(n52521) );
  NOR2X1 U55367 ( .A(n20978), .B(n20977), .Y(n52520) );
  NAND2X1 U55368 ( .A(n52521), .B(n52520), .Y(u_decode_u_regfile_N444) );
  NOR2X1 U55369 ( .A(n44560), .B(n43132), .Y(n52523) );
  NOR2X1 U55370 ( .A(n44557), .B(n37676), .Y(n52522) );
  NOR2X1 U55371 ( .A(n52523), .B(n52522), .Y(n52525) );
  NOR2X1 U55372 ( .A(n19406), .B(n19405), .Y(n52524) );
  NAND2X1 U55373 ( .A(n52525), .B(n52524), .Y(u_decode_u_regfile_N740) );
  NOR2X1 U55374 ( .A(n44383), .B(n43132), .Y(n52527) );
  NOR2X1 U55375 ( .A(n44380), .B(n43134), .Y(n52526) );
  NOR2X1 U55376 ( .A(n52527), .B(n52526), .Y(n52529) );
  NOR2X1 U55377 ( .A(n22548), .B(n22547), .Y(n52528) );
  NAND2X1 U55378 ( .A(n52529), .B(n52528), .Y(u_decode_u_regfile_N148) );
  NOR2X1 U55379 ( .A(n44305), .B(n43132), .Y(n52531) );
  NOR2X1 U55380 ( .A(n44302), .B(n43134), .Y(n52530) );
  NOR2X1 U55381 ( .A(n52531), .B(n52530), .Y(n52533) );
  NOR2X1 U55382 ( .A(n23896), .B(n23895), .Y(n52532) );
  NAND2X1 U55383 ( .A(n52533), .B(n52532), .Y(u_decode_u_regfile_N1036) );
  NOR2X1 U55384 ( .A(n44572), .B(n43132), .Y(n52535) );
  NOR2X1 U55385 ( .A(n44569), .B(n43134), .Y(n52534) );
  NOR2X1 U55386 ( .A(n52535), .B(n52534), .Y(n52537) );
  NOR2X1 U55387 ( .A(n19014), .B(n19013), .Y(n52536) );
  NAND2X1 U55388 ( .A(n52537), .B(n52536), .Y(u_decode_u_regfile_N814) );
  NOR2X1 U55389 ( .A(n43130), .B(n43277), .Y(n52539) );
  NOR2X1 U55390 ( .A(n43133), .B(n43384), .Y(n52538) );
  NOR2X1 U55391 ( .A(n52539), .B(n52538), .Y(n52541) );
  NOR2X1 U55392 ( .A(n20586), .B(n20585), .Y(n52540) );
  NAND2X1 U55393 ( .A(n52541), .B(n52540), .Y(u_decode_u_regfile_N518) );
  NOR2X1 U55394 ( .A(n44407), .B(n43131), .Y(n52543) );
  NOR2X1 U55395 ( .A(n44404), .B(n43134), .Y(n52542) );
  NOR2X1 U55396 ( .A(n52543), .B(n52542), .Y(n52545) );
  NOR2X1 U55397 ( .A(n22156), .B(n22155), .Y(n52544) );
  NAND2X1 U55398 ( .A(n52545), .B(n52544), .Y(u_decode_u_regfile_N222) );
  NOR2X1 U55399 ( .A(n44329), .B(n43131), .Y(n52547) );
  NOR2X1 U55400 ( .A(n44326), .B(n43134), .Y(n52546) );
  NOR2X1 U55401 ( .A(n52547), .B(n52546), .Y(n52549) );
  NOR2X1 U55402 ( .A(n23456), .B(n23455), .Y(n52548) );
  NAND2X1 U55403 ( .A(n52549), .B(n52548), .Y(u_decode_u_regfile_N1110) );
  NOR2X1 U55404 ( .A(n44584), .B(n43131), .Y(n52551) );
  NOR2X1 U55405 ( .A(n44581), .B(n43134), .Y(n52550) );
  NOR2X1 U55406 ( .A(n52551), .B(n52550), .Y(n52553) );
  NOR2X1 U55407 ( .A(n18622), .B(n18621), .Y(n52552) );
  NAND2X1 U55408 ( .A(n52553), .B(n52552), .Y(u_decode_u_regfile_N888) );
  NOR2X1 U55409 ( .A(n44431), .B(n43131), .Y(n52555) );
  NOR2X1 U55410 ( .A(n44428), .B(n43134), .Y(n52554) );
  NOR2X1 U55411 ( .A(n52555), .B(n52554), .Y(n52557) );
  NOR2X1 U55412 ( .A(n21764), .B(n21763), .Y(n52556) );
  NAND2X1 U55413 ( .A(n52557), .B(n52556), .Y(u_decode_u_regfile_N296) );
  NOR2X1 U55414 ( .A(n44515), .B(n43131), .Y(n52559) );
  NOR2X1 U55415 ( .A(n44512), .B(n43134), .Y(n52558) );
  NOR2X1 U55416 ( .A(n52559), .B(n52558), .Y(n52561) );
  NOR2X1 U55417 ( .A(n20194), .B(n20193), .Y(n52560) );
  NAND2X1 U55418 ( .A(n52561), .B(n52560), .Y(u_decode_u_regfile_N592) );
  NOR2X1 U55419 ( .A(n44353), .B(n43131), .Y(n52563) );
  NOR2X1 U55420 ( .A(n44350), .B(n43134), .Y(n52562) );
  NOR2X1 U55421 ( .A(n52563), .B(n52562), .Y(n52565) );
  NOR2X1 U55422 ( .A(n23022), .B(n23021), .Y(n52564) );
  NAND2X1 U55423 ( .A(n52565), .B(n52564), .Y(u_decode_u_regfile_N1184) );
  NOR2X1 U55424 ( .A(n44608), .B(n43131), .Y(n52567) );
  NOR2X1 U55425 ( .A(n44605), .B(n43134), .Y(n52566) );
  NOR2X1 U55426 ( .A(n52567), .B(n52566), .Y(n52569) );
  NOR2X1 U55427 ( .A(n18003), .B(n18000), .Y(n52568) );
  NAND2X1 U55428 ( .A(n52569), .B(n52568), .Y(u_decode_u_regfile_N999) );
  NOR2X1 U55429 ( .A(n43130), .B(n43274), .Y(n52571) );
  NOR2X1 U55430 ( .A(n43133), .B(n43390), .Y(n52570) );
  NOR2X1 U55431 ( .A(n52571), .B(n52570), .Y(n52573) );
  NOR2X1 U55432 ( .A(n23462), .B(n23461), .Y(n52572) );
  NAND2X1 U55433 ( .A(n52573), .B(n52572), .Y(u_decode_u_regfile_N111) );
  NOR2X1 U55434 ( .A(n44461), .B(n43131), .Y(n52575) );
  NOR2X1 U55435 ( .A(n44458), .B(n43134), .Y(n52574) );
  NOR2X1 U55436 ( .A(n52575), .B(n52574), .Y(n52577) );
  NOR2X1 U55437 ( .A(n21174), .B(n21173), .Y(n52576) );
  NAND2X1 U55438 ( .A(n52577), .B(n52576), .Y(u_decode_u_regfile_N407) );
  NOR2X1 U55439 ( .A(n44551), .B(n43131), .Y(n52579) );
  NOR2X1 U55440 ( .A(n44548), .B(n43134), .Y(n52578) );
  NOR2X1 U55441 ( .A(n52579), .B(n52578), .Y(n52581) );
  NOR2X1 U55442 ( .A(n19604), .B(n19603), .Y(n52580) );
  NAND2X1 U55443 ( .A(n52581), .B(n52580), .Y(u_decode_u_regfile_N703) );
  NOR2X1 U55444 ( .A(n44566), .B(n43131), .Y(n52583) );
  NOR2X1 U55445 ( .A(n44563), .B(n43133), .Y(n52582) );
  NOR2X1 U55446 ( .A(n52583), .B(n52582), .Y(n52585) );
  NOR2X1 U55447 ( .A(n19210), .B(n19209), .Y(n52584) );
  NAND2X1 U55448 ( .A(n52585), .B(n52584), .Y(u_decode_u_regfile_N777) );
  NOR2X1 U55449 ( .A(n44317), .B(n43131), .Y(n52587) );
  NOR2X1 U55450 ( .A(n44314), .B(n43133), .Y(n52586) );
  NOR2X1 U55451 ( .A(n52587), .B(n52586), .Y(n52589) );
  NOR2X1 U55452 ( .A(n23676), .B(n23675), .Y(n52588) );
  NAND2X1 U55453 ( .A(n52589), .B(n52588), .Y(u_decode_u_regfile_N1073) );
  NOR2X1 U55454 ( .A(n44395), .B(n43131), .Y(n52591) );
  NOR2X1 U55455 ( .A(n44392), .B(n43133), .Y(n52590) );
  NOR2X1 U55456 ( .A(n52591), .B(n52590), .Y(n52593) );
  NOR2X1 U55457 ( .A(n22352), .B(n22351), .Y(n52592) );
  NAND2X1 U55458 ( .A(n52593), .B(n52592), .Y(u_decode_u_regfile_N185) );
  NOR2X1 U55459 ( .A(n44485), .B(n43130), .Y(n52595) );
  NOR2X1 U55460 ( .A(n44482), .B(n43133), .Y(n52594) );
  NOR2X1 U55461 ( .A(n52595), .B(n52594), .Y(n52597) );
  NOR2X1 U55462 ( .A(n20782), .B(n20781), .Y(n52596) );
  NAND2X1 U55463 ( .A(n52597), .B(n52596), .Y(u_decode_u_regfile_N481) );
  NOR2X1 U55464 ( .A(n44419), .B(n43130), .Y(n52599) );
  NOR2X1 U55465 ( .A(n44416), .B(n43133), .Y(n52598) );
  NOR2X1 U55466 ( .A(n52599), .B(n52598), .Y(n52601) );
  NOR2X1 U55467 ( .A(n21960), .B(n21959), .Y(n52600) );
  NAND2X1 U55468 ( .A(n52601), .B(n52600), .Y(u_decode_u_regfile_N259) );
  NOR2X1 U55469 ( .A(n44341), .B(n43130), .Y(n52603) );
  NOR2X1 U55470 ( .A(n44338), .B(n43133), .Y(n52602) );
  NOR2X1 U55471 ( .A(n52603), .B(n52602), .Y(n52605) );
  NOR2X1 U55472 ( .A(n23242), .B(n23241), .Y(n52604) );
  NAND2X1 U55473 ( .A(n52605), .B(n52604), .Y(u_decode_u_regfile_N1147) );
  NOR2X1 U55474 ( .A(n44503), .B(n43130), .Y(n52607) );
  NOR2X1 U55475 ( .A(n44500), .B(n43133), .Y(n52606) );
  NOR2X1 U55476 ( .A(n52607), .B(n52606), .Y(n52609) );
  NOR2X1 U55477 ( .A(n20390), .B(n20389), .Y(n52608) );
  NAND2X1 U55478 ( .A(n52609), .B(n52608), .Y(u_decode_u_regfile_N555) );
  NOR2X1 U55479 ( .A(n44578), .B(n43130), .Y(n52611) );
  NOR2X1 U55480 ( .A(n44575), .B(n43133), .Y(n52610) );
  NOR2X1 U55481 ( .A(n52611), .B(n52610), .Y(n52613) );
  NOR2X1 U55482 ( .A(n18818), .B(n18817), .Y(n52612) );
  NAND2X1 U55483 ( .A(n52613), .B(n52612), .Y(u_decode_u_regfile_N851) );
  NOR2X1 U55484 ( .A(n44527), .B(n43130), .Y(n52615) );
  NOR2X1 U55485 ( .A(n44524), .B(n43133), .Y(n52614) );
  NOR2X1 U55486 ( .A(n52615), .B(n52614), .Y(n52617) );
  NOR2X1 U55487 ( .A(n19998), .B(n19997), .Y(n52616) );
  NAND2X1 U55488 ( .A(n52617), .B(n52616), .Y(u_decode_u_regfile_N629) );
  NOR2X1 U55489 ( .A(n44593), .B(n43130), .Y(n52619) );
  NOR2X1 U55490 ( .A(n44590), .B(n43134), .Y(n52618) );
  NOR2X1 U55491 ( .A(n52619), .B(n52618), .Y(n52621) );
  NOR2X1 U55492 ( .A(n18428), .B(n18427), .Y(n52620) );
  NAND2X1 U55493 ( .A(n52621), .B(n52620), .Y(u_decode_u_regfile_N925) );
  NOR2X1 U55494 ( .A(n44364), .B(n43130), .Y(n52623) );
  NOR2X1 U55495 ( .A(n44361), .B(n43133), .Y(n52622) );
  NOR2X1 U55496 ( .A(n52623), .B(n52622), .Y(n52625) );
  NOR2X1 U55497 ( .A(n22802), .B(n22801), .Y(n52624) );
  NAND2X1 U55498 ( .A(n52625), .B(n52624), .Y(u_decode_u_regfile_N1221) );
  NOR2X1 U55499 ( .A(n44443), .B(n43131), .Y(n52627) );
  NOR2X1 U55500 ( .A(n44440), .B(n43134), .Y(n52626) );
  NOR2X1 U55501 ( .A(n52627), .B(n52626), .Y(n52629) );
  NOR2X1 U55502 ( .A(n21568), .B(n21567), .Y(n52628) );
  NAND2X1 U55503 ( .A(n52629), .B(n52628), .Y(u_decode_u_regfile_N333) );
  NAND2X1 U55504 ( .A(n42315), .B(n73573), .Y(n15847) );
  NAND2X1 U55505 ( .A(n56797), .B(n42958), .Y(n52630) );
  NAND2X1 U55506 ( .A(n17052), .B(n52630), .Y(n52631) );
  NOR2X1 U55507 ( .A(n17096), .B(n52631), .Y(n52633) );
  NOR2X1 U55508 ( .A(n17050), .B(n17097), .Y(n52632) );
  NAND2X1 U55509 ( .A(n52633), .B(n52632), .Y(u_exec_alu_p_w[12]) );
  NOR2X1 U55510 ( .A(n44538), .B(n43137), .Y(n52635) );
  NOR2X1 U55511 ( .A(n44536), .B(n37677), .Y(n52634) );
  NOR2X1 U55512 ( .A(n52635), .B(n52634), .Y(n52637) );
  NOR2X1 U55513 ( .A(n19795), .B(n19794), .Y(n52636) );
  NAND2X1 U55514 ( .A(n52637), .B(n52636), .Y(u_decode_u_regfile_N667) );
  NOR2X1 U55515 ( .A(n44602), .B(n43138), .Y(n52639) );
  NOR2X1 U55516 ( .A(n44599), .B(n37677), .Y(n52638) );
  NOR2X1 U55517 ( .A(n52639), .B(n52638), .Y(n52641) );
  NOR2X1 U55518 ( .A(n18223), .B(n18221), .Y(n52640) );
  NAND2X1 U55519 ( .A(n52641), .B(n52640), .Y(u_decode_u_regfile_N963) );
  NOR2X1 U55520 ( .A(n43136), .B(n43271), .Y(n52643) );
  NOR2X1 U55521 ( .A(n43139), .B(n43387), .Y(n52642) );
  NOR2X1 U55522 ( .A(n52643), .B(n52642), .Y(n52645) );
  NOR2X1 U55523 ( .A(n21365), .B(n21364), .Y(n52644) );
  NAND2X1 U55524 ( .A(n52645), .B(n52644), .Y(u_decode_u_regfile_N371) );
  NOR2X1 U55525 ( .A(n44473), .B(n43138), .Y(n52647) );
  NOR2X1 U55526 ( .A(n44470), .B(n37677), .Y(n52646) );
  NOR2X1 U55527 ( .A(n52647), .B(n52646), .Y(n52649) );
  NOR2X1 U55528 ( .A(n20972), .B(n20971), .Y(n52648) );
  NAND2X1 U55529 ( .A(n52649), .B(n52648), .Y(u_decode_u_regfile_N445) );
  NOR2X1 U55530 ( .A(n44560), .B(n43138), .Y(n52651) );
  NOR2X1 U55531 ( .A(n44557), .B(n37677), .Y(n52650) );
  NOR2X1 U55532 ( .A(n52651), .B(n52650), .Y(n52653) );
  NOR2X1 U55533 ( .A(n19400), .B(n19399), .Y(n52652) );
  NAND2X1 U55534 ( .A(n52653), .B(n52652), .Y(u_decode_u_regfile_N741) );
  NOR2X1 U55535 ( .A(n44383), .B(n43138), .Y(n52655) );
  NOR2X1 U55536 ( .A(n44380), .B(n43140), .Y(n52654) );
  NOR2X1 U55537 ( .A(n52655), .B(n52654), .Y(n52657) );
  NOR2X1 U55538 ( .A(n22542), .B(n22541), .Y(n52656) );
  NAND2X1 U55539 ( .A(n52657), .B(n52656), .Y(u_decode_u_regfile_N149) );
  NOR2X1 U55540 ( .A(n44305), .B(n43138), .Y(n52659) );
  NOR2X1 U55541 ( .A(n44302), .B(n43140), .Y(n52658) );
  NOR2X1 U55542 ( .A(n52659), .B(n52658), .Y(n52661) );
  NOR2X1 U55543 ( .A(n23890), .B(n23889), .Y(n52660) );
  NAND2X1 U55544 ( .A(n52661), .B(n52660), .Y(u_decode_u_regfile_N1037) );
  NOR2X1 U55545 ( .A(n44572), .B(n43138), .Y(n52663) );
  NOR2X1 U55546 ( .A(n44569), .B(n43140), .Y(n52662) );
  NOR2X1 U55547 ( .A(n52663), .B(n52662), .Y(n52665) );
  NOR2X1 U55548 ( .A(n19008), .B(n19007), .Y(n52664) );
  NAND2X1 U55549 ( .A(n52665), .B(n52664), .Y(u_decode_u_regfile_N815) );
  NOR2X1 U55550 ( .A(n43136), .B(n43277), .Y(n52667) );
  NOR2X1 U55551 ( .A(n43139), .B(n43384), .Y(n52666) );
  NOR2X1 U55552 ( .A(n52667), .B(n52666), .Y(n52669) );
  NOR2X1 U55553 ( .A(n20580), .B(n20579), .Y(n52668) );
  NAND2X1 U55554 ( .A(n52669), .B(n52668), .Y(u_decode_u_regfile_N519) );
  NOR2X1 U55555 ( .A(n44407), .B(n43137), .Y(n52671) );
  NOR2X1 U55556 ( .A(n44404), .B(n43140), .Y(n52670) );
  NOR2X1 U55557 ( .A(n52671), .B(n52670), .Y(n52673) );
  NOR2X1 U55558 ( .A(n22150), .B(n22149), .Y(n52672) );
  NAND2X1 U55559 ( .A(n52673), .B(n52672), .Y(u_decode_u_regfile_N223) );
  NOR2X1 U55560 ( .A(n44329), .B(n43137), .Y(n52675) );
  NOR2X1 U55561 ( .A(n44326), .B(n43140), .Y(n52674) );
  NOR2X1 U55562 ( .A(n52675), .B(n52674), .Y(n52677) );
  NOR2X1 U55563 ( .A(n23450), .B(n23449), .Y(n52676) );
  NAND2X1 U55564 ( .A(n52677), .B(n52676), .Y(u_decode_u_regfile_N1111) );
  NOR2X1 U55565 ( .A(n44584), .B(n43137), .Y(n52679) );
  NOR2X1 U55566 ( .A(n44581), .B(n43140), .Y(n52678) );
  NOR2X1 U55567 ( .A(n52679), .B(n52678), .Y(n52681) );
  NOR2X1 U55568 ( .A(n18616), .B(n18615), .Y(n52680) );
  NAND2X1 U55569 ( .A(n52681), .B(n52680), .Y(u_decode_u_regfile_N889) );
  NOR2X1 U55570 ( .A(n44431), .B(n43137), .Y(n52683) );
  NOR2X1 U55571 ( .A(n44428), .B(n43140), .Y(n52682) );
  NOR2X1 U55572 ( .A(n52683), .B(n52682), .Y(n52685) );
  NOR2X1 U55573 ( .A(n21758), .B(n21757), .Y(n52684) );
  NAND2X1 U55574 ( .A(n52685), .B(n52684), .Y(u_decode_u_regfile_N297) );
  NOR2X1 U55575 ( .A(n44515), .B(n43137), .Y(n52687) );
  NOR2X1 U55576 ( .A(n44512), .B(n43140), .Y(n52686) );
  NOR2X1 U55577 ( .A(n52687), .B(n52686), .Y(n52689) );
  NOR2X1 U55578 ( .A(n20188), .B(n20187), .Y(n52688) );
  NAND2X1 U55579 ( .A(n52689), .B(n52688), .Y(u_decode_u_regfile_N593) );
  NOR2X1 U55580 ( .A(n44353), .B(n43137), .Y(n52691) );
  NOR2X1 U55581 ( .A(n44350), .B(n43140), .Y(n52690) );
  NOR2X1 U55582 ( .A(n52691), .B(n52690), .Y(n52693) );
  NOR2X1 U55583 ( .A(n23016), .B(n23015), .Y(n52692) );
  NAND2X1 U55584 ( .A(n52693), .B(n52692), .Y(u_decode_u_regfile_N1185) );
  NOR2X1 U55585 ( .A(n44608), .B(n43137), .Y(n52695) );
  NOR2X1 U55586 ( .A(n44605), .B(n43140), .Y(n52694) );
  NOR2X1 U55587 ( .A(n52695), .B(n52694), .Y(n52697) );
  NOR2X1 U55588 ( .A(n24102), .B(n24099), .Y(n52696) );
  NAND2X1 U55589 ( .A(n52697), .B(n52696), .Y(u_decode_u_regfile_N1000) );
  NOR2X1 U55590 ( .A(n43136), .B(n43274), .Y(n52699) );
  NOR2X1 U55591 ( .A(n43139), .B(n43390), .Y(n52698) );
  NOR2X1 U55592 ( .A(n52699), .B(n52698), .Y(n52701) );
  NOR2X1 U55593 ( .A(n23396), .B(n23395), .Y(n52700) );
  NAND2X1 U55594 ( .A(n52701), .B(n52700), .Y(u_decode_u_regfile_N112) );
  NOR2X1 U55595 ( .A(n44461), .B(n43137), .Y(n52703) );
  NOR2X1 U55596 ( .A(n44458), .B(n43140), .Y(n52702) );
  NOR2X1 U55597 ( .A(n52703), .B(n52702), .Y(n52705) );
  NOR2X1 U55598 ( .A(n21168), .B(n21167), .Y(n52704) );
  NAND2X1 U55599 ( .A(n52705), .B(n52704), .Y(u_decode_u_regfile_N408) );
  NOR2X1 U55600 ( .A(n44551), .B(n43137), .Y(n52707) );
  NOR2X1 U55601 ( .A(n44548), .B(n43140), .Y(n52706) );
  NOR2X1 U55602 ( .A(n52707), .B(n52706), .Y(n52709) );
  NOR2X1 U55603 ( .A(n19598), .B(n19597), .Y(n52708) );
  NAND2X1 U55604 ( .A(n52709), .B(n52708), .Y(u_decode_u_regfile_N704) );
  NOR2X1 U55605 ( .A(n44566), .B(n43137), .Y(n52711) );
  NOR2X1 U55606 ( .A(n44563), .B(n43139), .Y(n52710) );
  NOR2X1 U55607 ( .A(n52711), .B(n52710), .Y(n52713) );
  NOR2X1 U55608 ( .A(n19204), .B(n19203), .Y(n52712) );
  NAND2X1 U55609 ( .A(n52713), .B(n52712), .Y(u_decode_u_regfile_N778) );
  NOR2X1 U55610 ( .A(n44317), .B(n43137), .Y(n52715) );
  NOR2X1 U55611 ( .A(n44314), .B(n43139), .Y(n52714) );
  NOR2X1 U55612 ( .A(n52715), .B(n52714), .Y(n52717) );
  NOR2X1 U55613 ( .A(n23670), .B(n23669), .Y(n52716) );
  NAND2X1 U55614 ( .A(n52717), .B(n52716), .Y(u_decode_u_regfile_N1074) );
  NOR2X1 U55615 ( .A(n44395), .B(n43137), .Y(n52719) );
  NOR2X1 U55616 ( .A(n44392), .B(n43139), .Y(n52718) );
  NOR2X1 U55617 ( .A(n52719), .B(n52718), .Y(n52721) );
  NOR2X1 U55618 ( .A(n22346), .B(n22345), .Y(n52720) );
  NAND2X1 U55619 ( .A(n52721), .B(n52720), .Y(u_decode_u_regfile_N186) );
  NOR2X1 U55620 ( .A(n44485), .B(n43136), .Y(n52723) );
  NOR2X1 U55621 ( .A(n44482), .B(n43139), .Y(n52722) );
  NOR2X1 U55622 ( .A(n52723), .B(n52722), .Y(n52725) );
  NOR2X1 U55623 ( .A(n20776), .B(n20775), .Y(n52724) );
  NAND2X1 U55624 ( .A(n52725), .B(n52724), .Y(u_decode_u_regfile_N482) );
  NOR2X1 U55625 ( .A(n44419), .B(n43136), .Y(n52727) );
  NOR2X1 U55626 ( .A(n44416), .B(n43139), .Y(n52726) );
  NOR2X1 U55627 ( .A(n52727), .B(n52726), .Y(n52729) );
  NOR2X1 U55628 ( .A(n21954), .B(n21953), .Y(n52728) );
  NAND2X1 U55629 ( .A(n52729), .B(n52728), .Y(u_decode_u_regfile_N260) );
  NOR2X1 U55630 ( .A(n44341), .B(n43136), .Y(n52731) );
  NOR2X1 U55631 ( .A(n44338), .B(n43139), .Y(n52730) );
  NOR2X1 U55632 ( .A(n52731), .B(n52730), .Y(n52733) );
  NOR2X1 U55633 ( .A(n23236), .B(n23235), .Y(n52732) );
  NAND2X1 U55634 ( .A(n52733), .B(n52732), .Y(u_decode_u_regfile_N1148) );
  NOR2X1 U55635 ( .A(n44503), .B(n43136), .Y(n52735) );
  NOR2X1 U55636 ( .A(n44500), .B(n43139), .Y(n52734) );
  NOR2X1 U55637 ( .A(n52735), .B(n52734), .Y(n52737) );
  NOR2X1 U55638 ( .A(n20384), .B(n20383), .Y(n52736) );
  NAND2X1 U55639 ( .A(n52737), .B(n52736), .Y(u_decode_u_regfile_N556) );
  NOR2X1 U55640 ( .A(n44578), .B(n43136), .Y(n52739) );
  NOR2X1 U55641 ( .A(n44575), .B(n43139), .Y(n52738) );
  NOR2X1 U55642 ( .A(n52739), .B(n52738), .Y(n52741) );
  NOR2X1 U55643 ( .A(n18812), .B(n18811), .Y(n52740) );
  NAND2X1 U55644 ( .A(n52741), .B(n52740), .Y(u_decode_u_regfile_N852) );
  NOR2X1 U55645 ( .A(n44527), .B(n43136), .Y(n52743) );
  NOR2X1 U55646 ( .A(n44524), .B(n43139), .Y(n52742) );
  NOR2X1 U55647 ( .A(n52743), .B(n52742), .Y(n52745) );
  NOR2X1 U55648 ( .A(n19992), .B(n19991), .Y(n52744) );
  NAND2X1 U55649 ( .A(n52745), .B(n52744), .Y(u_decode_u_regfile_N630) );
  NOR2X1 U55650 ( .A(n44593), .B(n43136), .Y(n52747) );
  NOR2X1 U55651 ( .A(n44590), .B(n43140), .Y(n52746) );
  NOR2X1 U55652 ( .A(n52747), .B(n52746), .Y(n52749) );
  NOR2X1 U55653 ( .A(n18422), .B(n18421), .Y(n52748) );
  NAND2X1 U55654 ( .A(n52749), .B(n52748), .Y(u_decode_u_regfile_N926) );
  NOR2X1 U55655 ( .A(n44365), .B(n43136), .Y(n52751) );
  NOR2X1 U55656 ( .A(n44362), .B(n43139), .Y(n52750) );
  NOR2X1 U55657 ( .A(n52751), .B(n52750), .Y(n52753) );
  NOR2X1 U55658 ( .A(n22796), .B(n22795), .Y(n52752) );
  NAND2X1 U55659 ( .A(n52753), .B(n52752), .Y(u_decode_u_regfile_N1222) );
  NOR2X1 U55660 ( .A(n44443), .B(n43137), .Y(n52755) );
  NOR2X1 U55661 ( .A(n44440), .B(n43140), .Y(n52754) );
  NOR2X1 U55662 ( .A(n52755), .B(n52754), .Y(n52757) );
  NOR2X1 U55663 ( .A(n21562), .B(n21561), .Y(n52756) );
  NAND2X1 U55664 ( .A(n52757), .B(n52756), .Y(u_decode_u_regfile_N334) );
  NOR2X1 U55665 ( .A(n16915), .B(n16916), .Y(n52759) );
  NOR2X1 U55666 ( .A(n16955), .B(n16956), .Y(n52758) );
  NAND2X1 U55667 ( .A(n52759), .B(n52758), .Y(u_exec_alu_p_w[14]) );
  NOR2X1 U55668 ( .A(n44538), .B(n43143), .Y(n52761) );
  NOR2X1 U55669 ( .A(n44536), .B(n37678), .Y(n52760) );
  NOR2X1 U55670 ( .A(n52761), .B(n52760), .Y(n52763) );
  NOR2X1 U55671 ( .A(n19783), .B(n19782), .Y(n52762) );
  NAND2X1 U55672 ( .A(n52763), .B(n52762), .Y(u_decode_u_regfile_N669) );
  NOR2X1 U55673 ( .A(n44602), .B(n43144), .Y(n52765) );
  NOR2X1 U55674 ( .A(n44599), .B(n37678), .Y(n52764) );
  NOR2X1 U55675 ( .A(n52765), .B(n52764), .Y(n52767) );
  NOR2X1 U55676 ( .A(n18209), .B(n18207), .Y(n52766) );
  NAND2X1 U55677 ( .A(n52767), .B(n52766), .Y(u_decode_u_regfile_N965) );
  NOR2X1 U55678 ( .A(n43142), .B(n43271), .Y(n52769) );
  NOR2X1 U55679 ( .A(n43145), .B(n43387), .Y(n52768) );
  NOR2X1 U55680 ( .A(n52769), .B(n52768), .Y(n52771) );
  NOR2X1 U55681 ( .A(n21353), .B(n21352), .Y(n52770) );
  NAND2X1 U55682 ( .A(n52771), .B(n52770), .Y(u_decode_u_regfile_N373) );
  NOR2X1 U55683 ( .A(n44473), .B(n43144), .Y(n52773) );
  NOR2X1 U55684 ( .A(n44470), .B(n37678), .Y(n52772) );
  NOR2X1 U55685 ( .A(n52773), .B(n52772), .Y(n52775) );
  NOR2X1 U55686 ( .A(n20960), .B(n20959), .Y(n52774) );
  NAND2X1 U55687 ( .A(n52775), .B(n52774), .Y(u_decode_u_regfile_N447) );
  NOR2X1 U55688 ( .A(n44560), .B(n43144), .Y(n52777) );
  NOR2X1 U55689 ( .A(n44557), .B(n37678), .Y(n52776) );
  NOR2X1 U55690 ( .A(n52777), .B(n52776), .Y(n52779) );
  NOR2X1 U55691 ( .A(n19388), .B(n19387), .Y(n52778) );
  NAND2X1 U55692 ( .A(n52779), .B(n52778), .Y(u_decode_u_regfile_N743) );
  NOR2X1 U55693 ( .A(n44383), .B(n43144), .Y(n52781) );
  NOR2X1 U55694 ( .A(n44380), .B(n43146), .Y(n52780) );
  NOR2X1 U55695 ( .A(n52781), .B(n52780), .Y(n52783) );
  NOR2X1 U55696 ( .A(n22530), .B(n22529), .Y(n52782) );
  NAND2X1 U55697 ( .A(n52783), .B(n52782), .Y(u_decode_u_regfile_N151) );
  NOR2X1 U55698 ( .A(n44305), .B(n43144), .Y(n52785) );
  NOR2X1 U55699 ( .A(n44302), .B(n43146), .Y(n52784) );
  NOR2X1 U55700 ( .A(n52785), .B(n52784), .Y(n52787) );
  NOR2X1 U55701 ( .A(n23878), .B(n23877), .Y(n52786) );
  NAND2X1 U55702 ( .A(n52787), .B(n52786), .Y(u_decode_u_regfile_N1039) );
  NOR2X1 U55703 ( .A(n44572), .B(n43144), .Y(n52789) );
  NOR2X1 U55704 ( .A(n44569), .B(n43146), .Y(n52788) );
  NOR2X1 U55705 ( .A(n52789), .B(n52788), .Y(n52791) );
  NOR2X1 U55706 ( .A(n18996), .B(n18995), .Y(n52790) );
  NAND2X1 U55707 ( .A(n52791), .B(n52790), .Y(u_decode_u_regfile_N817) );
  NOR2X1 U55708 ( .A(n43142), .B(n43277), .Y(n52793) );
  NOR2X1 U55709 ( .A(n43145), .B(n43384), .Y(n52792) );
  NOR2X1 U55710 ( .A(n52793), .B(n52792), .Y(n52795) );
  NOR2X1 U55711 ( .A(n20568), .B(n20567), .Y(n52794) );
  NAND2X1 U55712 ( .A(n52795), .B(n52794), .Y(u_decode_u_regfile_N521) );
  NOR2X1 U55713 ( .A(n44407), .B(n43143), .Y(n52797) );
  NOR2X1 U55714 ( .A(n44404), .B(n43146), .Y(n52796) );
  NOR2X1 U55715 ( .A(n52797), .B(n52796), .Y(n52799) );
  NOR2X1 U55716 ( .A(n22138), .B(n22137), .Y(n52798) );
  NAND2X1 U55717 ( .A(n52799), .B(n52798), .Y(u_decode_u_regfile_N225) );
  NOR2X1 U55718 ( .A(n44329), .B(n43143), .Y(n52801) );
  NOR2X1 U55719 ( .A(n44326), .B(n43146), .Y(n52800) );
  NOR2X1 U55720 ( .A(n52801), .B(n52800), .Y(n52803) );
  NOR2X1 U55721 ( .A(n23438), .B(n23437), .Y(n52802) );
  NAND2X1 U55722 ( .A(n52803), .B(n52802), .Y(u_decode_u_regfile_N1113) );
  NOR2X1 U55723 ( .A(n44584), .B(n43143), .Y(n52805) );
  NOR2X1 U55724 ( .A(n44581), .B(n43146), .Y(n52804) );
  NOR2X1 U55725 ( .A(n52805), .B(n52804), .Y(n52807) );
  NOR2X1 U55726 ( .A(n18604), .B(n18603), .Y(n52806) );
  NAND2X1 U55727 ( .A(n52807), .B(n52806), .Y(u_decode_u_regfile_N891) );
  NOR2X1 U55728 ( .A(n44431), .B(n43143), .Y(n52809) );
  NOR2X1 U55729 ( .A(n44428), .B(n43146), .Y(n52808) );
  NOR2X1 U55730 ( .A(n52809), .B(n52808), .Y(n52811) );
  NOR2X1 U55731 ( .A(n21746), .B(n21745), .Y(n52810) );
  NAND2X1 U55732 ( .A(n52811), .B(n52810), .Y(u_decode_u_regfile_N299) );
  NOR2X1 U55733 ( .A(n44515), .B(n43143), .Y(n52813) );
  NOR2X1 U55734 ( .A(n44512), .B(n43146), .Y(n52812) );
  NOR2X1 U55735 ( .A(n52813), .B(n52812), .Y(n52815) );
  NOR2X1 U55736 ( .A(n20176), .B(n20175), .Y(n52814) );
  NAND2X1 U55737 ( .A(n52815), .B(n52814), .Y(u_decode_u_regfile_N595) );
  NOR2X1 U55738 ( .A(n44353), .B(n43143), .Y(n52817) );
  NOR2X1 U55739 ( .A(n44350), .B(n43146), .Y(n52816) );
  NOR2X1 U55740 ( .A(n52817), .B(n52816), .Y(n52819) );
  NOR2X1 U55741 ( .A(n23004), .B(n23003), .Y(n52818) );
  NAND2X1 U55742 ( .A(n52819), .B(n52818), .Y(u_decode_u_regfile_N1187) );
  NOR2X1 U55743 ( .A(n44608), .B(n43143), .Y(n52821) );
  NOR2X1 U55744 ( .A(n44605), .B(n43146), .Y(n52820) );
  NOR2X1 U55745 ( .A(n52821), .B(n52820), .Y(n52823) );
  NOR2X1 U55746 ( .A(n24088), .B(n24087), .Y(n52822) );
  NAND2X1 U55747 ( .A(n52823), .B(n52822), .Y(u_decode_u_regfile_N1002) );
  NOR2X1 U55748 ( .A(n43142), .B(n43274), .Y(n52825) );
  NOR2X1 U55749 ( .A(n43145), .B(n43390), .Y(n52824) );
  NOR2X1 U55750 ( .A(n52825), .B(n52824), .Y(n52827) );
  NOR2X1 U55751 ( .A(n23290), .B(n23289), .Y(n52826) );
  NAND2X1 U55752 ( .A(n52827), .B(n52826), .Y(u_decode_u_regfile_N114) );
  NOR2X1 U55753 ( .A(n44461), .B(n43143), .Y(n52829) );
  NOR2X1 U55754 ( .A(n44458), .B(n43146), .Y(n52828) );
  NOR2X1 U55755 ( .A(n52829), .B(n52828), .Y(n52831) );
  NOR2X1 U55756 ( .A(n21156), .B(n21155), .Y(n52830) );
  NAND2X1 U55757 ( .A(n52831), .B(n52830), .Y(u_decode_u_regfile_N410) );
  NOR2X1 U55758 ( .A(n44551), .B(n43143), .Y(n52833) );
  NOR2X1 U55759 ( .A(n44548), .B(n43146), .Y(n52832) );
  NOR2X1 U55760 ( .A(n52833), .B(n52832), .Y(n52835) );
  NOR2X1 U55761 ( .A(n19586), .B(n19585), .Y(n52834) );
  NAND2X1 U55762 ( .A(n52835), .B(n52834), .Y(u_decode_u_regfile_N706) );
  NOR2X1 U55763 ( .A(n44566), .B(n43143), .Y(n52837) );
  NOR2X1 U55764 ( .A(n44563), .B(n43145), .Y(n52836) );
  NOR2X1 U55765 ( .A(n52837), .B(n52836), .Y(n52839) );
  NOR2X1 U55766 ( .A(n19192), .B(n19191), .Y(n52838) );
  NAND2X1 U55767 ( .A(n52839), .B(n52838), .Y(u_decode_u_regfile_N780) );
  NOR2X1 U55768 ( .A(n44317), .B(n43143), .Y(n52841) );
  NOR2X1 U55769 ( .A(n44314), .B(n43145), .Y(n52840) );
  NOR2X1 U55770 ( .A(n52841), .B(n52840), .Y(n52843) );
  NOR2X1 U55771 ( .A(n23658), .B(n23657), .Y(n52842) );
  NAND2X1 U55772 ( .A(n52843), .B(n52842), .Y(u_decode_u_regfile_N1076) );
  NOR2X1 U55773 ( .A(n44395), .B(n43143), .Y(n52845) );
  NOR2X1 U55774 ( .A(n44392), .B(n43145), .Y(n52844) );
  NOR2X1 U55775 ( .A(n52845), .B(n52844), .Y(n52847) );
  NOR2X1 U55776 ( .A(n22334), .B(n22333), .Y(n52846) );
  NAND2X1 U55777 ( .A(n52847), .B(n52846), .Y(u_decode_u_regfile_N188) );
  NOR2X1 U55778 ( .A(n44485), .B(n43142), .Y(n52849) );
  NOR2X1 U55779 ( .A(n44482), .B(n43145), .Y(n52848) );
  NOR2X1 U55780 ( .A(n52849), .B(n52848), .Y(n52851) );
  NOR2X1 U55781 ( .A(n20764), .B(n20763), .Y(n52850) );
  NAND2X1 U55782 ( .A(n52851), .B(n52850), .Y(u_decode_u_regfile_N484) );
  NOR2X1 U55783 ( .A(n44419), .B(n43142), .Y(n52853) );
  NOR2X1 U55784 ( .A(n44416), .B(n43145), .Y(n52852) );
  NOR2X1 U55785 ( .A(n52853), .B(n52852), .Y(n52855) );
  NOR2X1 U55786 ( .A(n21942), .B(n21941), .Y(n52854) );
  NAND2X1 U55787 ( .A(n52855), .B(n52854), .Y(u_decode_u_regfile_N262) );
  NOR2X1 U55788 ( .A(n44341), .B(n43142), .Y(n52857) );
  NOR2X1 U55789 ( .A(n44338), .B(n43145), .Y(n52856) );
  NOR2X1 U55790 ( .A(n52857), .B(n52856), .Y(n52859) );
  NOR2X1 U55791 ( .A(n23218), .B(n23217), .Y(n52858) );
  NAND2X1 U55792 ( .A(n52859), .B(n52858), .Y(u_decode_u_regfile_N1150) );
  NOR2X1 U55793 ( .A(n44503), .B(n43142), .Y(n52861) );
  NOR2X1 U55794 ( .A(n44500), .B(n43145), .Y(n52860) );
  NOR2X1 U55795 ( .A(n52861), .B(n52860), .Y(n52863) );
  NOR2X1 U55796 ( .A(n20372), .B(n20371), .Y(n52862) );
  NAND2X1 U55797 ( .A(n52863), .B(n52862), .Y(u_decode_u_regfile_N558) );
  NOR2X1 U55798 ( .A(n44578), .B(n43142), .Y(n52865) );
  NOR2X1 U55799 ( .A(n44575), .B(n43145), .Y(n52864) );
  NOR2X1 U55800 ( .A(n52865), .B(n52864), .Y(n52867) );
  NOR2X1 U55801 ( .A(n18800), .B(n18799), .Y(n52866) );
  NAND2X1 U55802 ( .A(n52867), .B(n52866), .Y(u_decode_u_regfile_N854) );
  NOR2X1 U55803 ( .A(n44527), .B(n43142), .Y(n52869) );
  NOR2X1 U55804 ( .A(n44524), .B(n43145), .Y(n52868) );
  NOR2X1 U55805 ( .A(n52869), .B(n52868), .Y(n52871) );
  NOR2X1 U55806 ( .A(n19980), .B(n19979), .Y(n52870) );
  NAND2X1 U55807 ( .A(n52871), .B(n52870), .Y(u_decode_u_regfile_N632) );
  NOR2X1 U55808 ( .A(n44593), .B(n43142), .Y(n52873) );
  NOR2X1 U55809 ( .A(n44590), .B(n43146), .Y(n52872) );
  NOR2X1 U55810 ( .A(n52873), .B(n52872), .Y(n52875) );
  NOR2X1 U55811 ( .A(n18410), .B(n18409), .Y(n52874) );
  NAND2X1 U55812 ( .A(n52875), .B(n52874), .Y(u_decode_u_regfile_N928) );
  NOR2X1 U55813 ( .A(n44365), .B(n43142), .Y(n52877) );
  NOR2X1 U55814 ( .A(n44362), .B(n43145), .Y(n52876) );
  NOR2X1 U55815 ( .A(n52877), .B(n52876), .Y(n52879) );
  NOR2X1 U55816 ( .A(n22784), .B(n22783), .Y(n52878) );
  NAND2X1 U55817 ( .A(n52879), .B(n52878), .Y(u_decode_u_regfile_N1224) );
  NOR2X1 U55818 ( .A(n44443), .B(n43143), .Y(n52881) );
  NOR2X1 U55819 ( .A(n44440), .B(n43146), .Y(n52880) );
  NOR2X1 U55820 ( .A(n52881), .B(n52880), .Y(n52883) );
  NOR2X1 U55821 ( .A(n21550), .B(n21549), .Y(n52882) );
  NAND2X1 U55822 ( .A(n52883), .B(n52882), .Y(u_decode_u_regfile_N336) );
  NOR2X1 U55823 ( .A(n16808), .B(n16809), .Y(n52885) );
  NOR2X1 U55824 ( .A(n16846), .B(n16847), .Y(n52884) );
  NAND2X1 U55825 ( .A(n52885), .B(n52884), .Y(u_exec_alu_p_w[16]) );
  NOR2X1 U55826 ( .A(n44538), .B(n43150), .Y(n52887) );
  NOR2X1 U55827 ( .A(n44536), .B(n37679), .Y(n52886) );
  NOR2X1 U55828 ( .A(n52887), .B(n52886), .Y(n52889) );
  NOR2X1 U55829 ( .A(n19771), .B(n19770), .Y(n52888) );
  NAND2X1 U55830 ( .A(n52889), .B(n52888), .Y(u_decode_u_regfile_N671) );
  NOR2X1 U55831 ( .A(n44602), .B(n43150), .Y(n52891) );
  NOR2X1 U55832 ( .A(n44599), .B(n37679), .Y(n52890) );
  NOR2X1 U55833 ( .A(n52891), .B(n52890), .Y(n52893) );
  NOR2X1 U55834 ( .A(n18195), .B(n18193), .Y(n52892) );
  NAND2X1 U55835 ( .A(n52893), .B(n52892), .Y(u_decode_u_regfile_N967) );
  NOR2X1 U55836 ( .A(n43148), .B(n43271), .Y(n52895) );
  NOR2X1 U55837 ( .A(n43151), .B(n43387), .Y(n52894) );
  NOR2X1 U55838 ( .A(n52895), .B(n52894), .Y(n52897) );
  NOR2X1 U55839 ( .A(n21341), .B(n21340), .Y(n52896) );
  NAND2X1 U55840 ( .A(n52897), .B(n52896), .Y(u_decode_u_regfile_N375) );
  NOR2X1 U55841 ( .A(n44473), .B(n43150), .Y(n52899) );
  NOR2X1 U55842 ( .A(n44470), .B(n37679), .Y(n52898) );
  NOR2X1 U55843 ( .A(n52899), .B(n52898), .Y(n52901) );
  NOR2X1 U55844 ( .A(n20948), .B(n20947), .Y(n52900) );
  NAND2X1 U55845 ( .A(n52901), .B(n52900), .Y(u_decode_u_regfile_N449) );
  NOR2X1 U55846 ( .A(n44560), .B(n43150), .Y(n52903) );
  NOR2X1 U55847 ( .A(n44557), .B(n37679), .Y(n52902) );
  NOR2X1 U55848 ( .A(n52903), .B(n52902), .Y(n52905) );
  NOR2X1 U55849 ( .A(n19376), .B(n19375), .Y(n52904) );
  NAND2X1 U55850 ( .A(n52905), .B(n52904), .Y(u_decode_u_regfile_N745) );
  NOR2X1 U55851 ( .A(n44383), .B(n43149), .Y(n52907) );
  NOR2X1 U55852 ( .A(n44380), .B(n43152), .Y(n52906) );
  NOR2X1 U55853 ( .A(n52907), .B(n52906), .Y(n52909) );
  NOR2X1 U55854 ( .A(n22518), .B(n22517), .Y(n52908) );
  NAND2X1 U55855 ( .A(n52909), .B(n52908), .Y(u_decode_u_regfile_N153) );
  NOR2X1 U55856 ( .A(n44305), .B(n43149), .Y(n52911) );
  NOR2X1 U55857 ( .A(n44302), .B(n43152), .Y(n52910) );
  NOR2X1 U55858 ( .A(n52911), .B(n52910), .Y(n52913) );
  NOR2X1 U55859 ( .A(n23860), .B(n23859), .Y(n52912) );
  NAND2X1 U55860 ( .A(n52913), .B(n52912), .Y(u_decode_u_regfile_N1041) );
  NOR2X1 U55861 ( .A(n44572), .B(n43149), .Y(n52915) );
  NOR2X1 U55862 ( .A(n44569), .B(n43152), .Y(n52914) );
  NOR2X1 U55863 ( .A(n52915), .B(n52914), .Y(n52917) );
  NOR2X1 U55864 ( .A(n18984), .B(n18983), .Y(n52916) );
  NAND2X1 U55865 ( .A(n52917), .B(n52916), .Y(u_decode_u_regfile_N819) );
  NOR2X1 U55866 ( .A(n43148), .B(n43277), .Y(n52919) );
  NOR2X1 U55867 ( .A(n43151), .B(n43384), .Y(n52918) );
  NOR2X1 U55868 ( .A(n52919), .B(n52918), .Y(n52921) );
  NOR2X1 U55869 ( .A(n20556), .B(n20555), .Y(n52920) );
  NAND2X1 U55870 ( .A(n52921), .B(n52920), .Y(u_decode_u_regfile_N523) );
  NOR2X1 U55871 ( .A(n44407), .B(n43149), .Y(n52923) );
  NOR2X1 U55872 ( .A(n44404), .B(n43152), .Y(n52922) );
  NOR2X1 U55873 ( .A(n52923), .B(n52922), .Y(n52925) );
  NOR2X1 U55874 ( .A(n22126), .B(n22125), .Y(n52924) );
  NAND2X1 U55875 ( .A(n52925), .B(n52924), .Y(u_decode_u_regfile_N227) );
  NOR2X1 U55876 ( .A(n44329), .B(n43149), .Y(n52927) );
  NOR2X1 U55877 ( .A(n44326), .B(n43152), .Y(n52926) );
  NOR2X1 U55878 ( .A(n52927), .B(n52926), .Y(n52929) );
  NOR2X1 U55879 ( .A(n23426), .B(n23425), .Y(n52928) );
  NAND2X1 U55880 ( .A(n52929), .B(n52928), .Y(u_decode_u_regfile_N1115) );
  NOR2X1 U55881 ( .A(n44584), .B(n43149), .Y(n52931) );
  NOR2X1 U55882 ( .A(n44581), .B(n43152), .Y(n52930) );
  NOR2X1 U55883 ( .A(n52931), .B(n52930), .Y(n52933) );
  NOR2X1 U55884 ( .A(n18592), .B(n18591), .Y(n52932) );
  NAND2X1 U55885 ( .A(n52933), .B(n52932), .Y(u_decode_u_regfile_N893) );
  NOR2X1 U55886 ( .A(n44431), .B(n43149), .Y(n52935) );
  NOR2X1 U55887 ( .A(n44428), .B(n43152), .Y(n52934) );
  NOR2X1 U55888 ( .A(n52935), .B(n52934), .Y(n52937) );
  NOR2X1 U55889 ( .A(n21734), .B(n21733), .Y(n52936) );
  NAND2X1 U55890 ( .A(n52937), .B(n52936), .Y(u_decode_u_regfile_N301) );
  NOR2X1 U55891 ( .A(n44515), .B(n43149), .Y(n52939) );
  NOR2X1 U55892 ( .A(n44512), .B(n43152), .Y(n52938) );
  NOR2X1 U55893 ( .A(n52939), .B(n52938), .Y(n52941) );
  NOR2X1 U55894 ( .A(n20164), .B(n20163), .Y(n52940) );
  NAND2X1 U55895 ( .A(n52941), .B(n52940), .Y(u_decode_u_regfile_N597) );
  NOR2X1 U55896 ( .A(n44353), .B(n43149), .Y(n52943) );
  NOR2X1 U55897 ( .A(n44350), .B(n43152), .Y(n52942) );
  NOR2X1 U55898 ( .A(n52943), .B(n52942), .Y(n52945) );
  NOR2X1 U55899 ( .A(n22992), .B(n22991), .Y(n52944) );
  NAND2X1 U55900 ( .A(n52945), .B(n52944), .Y(u_decode_u_regfile_N1189) );
  NOR2X1 U55901 ( .A(n44608), .B(n43149), .Y(n52947) );
  NOR2X1 U55902 ( .A(n44605), .B(n43152), .Y(n52946) );
  NOR2X1 U55903 ( .A(n52947), .B(n52946), .Y(n52949) );
  NOR2X1 U55904 ( .A(n24076), .B(n24075), .Y(n52948) );
  NAND2X1 U55905 ( .A(n52949), .B(n52948), .Y(u_decode_u_regfile_N1004) );
  NOR2X1 U55906 ( .A(n43148), .B(n43274), .Y(n52951) );
  NOR2X1 U55907 ( .A(n43151), .B(n43390), .Y(n52950) );
  NOR2X1 U55908 ( .A(n52951), .B(n52950), .Y(n52953) );
  NOR2X1 U55909 ( .A(n23158), .B(n23157), .Y(n52952) );
  NAND2X1 U55910 ( .A(n52953), .B(n52952), .Y(u_decode_u_regfile_N116) );
  NOR2X1 U55911 ( .A(n44461), .B(n43149), .Y(n52955) );
  NOR2X1 U55912 ( .A(n44458), .B(n43152), .Y(n52954) );
  NOR2X1 U55913 ( .A(n52955), .B(n52954), .Y(n52957) );
  NOR2X1 U55914 ( .A(n21144), .B(n21143), .Y(n52956) );
  NAND2X1 U55915 ( .A(n52957), .B(n52956), .Y(u_decode_u_regfile_N412) );
  NOR2X1 U55916 ( .A(n44551), .B(n43149), .Y(n52959) );
  NOR2X1 U55917 ( .A(n44548), .B(n43152), .Y(n52958) );
  NOR2X1 U55918 ( .A(n52959), .B(n52958), .Y(n52961) );
  NOR2X1 U55919 ( .A(n19574), .B(n19573), .Y(n52960) );
  NAND2X1 U55920 ( .A(n52961), .B(n52960), .Y(u_decode_u_regfile_N708) );
  NOR2X1 U55921 ( .A(n44566), .B(n43148), .Y(n52963) );
  NOR2X1 U55922 ( .A(n44563), .B(n43151), .Y(n52962) );
  NOR2X1 U55923 ( .A(n52963), .B(n52962), .Y(n52965) );
  NOR2X1 U55924 ( .A(n19180), .B(n19179), .Y(n52964) );
  NAND2X1 U55925 ( .A(n52965), .B(n52964), .Y(u_decode_u_regfile_N782) );
  NOR2X1 U55926 ( .A(n44317), .B(n43148), .Y(n52967) );
  NOR2X1 U55927 ( .A(n44314), .B(n43151), .Y(n52966) );
  NOR2X1 U55928 ( .A(n52967), .B(n52966), .Y(n52969) );
  NOR2X1 U55929 ( .A(n23646), .B(n23645), .Y(n52968) );
  NAND2X1 U55930 ( .A(n52969), .B(n52968), .Y(u_decode_u_regfile_N1078) );
  NOR2X1 U55931 ( .A(n44395), .B(n43148), .Y(n52971) );
  NOR2X1 U55932 ( .A(n44392), .B(n43151), .Y(n52970) );
  NOR2X1 U55933 ( .A(n52971), .B(n52970), .Y(n52973) );
  NOR2X1 U55934 ( .A(n22322), .B(n22321), .Y(n52972) );
  NAND2X1 U55935 ( .A(n52973), .B(n52972), .Y(u_decode_u_regfile_N190) );
  NOR2X1 U55936 ( .A(n44485), .B(n43149), .Y(n52975) );
  NOR2X1 U55937 ( .A(n44482), .B(n43151), .Y(n52974) );
  NOR2X1 U55938 ( .A(n52975), .B(n52974), .Y(n52977) );
  NOR2X1 U55939 ( .A(n20752), .B(n20751), .Y(n52976) );
  NAND2X1 U55940 ( .A(n52977), .B(n52976), .Y(u_decode_u_regfile_N486) );
  NOR2X1 U55941 ( .A(n44419), .B(n43148), .Y(n52979) );
  NOR2X1 U55942 ( .A(n44416), .B(n43151), .Y(n52978) );
  NOR2X1 U55943 ( .A(n52979), .B(n52978), .Y(n52981) );
  NOR2X1 U55944 ( .A(n21930), .B(n21929), .Y(n52980) );
  NAND2X1 U55945 ( .A(n52981), .B(n52980), .Y(u_decode_u_regfile_N264) );
  NOR2X1 U55946 ( .A(n44341), .B(n43148), .Y(n52983) );
  NOR2X1 U55947 ( .A(n44338), .B(n43151), .Y(n52982) );
  NOR2X1 U55948 ( .A(n52983), .B(n52982), .Y(n52985) );
  NOR2X1 U55949 ( .A(n23206), .B(n23205), .Y(n52984) );
  NAND2X1 U55950 ( .A(n52985), .B(n52984), .Y(u_decode_u_regfile_N1152) );
  NOR2X1 U55951 ( .A(n44503), .B(n43148), .Y(n52987) );
  NOR2X1 U55952 ( .A(n44500), .B(n43151), .Y(n52986) );
  NOR2X1 U55953 ( .A(n52987), .B(n52986), .Y(n52989) );
  NOR2X1 U55954 ( .A(n20360), .B(n20359), .Y(n52988) );
  NAND2X1 U55955 ( .A(n52989), .B(n52988), .Y(u_decode_u_regfile_N560) );
  NOR2X1 U55956 ( .A(n44578), .B(n43148), .Y(n52991) );
  NOR2X1 U55957 ( .A(n44575), .B(n43151), .Y(n52990) );
  NOR2X1 U55958 ( .A(n52991), .B(n52990), .Y(n52993) );
  NOR2X1 U55959 ( .A(n18788), .B(n18787), .Y(n52992) );
  NAND2X1 U55960 ( .A(n52993), .B(n52992), .Y(u_decode_u_regfile_N856) );
  NOR2X1 U55961 ( .A(n44527), .B(n43148), .Y(n52995) );
  NOR2X1 U55962 ( .A(n44524), .B(n43151), .Y(n52994) );
  NOR2X1 U55963 ( .A(n52995), .B(n52994), .Y(n52997) );
  NOR2X1 U55964 ( .A(n19968), .B(n19967), .Y(n52996) );
  NAND2X1 U55965 ( .A(n52997), .B(n52996), .Y(u_decode_u_regfile_N634) );
  NOR2X1 U55966 ( .A(n44593), .B(n43148), .Y(n52999) );
  NOR2X1 U55967 ( .A(n44590), .B(n43152), .Y(n52998) );
  NOR2X1 U55968 ( .A(n52999), .B(n52998), .Y(n53001) );
  NOR2X1 U55969 ( .A(n18398), .B(n18397), .Y(n53000) );
  NAND2X1 U55970 ( .A(n53001), .B(n53000), .Y(u_decode_u_regfile_N930) );
  NOR2X1 U55971 ( .A(n44365), .B(n43148), .Y(n53003) );
  NOR2X1 U55972 ( .A(n44362), .B(n43151), .Y(n53002) );
  NOR2X1 U55973 ( .A(n53003), .B(n53002), .Y(n53005) );
  NOR2X1 U55974 ( .A(n22772), .B(n22771), .Y(n53004) );
  NAND2X1 U55975 ( .A(n53005), .B(n53004), .Y(u_decode_u_regfile_N1226) );
  NOR2X1 U55976 ( .A(n44443), .B(n43149), .Y(n53007) );
  NOR2X1 U55977 ( .A(n44440), .B(n43152), .Y(n53006) );
  NOR2X1 U55978 ( .A(n53007), .B(n53006), .Y(n53009) );
  NOR2X1 U55979 ( .A(n21538), .B(n21537), .Y(n53008) );
  NAND2X1 U55980 ( .A(n53009), .B(n53008), .Y(u_decode_u_regfile_N338) );
  NOR2X1 U55981 ( .A(n16755), .B(n16756), .Y(n53011) );
  NOR2X1 U55982 ( .A(n16794), .B(n16795), .Y(n53010) );
  NAND2X1 U55983 ( .A(n53011), .B(n53010), .Y(u_exec_alu_p_w[17]) );
  NOR2X1 U55984 ( .A(n44538), .B(n43156), .Y(n53013) );
  NOR2X1 U55985 ( .A(n44536), .B(n37680), .Y(n53012) );
  NOR2X1 U55986 ( .A(n53013), .B(n53012), .Y(n53015) );
  NOR2X1 U55987 ( .A(n19765), .B(n19764), .Y(n53014) );
  NAND2X1 U55988 ( .A(n53015), .B(n53014), .Y(u_decode_u_regfile_N672) );
  NOR2X1 U55989 ( .A(n44602), .B(n43156), .Y(n53017) );
  NOR2X1 U55990 ( .A(n44599), .B(n37680), .Y(n53016) );
  NOR2X1 U55991 ( .A(n53017), .B(n53016), .Y(n53019) );
  NOR2X1 U55992 ( .A(n18188), .B(n18186), .Y(n53018) );
  NAND2X1 U55993 ( .A(n53019), .B(n53018), .Y(u_decode_u_regfile_N968) );
  NOR2X1 U55994 ( .A(n43154), .B(n43271), .Y(n53021) );
  NOR2X1 U55995 ( .A(n43157), .B(n43387), .Y(n53020) );
  NOR2X1 U55996 ( .A(n53021), .B(n53020), .Y(n53023) );
  NOR2X1 U55997 ( .A(n21335), .B(n21334), .Y(n53022) );
  NAND2X1 U55998 ( .A(n53023), .B(n53022), .Y(u_decode_u_regfile_N376) );
  NOR2X1 U55999 ( .A(n44473), .B(n43156), .Y(n53025) );
  NOR2X1 U56000 ( .A(n44470), .B(n37680), .Y(n53024) );
  NOR2X1 U56001 ( .A(n53025), .B(n53024), .Y(n53027) );
  NOR2X1 U56002 ( .A(n20942), .B(n20941), .Y(n53026) );
  NAND2X1 U56003 ( .A(n53027), .B(n53026), .Y(u_decode_u_regfile_N450) );
  NOR2X1 U56004 ( .A(n44560), .B(n43156), .Y(n53029) );
  NOR2X1 U56005 ( .A(n44557), .B(n37680), .Y(n53028) );
  NOR2X1 U56006 ( .A(n53029), .B(n53028), .Y(n53031) );
  NOR2X1 U56007 ( .A(n19370), .B(n19369), .Y(n53030) );
  NAND2X1 U56008 ( .A(n53031), .B(n53030), .Y(u_decode_u_regfile_N746) );
  NOR2X1 U56009 ( .A(n44383), .B(n43155), .Y(n53033) );
  NOR2X1 U56010 ( .A(n44380), .B(n43158), .Y(n53032) );
  NOR2X1 U56011 ( .A(n53033), .B(n53032), .Y(n53035) );
  NOR2X1 U56012 ( .A(n22512), .B(n22511), .Y(n53034) );
  NAND2X1 U56013 ( .A(n53035), .B(n53034), .Y(u_decode_u_regfile_N154) );
  NOR2X1 U56014 ( .A(n44305), .B(n43155), .Y(n53037) );
  NOR2X1 U56015 ( .A(n44302), .B(n43158), .Y(n53036) );
  NOR2X1 U56016 ( .A(n53037), .B(n53036), .Y(n53039) );
  NOR2X1 U56017 ( .A(n23854), .B(n23853), .Y(n53038) );
  NAND2X1 U56018 ( .A(n53039), .B(n53038), .Y(u_decode_u_regfile_N1042) );
  NOR2X1 U56019 ( .A(n44572), .B(n43155), .Y(n53041) );
  NOR2X1 U56020 ( .A(n44569), .B(n43158), .Y(n53040) );
  NOR2X1 U56021 ( .A(n53041), .B(n53040), .Y(n53043) );
  NOR2X1 U56022 ( .A(n18978), .B(n18977), .Y(n53042) );
  NAND2X1 U56023 ( .A(n53043), .B(n53042), .Y(u_decode_u_regfile_N820) );
  NOR2X1 U56024 ( .A(n43154), .B(n43277), .Y(n53045) );
  NOR2X1 U56025 ( .A(n43157), .B(n43384), .Y(n53044) );
  NOR2X1 U56026 ( .A(n53045), .B(n53044), .Y(n53047) );
  NOR2X1 U56027 ( .A(n20550), .B(n20549), .Y(n53046) );
  NAND2X1 U56028 ( .A(n53047), .B(n53046), .Y(u_decode_u_regfile_N524) );
  NOR2X1 U56029 ( .A(n44407), .B(n43155), .Y(n53049) );
  NOR2X1 U56030 ( .A(n44404), .B(n43158), .Y(n53048) );
  NOR2X1 U56031 ( .A(n53049), .B(n53048), .Y(n53051) );
  NOR2X1 U56032 ( .A(n22120), .B(n22119), .Y(n53050) );
  NAND2X1 U56033 ( .A(n53051), .B(n53050), .Y(u_decode_u_regfile_N228) );
  NOR2X1 U56034 ( .A(n44329), .B(n43155), .Y(n53053) );
  NOR2X1 U56035 ( .A(n44326), .B(n43158), .Y(n53052) );
  NOR2X1 U56036 ( .A(n53053), .B(n53052), .Y(n53055) );
  NOR2X1 U56037 ( .A(n23420), .B(n23419), .Y(n53054) );
  NAND2X1 U56038 ( .A(n53055), .B(n53054), .Y(u_decode_u_regfile_N1116) );
  NOR2X1 U56039 ( .A(n44584), .B(n43155), .Y(n53057) );
  NOR2X1 U56040 ( .A(n44581), .B(n43158), .Y(n53056) );
  NOR2X1 U56041 ( .A(n53057), .B(n53056), .Y(n53059) );
  NOR2X1 U56042 ( .A(n18586), .B(n18585), .Y(n53058) );
  NAND2X1 U56043 ( .A(n53059), .B(n53058), .Y(u_decode_u_regfile_N894) );
  NOR2X1 U56044 ( .A(n44431), .B(n43155), .Y(n53061) );
  NOR2X1 U56045 ( .A(n44428), .B(n43158), .Y(n53060) );
  NOR2X1 U56046 ( .A(n53061), .B(n53060), .Y(n53063) );
  NOR2X1 U56047 ( .A(n21728), .B(n21727), .Y(n53062) );
  NAND2X1 U56048 ( .A(n53063), .B(n53062), .Y(u_decode_u_regfile_N302) );
  NOR2X1 U56049 ( .A(n44515), .B(n43155), .Y(n53065) );
  NOR2X1 U56050 ( .A(n44512), .B(n43158), .Y(n53064) );
  NOR2X1 U56051 ( .A(n53065), .B(n53064), .Y(n53067) );
  NOR2X1 U56052 ( .A(n20158), .B(n20157), .Y(n53066) );
  NAND2X1 U56053 ( .A(n53067), .B(n53066), .Y(u_decode_u_regfile_N598) );
  NOR2X1 U56054 ( .A(n44353), .B(n43155), .Y(n53069) );
  NOR2X1 U56055 ( .A(n44350), .B(n43158), .Y(n53068) );
  NOR2X1 U56056 ( .A(n53069), .B(n53068), .Y(n53071) );
  NOR2X1 U56057 ( .A(n22980), .B(n22979), .Y(n53070) );
  NAND2X1 U56058 ( .A(n53071), .B(n53070), .Y(u_decode_u_regfile_N1190) );
  NOR2X1 U56059 ( .A(n44608), .B(n43155), .Y(n53073) );
  NOR2X1 U56060 ( .A(n44605), .B(n43158), .Y(n53072) );
  NOR2X1 U56061 ( .A(n53073), .B(n53072), .Y(n53075) );
  NOR2X1 U56062 ( .A(n24070), .B(n24069), .Y(n53074) );
  NAND2X1 U56063 ( .A(n53075), .B(n53074), .Y(u_decode_u_regfile_N1005) );
  NOR2X1 U56064 ( .A(n43154), .B(n43274), .Y(n53077) );
  NOR2X1 U56065 ( .A(n43157), .B(n43390), .Y(n53076) );
  NOR2X1 U56066 ( .A(n53077), .B(n53076), .Y(n53079) );
  NOR2X1 U56067 ( .A(n23100), .B(n23099), .Y(n53078) );
  NAND2X1 U56068 ( .A(n53079), .B(n53078), .Y(u_decode_u_regfile_N117) );
  NOR2X1 U56069 ( .A(n44461), .B(n43155), .Y(n53081) );
  NOR2X1 U56070 ( .A(n44458), .B(n43158), .Y(n53080) );
  NOR2X1 U56071 ( .A(n53081), .B(n53080), .Y(n53083) );
  NOR2X1 U56072 ( .A(n21138), .B(n21137), .Y(n53082) );
  NAND2X1 U56073 ( .A(n53083), .B(n53082), .Y(u_decode_u_regfile_N413) );
  NOR2X1 U56074 ( .A(n44551), .B(n43155), .Y(n53085) );
  NOR2X1 U56075 ( .A(n44548), .B(n43158), .Y(n53084) );
  NOR2X1 U56076 ( .A(n53085), .B(n53084), .Y(n53087) );
  NOR2X1 U56077 ( .A(n19568), .B(n19567), .Y(n53086) );
  NAND2X1 U56078 ( .A(n53087), .B(n53086), .Y(u_decode_u_regfile_N709) );
  NOR2X1 U56079 ( .A(n44566), .B(n43154), .Y(n53089) );
  NOR2X1 U56080 ( .A(n44563), .B(n43157), .Y(n53088) );
  NOR2X1 U56081 ( .A(n53089), .B(n53088), .Y(n53091) );
  NOR2X1 U56082 ( .A(n19174), .B(n19173), .Y(n53090) );
  NAND2X1 U56083 ( .A(n53091), .B(n53090), .Y(u_decode_u_regfile_N783) );
  NOR2X1 U56084 ( .A(n44317), .B(n43154), .Y(n53093) );
  NOR2X1 U56085 ( .A(n44314), .B(n43157), .Y(n53092) );
  NOR2X1 U56086 ( .A(n53093), .B(n53092), .Y(n53095) );
  NOR2X1 U56087 ( .A(n23640), .B(n23639), .Y(n53094) );
  NAND2X1 U56088 ( .A(n53095), .B(n53094), .Y(u_decode_u_regfile_N1079) );
  NOR2X1 U56089 ( .A(n44395), .B(n43154), .Y(n53097) );
  NOR2X1 U56090 ( .A(n44392), .B(n43157), .Y(n53096) );
  NOR2X1 U56091 ( .A(n53097), .B(n53096), .Y(n53099) );
  NOR2X1 U56092 ( .A(n22316), .B(n22315), .Y(n53098) );
  NAND2X1 U56093 ( .A(n53099), .B(n53098), .Y(u_decode_u_regfile_N191) );
  NOR2X1 U56094 ( .A(n44485), .B(n43155), .Y(n53101) );
  NOR2X1 U56095 ( .A(n44482), .B(n43157), .Y(n53100) );
  NOR2X1 U56096 ( .A(n53101), .B(n53100), .Y(n53103) );
  NOR2X1 U56097 ( .A(n20746), .B(n20745), .Y(n53102) );
  NAND2X1 U56098 ( .A(n53103), .B(n53102), .Y(u_decode_u_regfile_N487) );
  NOR2X1 U56099 ( .A(n44419), .B(n43154), .Y(n53105) );
  NOR2X1 U56100 ( .A(n44416), .B(n43157), .Y(n53104) );
  NOR2X1 U56101 ( .A(n53105), .B(n53104), .Y(n53107) );
  NOR2X1 U56102 ( .A(n21924), .B(n21923), .Y(n53106) );
  NAND2X1 U56103 ( .A(n53107), .B(n53106), .Y(u_decode_u_regfile_N265) );
  NOR2X1 U56104 ( .A(n44341), .B(n43154), .Y(n53109) );
  NOR2X1 U56105 ( .A(n44338), .B(n43157), .Y(n53108) );
  NOR2X1 U56106 ( .A(n53109), .B(n53108), .Y(n53111) );
  NOR2X1 U56107 ( .A(n23200), .B(n23199), .Y(n53110) );
  NAND2X1 U56108 ( .A(n53111), .B(n53110), .Y(u_decode_u_regfile_N1153) );
  NOR2X1 U56109 ( .A(n44503), .B(n43154), .Y(n53113) );
  NOR2X1 U56110 ( .A(n44500), .B(n43157), .Y(n53112) );
  NOR2X1 U56111 ( .A(n53113), .B(n53112), .Y(n53115) );
  NOR2X1 U56112 ( .A(n20354), .B(n20353), .Y(n53114) );
  NAND2X1 U56113 ( .A(n53115), .B(n53114), .Y(u_decode_u_regfile_N561) );
  NOR2X1 U56114 ( .A(n44578), .B(n43154), .Y(n53117) );
  NOR2X1 U56115 ( .A(n44575), .B(n43157), .Y(n53116) );
  NOR2X1 U56116 ( .A(n53117), .B(n53116), .Y(n53119) );
  NOR2X1 U56117 ( .A(n18782), .B(n18781), .Y(n53118) );
  NAND2X1 U56118 ( .A(n53119), .B(n53118), .Y(u_decode_u_regfile_N857) );
  NOR2X1 U56119 ( .A(n44527), .B(n43154), .Y(n53121) );
  NOR2X1 U56120 ( .A(n44524), .B(n43157), .Y(n53120) );
  NOR2X1 U56121 ( .A(n53121), .B(n53120), .Y(n53123) );
  NOR2X1 U56122 ( .A(n19962), .B(n19961), .Y(n53122) );
  NAND2X1 U56123 ( .A(n53123), .B(n53122), .Y(u_decode_u_regfile_N635) );
  NOR2X1 U56124 ( .A(n44593), .B(n43154), .Y(n53125) );
  NOR2X1 U56125 ( .A(n44590), .B(n43158), .Y(n53124) );
  NOR2X1 U56126 ( .A(n53125), .B(n53124), .Y(n53127) );
  NOR2X1 U56127 ( .A(n18392), .B(n18391), .Y(n53126) );
  NAND2X1 U56128 ( .A(n53127), .B(n53126), .Y(u_decode_u_regfile_N931) );
  NOR2X1 U56129 ( .A(n44365), .B(n43154), .Y(n53129) );
  NOR2X1 U56130 ( .A(n44362), .B(n43157), .Y(n53128) );
  NOR2X1 U56131 ( .A(n53129), .B(n53128), .Y(n53131) );
  NOR2X1 U56132 ( .A(n22766), .B(n22765), .Y(n53130) );
  NAND2X1 U56133 ( .A(n53131), .B(n53130), .Y(u_decode_u_regfile_N1227) );
  NOR2X1 U56134 ( .A(n44443), .B(n43155), .Y(n53133) );
  NOR2X1 U56135 ( .A(n44440), .B(n43158), .Y(n53132) );
  NOR2X1 U56136 ( .A(n53133), .B(n53132), .Y(n53135) );
  NOR2X1 U56137 ( .A(n21532), .B(n21531), .Y(n53134) );
  NAND2X1 U56138 ( .A(n53135), .B(n53134), .Y(u_decode_u_regfile_N339) );
  NOR2X1 U56139 ( .A(n16701), .B(n16702), .Y(n53137) );
  NOR2X1 U56140 ( .A(n16741), .B(n16742), .Y(n53136) );
  NAND2X1 U56141 ( .A(n53137), .B(n53136), .Y(u_exec_alu_p_w[18]) );
  NOR2X1 U56142 ( .A(n44538), .B(n43162), .Y(n53139) );
  NOR2X1 U56143 ( .A(n44536), .B(n37681), .Y(n53138) );
  NOR2X1 U56144 ( .A(n53139), .B(n53138), .Y(n53141) );
  NOR2X1 U56145 ( .A(n19759), .B(n19758), .Y(n53140) );
  NAND2X1 U56146 ( .A(n53141), .B(n53140), .Y(u_decode_u_regfile_N673) );
  NOR2X1 U56147 ( .A(n44602), .B(n43162), .Y(n53143) );
  NOR2X1 U56148 ( .A(n44599), .B(n37681), .Y(n53142) );
  NOR2X1 U56149 ( .A(n53143), .B(n53142), .Y(n53145) );
  NOR2X1 U56150 ( .A(n18181), .B(n18179), .Y(n53144) );
  NAND2X1 U56151 ( .A(n53145), .B(n53144), .Y(u_decode_u_regfile_N969) );
  NOR2X1 U56152 ( .A(n43160), .B(n43271), .Y(n53147) );
  NOR2X1 U56153 ( .A(n43163), .B(n43387), .Y(n53146) );
  NOR2X1 U56154 ( .A(n53147), .B(n53146), .Y(n53149) );
  NOR2X1 U56155 ( .A(n21329), .B(n21328), .Y(n53148) );
  NAND2X1 U56156 ( .A(n53149), .B(n53148), .Y(u_decode_u_regfile_N377) );
  NOR2X1 U56157 ( .A(n44473), .B(n43162), .Y(n53151) );
  NOR2X1 U56158 ( .A(n44470), .B(n37681), .Y(n53150) );
  NOR2X1 U56159 ( .A(n53151), .B(n53150), .Y(n53153) );
  NOR2X1 U56160 ( .A(n20936), .B(n20935), .Y(n53152) );
  NAND2X1 U56161 ( .A(n53153), .B(n53152), .Y(u_decode_u_regfile_N451) );
  NOR2X1 U56162 ( .A(n44560), .B(n43162), .Y(n53155) );
  NOR2X1 U56163 ( .A(n44557), .B(n37681), .Y(n53154) );
  NOR2X1 U56164 ( .A(n53155), .B(n53154), .Y(n53157) );
  NOR2X1 U56165 ( .A(n19364), .B(n19363), .Y(n53156) );
  NAND2X1 U56166 ( .A(n53157), .B(n53156), .Y(u_decode_u_regfile_N747) );
  NOR2X1 U56167 ( .A(n44383), .B(n43161), .Y(n53159) );
  NOR2X1 U56168 ( .A(n44380), .B(n43164), .Y(n53158) );
  NOR2X1 U56169 ( .A(n53159), .B(n53158), .Y(n53161) );
  NOR2X1 U56170 ( .A(n22506), .B(n22505), .Y(n53160) );
  NAND2X1 U56171 ( .A(n53161), .B(n53160), .Y(u_decode_u_regfile_N155) );
  NOR2X1 U56172 ( .A(n44305), .B(n43161), .Y(n53163) );
  NOR2X1 U56173 ( .A(n44302), .B(n43164), .Y(n53162) );
  NOR2X1 U56174 ( .A(n53163), .B(n53162), .Y(n53165) );
  NOR2X1 U56175 ( .A(n23848), .B(n23847), .Y(n53164) );
  NAND2X1 U56176 ( .A(n53165), .B(n53164), .Y(u_decode_u_regfile_N1043) );
  NOR2X1 U56177 ( .A(n44572), .B(n43161), .Y(n53167) );
  NOR2X1 U56178 ( .A(n44569), .B(n43164), .Y(n53166) );
  NOR2X1 U56179 ( .A(n53167), .B(n53166), .Y(n53169) );
  NOR2X1 U56180 ( .A(n18972), .B(n18971), .Y(n53168) );
  NAND2X1 U56181 ( .A(n53169), .B(n53168), .Y(u_decode_u_regfile_N821) );
  NOR2X1 U56182 ( .A(n43160), .B(n43277), .Y(n53171) );
  NOR2X1 U56183 ( .A(n43163), .B(n43384), .Y(n53170) );
  NOR2X1 U56184 ( .A(n53171), .B(n53170), .Y(n53173) );
  NOR2X1 U56185 ( .A(n20544), .B(n20543), .Y(n53172) );
  NAND2X1 U56186 ( .A(n53173), .B(n53172), .Y(u_decode_u_regfile_N525) );
  NOR2X1 U56187 ( .A(n44407), .B(n43161), .Y(n53175) );
  NOR2X1 U56188 ( .A(n44404), .B(n43164), .Y(n53174) );
  NOR2X1 U56189 ( .A(n53175), .B(n53174), .Y(n53177) );
  NOR2X1 U56190 ( .A(n22114), .B(n22113), .Y(n53176) );
  NAND2X1 U56191 ( .A(n53177), .B(n53176), .Y(u_decode_u_regfile_N229) );
  NOR2X1 U56192 ( .A(n44329), .B(n43161), .Y(n53179) );
  NOR2X1 U56193 ( .A(n44326), .B(n43164), .Y(n53178) );
  NOR2X1 U56194 ( .A(n53179), .B(n53178), .Y(n53181) );
  NOR2X1 U56195 ( .A(n23414), .B(n23413), .Y(n53180) );
  NAND2X1 U56196 ( .A(n53181), .B(n53180), .Y(u_decode_u_regfile_N1117) );
  NOR2X1 U56197 ( .A(n44584), .B(n43161), .Y(n53183) );
  NOR2X1 U56198 ( .A(n44581), .B(n43164), .Y(n53182) );
  NOR2X1 U56199 ( .A(n53183), .B(n53182), .Y(n53185) );
  NOR2X1 U56200 ( .A(n18580), .B(n18579), .Y(n53184) );
  NAND2X1 U56201 ( .A(n53185), .B(n53184), .Y(u_decode_u_regfile_N895) );
  NOR2X1 U56202 ( .A(n44431), .B(n43161), .Y(n53187) );
  NOR2X1 U56203 ( .A(n44428), .B(n43164), .Y(n53186) );
  NOR2X1 U56204 ( .A(n53187), .B(n53186), .Y(n53189) );
  NOR2X1 U56205 ( .A(n21722), .B(n21721), .Y(n53188) );
  NAND2X1 U56206 ( .A(n53189), .B(n53188), .Y(u_decode_u_regfile_N303) );
  NOR2X1 U56207 ( .A(n44515), .B(n43161), .Y(n53191) );
  NOR2X1 U56208 ( .A(n44512), .B(n43164), .Y(n53190) );
  NOR2X1 U56209 ( .A(n53191), .B(n53190), .Y(n53193) );
  NOR2X1 U56210 ( .A(n20152), .B(n20151), .Y(n53192) );
  NAND2X1 U56211 ( .A(n53193), .B(n53192), .Y(u_decode_u_regfile_N599) );
  NOR2X1 U56212 ( .A(n44353), .B(n43161), .Y(n53195) );
  NOR2X1 U56213 ( .A(n44350), .B(n43164), .Y(n53194) );
  NOR2X1 U56214 ( .A(n53195), .B(n53194), .Y(n53197) );
  NOR2X1 U56215 ( .A(n22974), .B(n22973), .Y(n53196) );
  NAND2X1 U56216 ( .A(n53197), .B(n53196), .Y(u_decode_u_regfile_N1191) );
  NOR2X1 U56217 ( .A(n44608), .B(n43161), .Y(n53199) );
  NOR2X1 U56218 ( .A(n44605), .B(n43164), .Y(n53198) );
  NOR2X1 U56219 ( .A(n53199), .B(n53198), .Y(n53201) );
  NOR2X1 U56220 ( .A(n24064), .B(n24063), .Y(n53200) );
  NAND2X1 U56221 ( .A(n53201), .B(n53200), .Y(u_decode_u_regfile_N1006) );
  NOR2X1 U56222 ( .A(n43160), .B(n43274), .Y(n53203) );
  NOR2X1 U56223 ( .A(n43163), .B(n43390), .Y(n53202) );
  NOR2X1 U56224 ( .A(n53203), .B(n53202), .Y(n53205) );
  NOR2X1 U56225 ( .A(n23052), .B(n23051), .Y(n53204) );
  NAND2X1 U56226 ( .A(n53205), .B(n53204), .Y(u_decode_u_regfile_N118) );
  NOR2X1 U56227 ( .A(n44461), .B(n43161), .Y(n53207) );
  NOR2X1 U56228 ( .A(n44458), .B(n43164), .Y(n53206) );
  NOR2X1 U56229 ( .A(n53207), .B(n53206), .Y(n53209) );
  NOR2X1 U56230 ( .A(n21132), .B(n21131), .Y(n53208) );
  NAND2X1 U56231 ( .A(n53209), .B(n53208), .Y(u_decode_u_regfile_N414) );
  NOR2X1 U56232 ( .A(n44551), .B(n43161), .Y(n53211) );
  NOR2X1 U56233 ( .A(n44548), .B(n43164), .Y(n53210) );
  NOR2X1 U56234 ( .A(n53211), .B(n53210), .Y(n53213) );
  NOR2X1 U56235 ( .A(n19562), .B(n19561), .Y(n53212) );
  NAND2X1 U56236 ( .A(n53213), .B(n53212), .Y(u_decode_u_regfile_N710) );
  NOR2X1 U56237 ( .A(n44566), .B(n43160), .Y(n53215) );
  NOR2X1 U56238 ( .A(n44563), .B(n43163), .Y(n53214) );
  NOR2X1 U56239 ( .A(n53215), .B(n53214), .Y(n53217) );
  NOR2X1 U56240 ( .A(n19168), .B(n19167), .Y(n53216) );
  NAND2X1 U56241 ( .A(n53217), .B(n53216), .Y(u_decode_u_regfile_N784) );
  NOR2X1 U56242 ( .A(n44317), .B(n43160), .Y(n53219) );
  NOR2X1 U56243 ( .A(n44314), .B(n43163), .Y(n53218) );
  NOR2X1 U56244 ( .A(n53219), .B(n53218), .Y(n53221) );
  NOR2X1 U56245 ( .A(n23628), .B(n23627), .Y(n53220) );
  NAND2X1 U56246 ( .A(n53221), .B(n53220), .Y(u_decode_u_regfile_N1080) );
  NOR2X1 U56247 ( .A(n44395), .B(n43160), .Y(n53223) );
  NOR2X1 U56248 ( .A(n44392), .B(n43163), .Y(n53222) );
  NOR2X1 U56249 ( .A(n53223), .B(n53222), .Y(n53225) );
  NOR2X1 U56250 ( .A(n22310), .B(n22309), .Y(n53224) );
  NAND2X1 U56251 ( .A(n53225), .B(n53224), .Y(u_decode_u_regfile_N192) );
  NOR2X1 U56252 ( .A(n44485), .B(n43161), .Y(n53227) );
  NOR2X1 U56253 ( .A(n44482), .B(n43163), .Y(n53226) );
  NOR2X1 U56254 ( .A(n53227), .B(n53226), .Y(n53229) );
  NOR2X1 U56255 ( .A(n20740), .B(n20739), .Y(n53228) );
  NAND2X1 U56256 ( .A(n53229), .B(n53228), .Y(u_decode_u_regfile_N488) );
  NOR2X1 U56257 ( .A(n44419), .B(n43160), .Y(n53231) );
  NOR2X1 U56258 ( .A(n44416), .B(n43163), .Y(n53230) );
  NOR2X1 U56259 ( .A(n53231), .B(n53230), .Y(n53233) );
  NOR2X1 U56260 ( .A(n21918), .B(n21917), .Y(n53232) );
  NAND2X1 U56261 ( .A(n53233), .B(n53232), .Y(u_decode_u_regfile_N266) );
  NOR2X1 U56262 ( .A(n44341), .B(n43160), .Y(n53235) );
  NOR2X1 U56263 ( .A(n44338), .B(n43163), .Y(n53234) );
  NOR2X1 U56264 ( .A(n53235), .B(n53234), .Y(n53237) );
  NOR2X1 U56265 ( .A(n23194), .B(n23193), .Y(n53236) );
  NAND2X1 U56266 ( .A(n53237), .B(n53236), .Y(u_decode_u_regfile_N1154) );
  NOR2X1 U56267 ( .A(n44503), .B(n43160), .Y(n53239) );
  NOR2X1 U56268 ( .A(n44500), .B(n43163), .Y(n53238) );
  NOR2X1 U56269 ( .A(n53239), .B(n53238), .Y(n53241) );
  NOR2X1 U56270 ( .A(n20348), .B(n20347), .Y(n53240) );
  NAND2X1 U56271 ( .A(n53241), .B(n53240), .Y(u_decode_u_regfile_N562) );
  NOR2X1 U56272 ( .A(n44578), .B(n43160), .Y(n53243) );
  NOR2X1 U56273 ( .A(n44575), .B(n43163), .Y(n53242) );
  NOR2X1 U56274 ( .A(n53243), .B(n53242), .Y(n53245) );
  NOR2X1 U56275 ( .A(n18776), .B(n18775), .Y(n53244) );
  NAND2X1 U56276 ( .A(n53245), .B(n53244), .Y(u_decode_u_regfile_N858) );
  NOR2X1 U56277 ( .A(n44527), .B(n43160), .Y(n53247) );
  NOR2X1 U56278 ( .A(n44524), .B(n43163), .Y(n53246) );
  NOR2X1 U56279 ( .A(n53247), .B(n53246), .Y(n53249) );
  NOR2X1 U56280 ( .A(n19956), .B(n19955), .Y(n53248) );
  NAND2X1 U56281 ( .A(n53249), .B(n53248), .Y(u_decode_u_regfile_N636) );
  NOR2X1 U56282 ( .A(n44593), .B(n43160), .Y(n53251) );
  NOR2X1 U56283 ( .A(n44590), .B(n43164), .Y(n53250) );
  NOR2X1 U56284 ( .A(n53251), .B(n53250), .Y(n53253) );
  NOR2X1 U56285 ( .A(n18386), .B(n18385), .Y(n53252) );
  NAND2X1 U56286 ( .A(n53253), .B(n53252), .Y(u_decode_u_regfile_N932) );
  NOR2X1 U56287 ( .A(n44365), .B(n43160), .Y(n53255) );
  NOR2X1 U56288 ( .A(n44362), .B(n43163), .Y(n53254) );
  NOR2X1 U56289 ( .A(n53255), .B(n53254), .Y(n53257) );
  NOR2X1 U56290 ( .A(n22760), .B(n22759), .Y(n53256) );
  NAND2X1 U56291 ( .A(n53257), .B(n53256), .Y(u_decode_u_regfile_N1228) );
  NOR2X1 U56292 ( .A(n44443), .B(n43161), .Y(n53259) );
  NOR2X1 U56293 ( .A(n44440), .B(n43164), .Y(n53258) );
  NOR2X1 U56294 ( .A(n53259), .B(n53258), .Y(n53261) );
  NOR2X1 U56295 ( .A(n21526), .B(n21525), .Y(n53260) );
  NAND2X1 U56296 ( .A(n53261), .B(n53260), .Y(u_decode_u_regfile_N340) );
  NOR2X1 U56297 ( .A(n16645), .B(n16646), .Y(n53263) );
  NOR2X1 U56298 ( .A(n16687), .B(n16688), .Y(n53262) );
  NAND2X1 U56299 ( .A(n53263), .B(n53262), .Y(u_exec_alu_p_w[19]) );
  NOR2X1 U56300 ( .A(n44538), .B(n43168), .Y(n53265) );
  NOR2X1 U56301 ( .A(n44536), .B(n43170), .Y(n53264) );
  NOR2X1 U56302 ( .A(n53265), .B(n53264), .Y(n53267) );
  NOR2X1 U56303 ( .A(n19753), .B(n19752), .Y(n53266) );
  NAND2X1 U56304 ( .A(n53267), .B(n53266), .Y(u_decode_u_regfile_N674) );
  NOR2X1 U56305 ( .A(n44602), .B(n43168), .Y(n53269) );
  NOR2X1 U56306 ( .A(n44599), .B(n43170), .Y(n53268) );
  NOR2X1 U56307 ( .A(n53269), .B(n53268), .Y(n53271) );
  NOR2X1 U56308 ( .A(n18174), .B(n18172), .Y(n53270) );
  NAND2X1 U56309 ( .A(n53271), .B(n53270), .Y(u_decode_u_regfile_N970) );
  NOR2X1 U56310 ( .A(n43166), .B(n43271), .Y(n53273) );
  NOR2X1 U56311 ( .A(n43169), .B(n43387), .Y(n53272) );
  NOR2X1 U56312 ( .A(n53273), .B(n53272), .Y(n53275) );
  NOR2X1 U56313 ( .A(n21323), .B(n21322), .Y(n53274) );
  NAND2X1 U56314 ( .A(n53275), .B(n53274), .Y(u_decode_u_regfile_N378) );
  NOR2X1 U56315 ( .A(n44473), .B(n43168), .Y(n53277) );
  NOR2X1 U56316 ( .A(n44470), .B(n43170), .Y(n53276) );
  NOR2X1 U56317 ( .A(n53277), .B(n53276), .Y(n53279) );
  NOR2X1 U56318 ( .A(n20930), .B(n20929), .Y(n53278) );
  NAND2X1 U56319 ( .A(n53279), .B(n53278), .Y(u_decode_u_regfile_N452) );
  NOR2X1 U56320 ( .A(n44560), .B(n43168), .Y(n53281) );
  NOR2X1 U56321 ( .A(n44557), .B(n43170), .Y(n53280) );
  NOR2X1 U56322 ( .A(n53281), .B(n53280), .Y(n53283) );
  NOR2X1 U56323 ( .A(n19358), .B(n19357), .Y(n53282) );
  NAND2X1 U56324 ( .A(n53283), .B(n53282), .Y(u_decode_u_regfile_N748) );
  NOR2X1 U56325 ( .A(n44383), .B(n43167), .Y(n53285) );
  NOR2X1 U56326 ( .A(n44380), .B(n37593), .Y(n53284) );
  NOR2X1 U56327 ( .A(n53285), .B(n53284), .Y(n53287) );
  NOR2X1 U56328 ( .A(n22500), .B(n22499), .Y(n53286) );
  NAND2X1 U56329 ( .A(n53287), .B(n53286), .Y(u_decode_u_regfile_N156) );
  NOR2X1 U56330 ( .A(n44305), .B(n43167), .Y(n53289) );
  NOR2X1 U56331 ( .A(n44302), .B(n37593), .Y(n53288) );
  NOR2X1 U56332 ( .A(n53289), .B(n53288), .Y(n53291) );
  NOR2X1 U56333 ( .A(n23842), .B(n23841), .Y(n53290) );
  NAND2X1 U56334 ( .A(n53291), .B(n53290), .Y(u_decode_u_regfile_N1044) );
  NOR2X1 U56335 ( .A(n44572), .B(n43167), .Y(n53293) );
  NOR2X1 U56336 ( .A(n44569), .B(n37593), .Y(n53292) );
  NOR2X1 U56337 ( .A(n53293), .B(n53292), .Y(n53295) );
  NOR2X1 U56338 ( .A(n18966), .B(n18965), .Y(n53294) );
  NAND2X1 U56339 ( .A(n53295), .B(n53294), .Y(u_decode_u_regfile_N822) );
  NOR2X1 U56340 ( .A(n43166), .B(n43277), .Y(n53297) );
  NOR2X1 U56341 ( .A(n43169), .B(n43384), .Y(n53296) );
  NOR2X1 U56342 ( .A(n53297), .B(n53296), .Y(n53299) );
  NOR2X1 U56343 ( .A(n20538), .B(n20537), .Y(n53298) );
  NAND2X1 U56344 ( .A(n53299), .B(n53298), .Y(u_decode_u_regfile_N526) );
  NOR2X1 U56345 ( .A(n44407), .B(n43167), .Y(n53301) );
  NOR2X1 U56346 ( .A(n44404), .B(n37593), .Y(n53300) );
  NOR2X1 U56347 ( .A(n53301), .B(n53300), .Y(n53303) );
  NOR2X1 U56348 ( .A(n22108), .B(n22107), .Y(n53302) );
  NAND2X1 U56349 ( .A(n53303), .B(n53302), .Y(u_decode_u_regfile_N230) );
  NOR2X1 U56350 ( .A(n44329), .B(n43167), .Y(n53305) );
  NOR2X1 U56351 ( .A(n44326), .B(n37593), .Y(n53304) );
  NOR2X1 U56352 ( .A(n53305), .B(n53304), .Y(n53307) );
  NOR2X1 U56353 ( .A(n23408), .B(n23407), .Y(n53306) );
  NAND2X1 U56354 ( .A(n53307), .B(n53306), .Y(u_decode_u_regfile_N1118) );
  NOR2X1 U56355 ( .A(n44584), .B(n43167), .Y(n53309) );
  NOR2X1 U56356 ( .A(n44581), .B(n37593), .Y(n53308) );
  NOR2X1 U56357 ( .A(n53309), .B(n53308), .Y(n53311) );
  NOR2X1 U56358 ( .A(n18574), .B(n18573), .Y(n53310) );
  NAND2X1 U56359 ( .A(n53311), .B(n53310), .Y(u_decode_u_regfile_N896) );
  NOR2X1 U56360 ( .A(n44431), .B(n43167), .Y(n53313) );
  NOR2X1 U56361 ( .A(n44428), .B(n37593), .Y(n53312) );
  NOR2X1 U56362 ( .A(n53313), .B(n53312), .Y(n53315) );
  NOR2X1 U56363 ( .A(n21716), .B(n21715), .Y(n53314) );
  NAND2X1 U56364 ( .A(n53315), .B(n53314), .Y(u_decode_u_regfile_N304) );
  NOR2X1 U56365 ( .A(n44515), .B(n43167), .Y(n53317) );
  NOR2X1 U56366 ( .A(n44512), .B(n37593), .Y(n53316) );
  NOR2X1 U56367 ( .A(n53317), .B(n53316), .Y(n53319) );
  NOR2X1 U56368 ( .A(n20146), .B(n20145), .Y(n53318) );
  NAND2X1 U56369 ( .A(n53319), .B(n53318), .Y(u_decode_u_regfile_N600) );
  NOR2X1 U56370 ( .A(n44353), .B(n43167), .Y(n53321) );
  NOR2X1 U56371 ( .A(n44350), .B(n37593), .Y(n53320) );
  NOR2X1 U56372 ( .A(n53321), .B(n53320), .Y(n53323) );
  NOR2X1 U56373 ( .A(n22968), .B(n22967), .Y(n53322) );
  NAND2X1 U56374 ( .A(n53323), .B(n53322), .Y(u_decode_u_regfile_N1192) );
  NOR2X1 U56375 ( .A(n44608), .B(n43167), .Y(n53325) );
  NOR2X1 U56376 ( .A(n44605), .B(n37593), .Y(n53324) );
  NOR2X1 U56377 ( .A(n53325), .B(n53324), .Y(n53327) );
  NOR2X1 U56378 ( .A(n24058), .B(n24057), .Y(n53326) );
  NAND2X1 U56379 ( .A(n53327), .B(n53326), .Y(u_decode_u_regfile_N1007) );
  NOR2X1 U56380 ( .A(n43166), .B(n43274), .Y(n53329) );
  NOR2X1 U56381 ( .A(n43169), .B(n43390), .Y(n53328) );
  NOR2X1 U56382 ( .A(n53329), .B(n53328), .Y(n53331) );
  NOR2X1 U56383 ( .A(n22986), .B(n22985), .Y(n53330) );
  NAND2X1 U56384 ( .A(n53331), .B(n53330), .Y(u_decode_u_regfile_N119) );
  NOR2X1 U56385 ( .A(n44461), .B(n43167), .Y(n53333) );
  NOR2X1 U56386 ( .A(n44458), .B(n37593), .Y(n53332) );
  NOR2X1 U56387 ( .A(n53333), .B(n53332), .Y(n53335) );
  NOR2X1 U56388 ( .A(n21126), .B(n21125), .Y(n53334) );
  NAND2X1 U56389 ( .A(n53335), .B(n53334), .Y(u_decode_u_regfile_N415) );
  NOR2X1 U56390 ( .A(n44551), .B(n43167), .Y(n53337) );
  NOR2X1 U56391 ( .A(n44548), .B(n37593), .Y(n53336) );
  NOR2X1 U56392 ( .A(n53337), .B(n53336), .Y(n53339) );
  NOR2X1 U56393 ( .A(n19556), .B(n19555), .Y(n53338) );
  NAND2X1 U56394 ( .A(n53339), .B(n53338), .Y(u_decode_u_regfile_N711) );
  NOR2X1 U56395 ( .A(n44566), .B(n43166), .Y(n53341) );
  NOR2X1 U56396 ( .A(n44563), .B(n43169), .Y(n53340) );
  NOR2X1 U56397 ( .A(n53341), .B(n53340), .Y(n53343) );
  NOR2X1 U56398 ( .A(n19162), .B(n19161), .Y(n53342) );
  NAND2X1 U56399 ( .A(n53343), .B(n53342), .Y(u_decode_u_regfile_N785) );
  NOR2X1 U56400 ( .A(n44317), .B(n43166), .Y(n53345) );
  NOR2X1 U56401 ( .A(n44314), .B(n43169), .Y(n53344) );
  NOR2X1 U56402 ( .A(n53345), .B(n53344), .Y(n53347) );
  NOR2X1 U56403 ( .A(n23622), .B(n23621), .Y(n53346) );
  NAND2X1 U56404 ( .A(n53347), .B(n53346), .Y(u_decode_u_regfile_N1081) );
  NOR2X1 U56405 ( .A(n44395), .B(n43166), .Y(n53349) );
  NOR2X1 U56406 ( .A(n44392), .B(n43169), .Y(n53348) );
  NOR2X1 U56407 ( .A(n53349), .B(n53348), .Y(n53351) );
  NOR2X1 U56408 ( .A(n22304), .B(n22303), .Y(n53350) );
  NAND2X1 U56409 ( .A(n53351), .B(n53350), .Y(u_decode_u_regfile_N193) );
  NOR2X1 U56410 ( .A(n44485), .B(n43166), .Y(n53353) );
  NOR2X1 U56411 ( .A(n44482), .B(n37593), .Y(n53352) );
  NOR2X1 U56412 ( .A(n53353), .B(n53352), .Y(n53355) );
  NOR2X1 U56413 ( .A(n20734), .B(n20733), .Y(n53354) );
  NAND2X1 U56414 ( .A(n53355), .B(n53354), .Y(u_decode_u_regfile_N489) );
  NOR2X1 U56415 ( .A(n44419), .B(n43166), .Y(n53357) );
  NOR2X1 U56416 ( .A(n44416), .B(n43169), .Y(n53356) );
  NOR2X1 U56417 ( .A(n53357), .B(n53356), .Y(n53359) );
  NOR2X1 U56418 ( .A(n21912), .B(n21911), .Y(n53358) );
  NAND2X1 U56419 ( .A(n53359), .B(n53358), .Y(u_decode_u_regfile_N267) );
  NOR2X1 U56420 ( .A(n44341), .B(n43166), .Y(n53361) );
  NOR2X1 U56421 ( .A(n44338), .B(n43169), .Y(n53360) );
  NOR2X1 U56422 ( .A(n53361), .B(n53360), .Y(n53363) );
  NOR2X1 U56423 ( .A(n23188), .B(n23187), .Y(n53362) );
  NAND2X1 U56424 ( .A(n53363), .B(n53362), .Y(u_decode_u_regfile_N1155) );
  NOR2X1 U56425 ( .A(n44503), .B(n43166), .Y(n53365) );
  NOR2X1 U56426 ( .A(n44500), .B(n43169), .Y(n53364) );
  NOR2X1 U56427 ( .A(n53365), .B(n53364), .Y(n53367) );
  NOR2X1 U56428 ( .A(n20342), .B(n20341), .Y(n53366) );
  NAND2X1 U56429 ( .A(n53367), .B(n53366), .Y(u_decode_u_regfile_N563) );
  NOR2X1 U56430 ( .A(n44578), .B(n43166), .Y(n53369) );
  NOR2X1 U56431 ( .A(n44575), .B(n43169), .Y(n53368) );
  NOR2X1 U56432 ( .A(n53369), .B(n53368), .Y(n53371) );
  NOR2X1 U56433 ( .A(n18770), .B(n18769), .Y(n53370) );
  NAND2X1 U56434 ( .A(n53371), .B(n53370), .Y(u_decode_u_regfile_N859) );
  NOR2X1 U56435 ( .A(n44527), .B(n43166), .Y(n53373) );
  NOR2X1 U56436 ( .A(n44524), .B(n43169), .Y(n53372) );
  NOR2X1 U56437 ( .A(n53373), .B(n53372), .Y(n53375) );
  NOR2X1 U56438 ( .A(n19950), .B(n19949), .Y(n53374) );
  NAND2X1 U56439 ( .A(n53375), .B(n53374), .Y(u_decode_u_regfile_N637) );
  NOR2X1 U56440 ( .A(n44593), .B(n43167), .Y(n53377) );
  NOR2X1 U56441 ( .A(n44590), .B(n43169), .Y(n53376) );
  NOR2X1 U56442 ( .A(n53377), .B(n53376), .Y(n53379) );
  NOR2X1 U56443 ( .A(n18380), .B(n18379), .Y(n53378) );
  NAND2X1 U56444 ( .A(n53379), .B(n53378), .Y(u_decode_u_regfile_N933) );
  NOR2X1 U56445 ( .A(n44365), .B(n43166), .Y(n53381) );
  NOR2X1 U56446 ( .A(n44362), .B(n43169), .Y(n53380) );
  NOR2X1 U56447 ( .A(n53381), .B(n53380), .Y(n53383) );
  NOR2X1 U56448 ( .A(n22754), .B(n22753), .Y(n53382) );
  NAND2X1 U56449 ( .A(n53383), .B(n53382), .Y(u_decode_u_regfile_N1229) );
  NOR2X1 U56450 ( .A(n44443), .B(n43167), .Y(n53385) );
  NOR2X1 U56451 ( .A(n44440), .B(n37593), .Y(n53384) );
  NOR2X1 U56452 ( .A(n53385), .B(n53384), .Y(n53387) );
  NOR2X1 U56453 ( .A(n21520), .B(n21519), .Y(n53386) );
  NAND2X1 U56454 ( .A(n53387), .B(n53386), .Y(u_decode_u_regfile_N341) );
  NOR2X1 U56455 ( .A(n16525), .B(n16526), .Y(n53389) );
  NOR2X1 U56456 ( .A(n16567), .B(n16568), .Y(n53388) );
  NAND2X1 U56457 ( .A(n53389), .B(n53388), .Y(u_exec_alu_p_w[20]) );
  NOR2X1 U56458 ( .A(n44538), .B(n43173), .Y(n53391) );
  NOR2X1 U56459 ( .A(n44536), .B(n43175), .Y(n53390) );
  NOR2X1 U56460 ( .A(n53391), .B(n53390), .Y(n53393) );
  NOR2X1 U56461 ( .A(n19747), .B(n19746), .Y(n53392) );
  NAND2X1 U56462 ( .A(n53393), .B(n53392), .Y(u_decode_u_regfile_N675) );
  NOR2X1 U56463 ( .A(n44602), .B(n43173), .Y(n53395) );
  NOR2X1 U56464 ( .A(n44599), .B(n43175), .Y(n53394) );
  NOR2X1 U56465 ( .A(n53395), .B(n53394), .Y(n53397) );
  NOR2X1 U56466 ( .A(n18167), .B(n18165), .Y(n53396) );
  NAND2X1 U56467 ( .A(n53397), .B(n53396), .Y(u_decode_u_regfile_N971) );
  NOR2X1 U56468 ( .A(n43171), .B(n43271), .Y(n53399) );
  NOR2X1 U56469 ( .A(n43174), .B(n43386), .Y(n53398) );
  NOR2X1 U56470 ( .A(n53399), .B(n53398), .Y(n53401) );
  NOR2X1 U56471 ( .A(n21317), .B(n21316), .Y(n53400) );
  NAND2X1 U56472 ( .A(n53401), .B(n53400), .Y(u_decode_u_regfile_N379) );
  NOR2X1 U56473 ( .A(n44473), .B(n43173), .Y(n53403) );
  NOR2X1 U56474 ( .A(n44470), .B(n43175), .Y(n53402) );
  NOR2X1 U56475 ( .A(n53403), .B(n53402), .Y(n53405) );
  NOR2X1 U56476 ( .A(n20924), .B(n20923), .Y(n53404) );
  NAND2X1 U56477 ( .A(n53405), .B(n53404), .Y(u_decode_u_regfile_N453) );
  NOR2X1 U56478 ( .A(n44560), .B(n43173), .Y(n53407) );
  NOR2X1 U56479 ( .A(n44557), .B(n43175), .Y(n53406) );
  NOR2X1 U56480 ( .A(n53407), .B(n53406), .Y(n53409) );
  NOR2X1 U56481 ( .A(n19352), .B(n19351), .Y(n53408) );
  NAND2X1 U56482 ( .A(n53409), .B(n53408), .Y(u_decode_u_regfile_N749) );
  NOR2X1 U56483 ( .A(n44383), .B(n43172), .Y(n53411) );
  NOR2X1 U56484 ( .A(n44380), .B(n37594), .Y(n53410) );
  NOR2X1 U56485 ( .A(n53411), .B(n53410), .Y(n53413) );
  NOR2X1 U56486 ( .A(n22494), .B(n22493), .Y(n53412) );
  NAND2X1 U56487 ( .A(n53413), .B(n53412), .Y(u_decode_u_regfile_N157) );
  NOR2X1 U56488 ( .A(n44305), .B(n43172), .Y(n53415) );
  NOR2X1 U56489 ( .A(n44302), .B(n37594), .Y(n53414) );
  NOR2X1 U56490 ( .A(n53415), .B(n53414), .Y(n53417) );
  NOR2X1 U56491 ( .A(n23836), .B(n23835), .Y(n53416) );
  NAND2X1 U56492 ( .A(n53417), .B(n53416), .Y(u_decode_u_regfile_N1045) );
  NOR2X1 U56493 ( .A(n44572), .B(n43172), .Y(n53419) );
  NOR2X1 U56494 ( .A(n44569), .B(n37594), .Y(n53418) );
  NOR2X1 U56495 ( .A(n53419), .B(n53418), .Y(n53421) );
  NOR2X1 U56496 ( .A(n18960), .B(n18959), .Y(n53420) );
  NAND2X1 U56497 ( .A(n53421), .B(n53420), .Y(u_decode_u_regfile_N823) );
  NOR2X1 U56498 ( .A(n43171), .B(n43277), .Y(n53423) );
  NOR2X1 U56499 ( .A(n43174), .B(n43383), .Y(n53422) );
  NOR2X1 U56500 ( .A(n53423), .B(n53422), .Y(n53425) );
  NOR2X1 U56501 ( .A(n20532), .B(n20531), .Y(n53424) );
  NAND2X1 U56502 ( .A(n53425), .B(n53424), .Y(u_decode_u_regfile_N527) );
  NOR2X1 U56503 ( .A(n44407), .B(n43172), .Y(n53427) );
  NOR2X1 U56504 ( .A(n44404), .B(n37594), .Y(n53426) );
  NOR2X1 U56505 ( .A(n53427), .B(n53426), .Y(n53429) );
  NOR2X1 U56506 ( .A(n22102), .B(n22101), .Y(n53428) );
  NAND2X1 U56507 ( .A(n53429), .B(n53428), .Y(u_decode_u_regfile_N231) );
  NOR2X1 U56508 ( .A(n44329), .B(n43172), .Y(n53431) );
  NOR2X1 U56509 ( .A(n44326), .B(n37594), .Y(n53430) );
  NOR2X1 U56510 ( .A(n53431), .B(n53430), .Y(n53433) );
  NOR2X1 U56511 ( .A(n23402), .B(n23401), .Y(n53432) );
  NAND2X1 U56512 ( .A(n53433), .B(n53432), .Y(u_decode_u_regfile_N1119) );
  NOR2X1 U56513 ( .A(n44584), .B(n43172), .Y(n53435) );
  NOR2X1 U56514 ( .A(n44581), .B(n37594), .Y(n53434) );
  NOR2X1 U56515 ( .A(n53435), .B(n53434), .Y(n53437) );
  NOR2X1 U56516 ( .A(n18568), .B(n18567), .Y(n53436) );
  NAND2X1 U56517 ( .A(n53437), .B(n53436), .Y(u_decode_u_regfile_N897) );
  NOR2X1 U56518 ( .A(n44431), .B(n43172), .Y(n53439) );
  NOR2X1 U56519 ( .A(n44428), .B(n37594), .Y(n53438) );
  NOR2X1 U56520 ( .A(n53439), .B(n53438), .Y(n53441) );
  NOR2X1 U56521 ( .A(n21710), .B(n21709), .Y(n53440) );
  NAND2X1 U56522 ( .A(n53441), .B(n53440), .Y(u_decode_u_regfile_N305) );
  NOR2X1 U56523 ( .A(n44515), .B(n43172), .Y(n53443) );
  NOR2X1 U56524 ( .A(n44512), .B(n37594), .Y(n53442) );
  NOR2X1 U56525 ( .A(n53443), .B(n53442), .Y(n53445) );
  NOR2X1 U56526 ( .A(n20140), .B(n20139), .Y(n53444) );
  NAND2X1 U56527 ( .A(n53445), .B(n53444), .Y(u_decode_u_regfile_N601) );
  NOR2X1 U56528 ( .A(n44353), .B(n43172), .Y(n53447) );
  NOR2X1 U56529 ( .A(n44350), .B(n37594), .Y(n53446) );
  NOR2X1 U56530 ( .A(n53447), .B(n53446), .Y(n53449) );
  NOR2X1 U56531 ( .A(n22962), .B(n22961), .Y(n53448) );
  NAND2X1 U56532 ( .A(n53449), .B(n53448), .Y(u_decode_u_regfile_N1193) );
  NOR2X1 U56533 ( .A(n44608), .B(n43172), .Y(n53451) );
  NOR2X1 U56534 ( .A(n44605), .B(n37594), .Y(n53450) );
  NOR2X1 U56535 ( .A(n53451), .B(n53450), .Y(n53453) );
  NOR2X1 U56536 ( .A(n24052), .B(n24051), .Y(n53452) );
  NAND2X1 U56537 ( .A(n53453), .B(n53452), .Y(u_decode_u_regfile_N1008) );
  NOR2X1 U56538 ( .A(n43171), .B(n43274), .Y(n53455) );
  NOR2X1 U56539 ( .A(n43174), .B(n43389), .Y(n53454) );
  NOR2X1 U56540 ( .A(n53455), .B(n53454), .Y(n53457) );
  NOR2X1 U56541 ( .A(n22920), .B(n22919), .Y(n53456) );
  NAND2X1 U56542 ( .A(n53457), .B(n53456), .Y(u_decode_u_regfile_N120) );
  NOR2X1 U56543 ( .A(n44461), .B(n43172), .Y(n53459) );
  NOR2X1 U56544 ( .A(n44458), .B(n37594), .Y(n53458) );
  NOR2X1 U56545 ( .A(n53459), .B(n53458), .Y(n53461) );
  NOR2X1 U56546 ( .A(n21120), .B(n21119), .Y(n53460) );
  NAND2X1 U56547 ( .A(n53461), .B(n53460), .Y(u_decode_u_regfile_N416) );
  NOR2X1 U56548 ( .A(n44551), .B(n43172), .Y(n53463) );
  NOR2X1 U56549 ( .A(n44548), .B(n37594), .Y(n53462) );
  NOR2X1 U56550 ( .A(n53463), .B(n53462), .Y(n53465) );
  NOR2X1 U56551 ( .A(n19550), .B(n19549), .Y(n53464) );
  NAND2X1 U56552 ( .A(n53465), .B(n53464), .Y(u_decode_u_regfile_N712) );
  NOR2X1 U56553 ( .A(n44566), .B(n43171), .Y(n53467) );
  NOR2X1 U56554 ( .A(n44563), .B(n43174), .Y(n53466) );
  NOR2X1 U56555 ( .A(n53467), .B(n53466), .Y(n53469) );
  NOR2X1 U56556 ( .A(n19156), .B(n19155), .Y(n53468) );
  NAND2X1 U56557 ( .A(n53469), .B(n53468), .Y(u_decode_u_regfile_N786) );
  NOR2X1 U56558 ( .A(n44317), .B(n43171), .Y(n53471) );
  NOR2X1 U56559 ( .A(n44314), .B(n43174), .Y(n53470) );
  NOR2X1 U56560 ( .A(n53471), .B(n53470), .Y(n53473) );
  NOR2X1 U56561 ( .A(n23616), .B(n23615), .Y(n53472) );
  NAND2X1 U56562 ( .A(n53473), .B(n53472), .Y(u_decode_u_regfile_N1082) );
  NOR2X1 U56563 ( .A(n44395), .B(n43171), .Y(n53475) );
  NOR2X1 U56564 ( .A(n44392), .B(n43174), .Y(n53474) );
  NOR2X1 U56565 ( .A(n53475), .B(n53474), .Y(n53477) );
  NOR2X1 U56566 ( .A(n22298), .B(n22297), .Y(n53476) );
  NAND2X1 U56567 ( .A(n53477), .B(n53476), .Y(u_decode_u_regfile_N194) );
  NOR2X1 U56568 ( .A(n44485), .B(n43172), .Y(n53479) );
  NOR2X1 U56569 ( .A(n44482), .B(n37594), .Y(n53478) );
  NOR2X1 U56570 ( .A(n53479), .B(n53478), .Y(n53481) );
  NOR2X1 U56571 ( .A(n20728), .B(n20727), .Y(n53480) );
  NAND2X1 U56572 ( .A(n53481), .B(n53480), .Y(u_decode_u_regfile_N490) );
  NOR2X1 U56573 ( .A(n44419), .B(n43171), .Y(n53483) );
  NOR2X1 U56574 ( .A(n44416), .B(n43174), .Y(n53482) );
  NOR2X1 U56575 ( .A(n53483), .B(n53482), .Y(n53485) );
  NOR2X1 U56576 ( .A(n21906), .B(n21905), .Y(n53484) );
  NAND2X1 U56577 ( .A(n53485), .B(n53484), .Y(u_decode_u_regfile_N268) );
  NOR2X1 U56578 ( .A(n44341), .B(n43171), .Y(n53487) );
  NOR2X1 U56579 ( .A(n44338), .B(n43174), .Y(n53486) );
  NOR2X1 U56580 ( .A(n53487), .B(n53486), .Y(n53489) );
  NOR2X1 U56581 ( .A(n23182), .B(n23181), .Y(n53488) );
  NAND2X1 U56582 ( .A(n53489), .B(n53488), .Y(u_decode_u_regfile_N1156) );
  NOR2X1 U56583 ( .A(n44503), .B(n43171), .Y(n53491) );
  NOR2X1 U56584 ( .A(n44500), .B(n43174), .Y(n53490) );
  NOR2X1 U56585 ( .A(n53491), .B(n53490), .Y(n53493) );
  NOR2X1 U56586 ( .A(n20336), .B(n20335), .Y(n53492) );
  NAND2X1 U56587 ( .A(n53493), .B(n53492), .Y(u_decode_u_regfile_N564) );
  NOR2X1 U56588 ( .A(n44578), .B(n43171), .Y(n53495) );
  NOR2X1 U56589 ( .A(n44575), .B(n43174), .Y(n53494) );
  NOR2X1 U56590 ( .A(n53495), .B(n53494), .Y(n53497) );
  NOR2X1 U56591 ( .A(n18764), .B(n18763), .Y(n53496) );
  NAND2X1 U56592 ( .A(n53497), .B(n53496), .Y(u_decode_u_regfile_N860) );
  NOR2X1 U56593 ( .A(n44527), .B(n43171), .Y(n53499) );
  NOR2X1 U56594 ( .A(n44524), .B(n43174), .Y(n53498) );
  NOR2X1 U56595 ( .A(n53499), .B(n53498), .Y(n53501) );
  NOR2X1 U56596 ( .A(n19944), .B(n19943), .Y(n53500) );
  NAND2X1 U56597 ( .A(n53501), .B(n53500), .Y(u_decode_u_regfile_N638) );
  NOR2X1 U56598 ( .A(n44593), .B(n43171), .Y(n53503) );
  NOR2X1 U56599 ( .A(n44590), .B(n43174), .Y(n53502) );
  NOR2X1 U56600 ( .A(n53503), .B(n53502), .Y(n53505) );
  NOR2X1 U56601 ( .A(n18374), .B(n18373), .Y(n53504) );
  NAND2X1 U56602 ( .A(n53505), .B(n53504), .Y(u_decode_u_regfile_N934) );
  NOR2X1 U56603 ( .A(n44365), .B(n43171), .Y(n53507) );
  NOR2X1 U56604 ( .A(n44362), .B(n43174), .Y(n53506) );
  NOR2X1 U56605 ( .A(n53507), .B(n53506), .Y(n53509) );
  NOR2X1 U56606 ( .A(n22742), .B(n22741), .Y(n53508) );
  NAND2X1 U56607 ( .A(n53509), .B(n53508), .Y(u_decode_u_regfile_N1230) );
  NOR2X1 U56608 ( .A(n44443), .B(n43172), .Y(n53511) );
  NOR2X1 U56609 ( .A(n44440), .B(n37594), .Y(n53510) );
  NOR2X1 U56610 ( .A(n53511), .B(n53510), .Y(n53513) );
  NOR2X1 U56611 ( .A(n21514), .B(n21513), .Y(n53512) );
  NAND2X1 U56612 ( .A(n53513), .B(n53512), .Y(u_decode_u_regfile_N342) );
  NOR2X1 U56613 ( .A(n16471), .B(n16472), .Y(n53515) );
  NOR2X1 U56614 ( .A(n16510), .B(n16511), .Y(n53514) );
  NAND2X1 U56615 ( .A(n53515), .B(n53514), .Y(u_exec_alu_p_w[21]) );
  NOR2X1 U56616 ( .A(n44538), .B(n43178), .Y(n53517) );
  NOR2X1 U56617 ( .A(n44536), .B(n37682), .Y(n53516) );
  NOR2X1 U56618 ( .A(n53517), .B(n53516), .Y(n53519) );
  NOR2X1 U56619 ( .A(n19741), .B(n19740), .Y(n53518) );
  NAND2X1 U56620 ( .A(n53519), .B(n53518), .Y(u_decode_u_regfile_N676) );
  NOR2X1 U56621 ( .A(n44602), .B(n43178), .Y(n53521) );
  NOR2X1 U56622 ( .A(n44599), .B(n37682), .Y(n53520) );
  NOR2X1 U56623 ( .A(n53521), .B(n53520), .Y(n53523) );
  NOR2X1 U56624 ( .A(n18160), .B(n18158), .Y(n53522) );
  NAND2X1 U56625 ( .A(n53523), .B(n53522), .Y(u_decode_u_regfile_N972) );
  NOR2X1 U56626 ( .A(n43176), .B(n43271), .Y(n53525) );
  NOR2X1 U56627 ( .A(n43179), .B(n43386), .Y(n53524) );
  NOR2X1 U56628 ( .A(n53525), .B(n53524), .Y(n53527) );
  NOR2X1 U56629 ( .A(n21311), .B(n21310), .Y(n53526) );
  NAND2X1 U56630 ( .A(n53527), .B(n53526), .Y(u_decode_u_regfile_N380) );
  NOR2X1 U56631 ( .A(n44473), .B(n43178), .Y(n53529) );
  NOR2X1 U56632 ( .A(n44470), .B(n37682), .Y(n53528) );
  NOR2X1 U56633 ( .A(n53529), .B(n53528), .Y(n53531) );
  NOR2X1 U56634 ( .A(n20918), .B(n20917), .Y(n53530) );
  NAND2X1 U56635 ( .A(n53531), .B(n53530), .Y(u_decode_u_regfile_N454) );
  NOR2X1 U56636 ( .A(n44560), .B(n43178), .Y(n53533) );
  NOR2X1 U56637 ( .A(n44557), .B(n37682), .Y(n53532) );
  NOR2X1 U56638 ( .A(n53533), .B(n53532), .Y(n53535) );
  NOR2X1 U56639 ( .A(n19346), .B(n19345), .Y(n53534) );
  NAND2X1 U56640 ( .A(n53535), .B(n53534), .Y(u_decode_u_regfile_N750) );
  NOR2X1 U56641 ( .A(n44383), .B(n43177), .Y(n53537) );
  NOR2X1 U56642 ( .A(n44380), .B(n43180), .Y(n53536) );
  NOR2X1 U56643 ( .A(n53537), .B(n53536), .Y(n53539) );
  NOR2X1 U56644 ( .A(n22488), .B(n22487), .Y(n53538) );
  NAND2X1 U56645 ( .A(n53539), .B(n53538), .Y(u_decode_u_regfile_N158) );
  NOR2X1 U56646 ( .A(n44305), .B(n43177), .Y(n53541) );
  NOR2X1 U56647 ( .A(n44302), .B(n43180), .Y(n53540) );
  NOR2X1 U56648 ( .A(n53541), .B(n53540), .Y(n53543) );
  NOR2X1 U56649 ( .A(n23830), .B(n23829), .Y(n53542) );
  NAND2X1 U56650 ( .A(n53543), .B(n53542), .Y(u_decode_u_regfile_N1046) );
  NOR2X1 U56651 ( .A(n44572), .B(n43177), .Y(n53545) );
  NOR2X1 U56652 ( .A(n44569), .B(n43180), .Y(n53544) );
  NOR2X1 U56653 ( .A(n53545), .B(n53544), .Y(n53547) );
  NOR2X1 U56654 ( .A(n18954), .B(n18953), .Y(n53546) );
  NAND2X1 U56655 ( .A(n53547), .B(n53546), .Y(u_decode_u_regfile_N824) );
  NOR2X1 U56656 ( .A(n43176), .B(n43277), .Y(n53549) );
  NOR2X1 U56657 ( .A(n43179), .B(n43383), .Y(n53548) );
  NOR2X1 U56658 ( .A(n53549), .B(n53548), .Y(n53551) );
  NOR2X1 U56659 ( .A(n20526), .B(n20525), .Y(n53550) );
  NAND2X1 U56660 ( .A(n53551), .B(n53550), .Y(u_decode_u_regfile_N528) );
  NOR2X1 U56661 ( .A(n44407), .B(n43177), .Y(n53553) );
  NOR2X1 U56662 ( .A(n44404), .B(n43180), .Y(n53552) );
  NOR2X1 U56663 ( .A(n53553), .B(n53552), .Y(n53555) );
  NOR2X1 U56664 ( .A(n22096), .B(n22095), .Y(n53554) );
  NAND2X1 U56665 ( .A(n53555), .B(n53554), .Y(u_decode_u_regfile_N232) );
  NOR2X1 U56666 ( .A(n44329), .B(n43177), .Y(n53557) );
  NOR2X1 U56667 ( .A(n44326), .B(n43180), .Y(n53556) );
  NOR2X1 U56668 ( .A(n53557), .B(n53556), .Y(n53559) );
  NOR2X1 U56669 ( .A(n23390), .B(n23389), .Y(n53558) );
  NAND2X1 U56670 ( .A(n53559), .B(n53558), .Y(u_decode_u_regfile_N1120) );
  NOR2X1 U56671 ( .A(n44584), .B(n43177), .Y(n53561) );
  NOR2X1 U56672 ( .A(n44581), .B(n43180), .Y(n53560) );
  NOR2X1 U56673 ( .A(n53561), .B(n53560), .Y(n53563) );
  NOR2X1 U56674 ( .A(n18562), .B(n18561), .Y(n53562) );
  NAND2X1 U56675 ( .A(n53563), .B(n53562), .Y(u_decode_u_regfile_N898) );
  NOR2X1 U56676 ( .A(n44431), .B(n43177), .Y(n53565) );
  NOR2X1 U56677 ( .A(n44428), .B(n43180), .Y(n53564) );
  NOR2X1 U56678 ( .A(n53565), .B(n53564), .Y(n53567) );
  NOR2X1 U56679 ( .A(n21704), .B(n21703), .Y(n53566) );
  NAND2X1 U56680 ( .A(n53567), .B(n53566), .Y(u_decode_u_regfile_N306) );
  NOR2X1 U56681 ( .A(n44515), .B(n43177), .Y(n53569) );
  NOR2X1 U56682 ( .A(n44512), .B(n43180), .Y(n53568) );
  NOR2X1 U56683 ( .A(n53569), .B(n53568), .Y(n53571) );
  NOR2X1 U56684 ( .A(n20134), .B(n20133), .Y(n53570) );
  NAND2X1 U56685 ( .A(n53571), .B(n53570), .Y(u_decode_u_regfile_N602) );
  NOR2X1 U56686 ( .A(n44353), .B(n43177), .Y(n53573) );
  NOR2X1 U56687 ( .A(n44350), .B(n43180), .Y(n53572) );
  NOR2X1 U56688 ( .A(n53573), .B(n53572), .Y(n53575) );
  NOR2X1 U56689 ( .A(n22956), .B(n22955), .Y(n53574) );
  NAND2X1 U56690 ( .A(n53575), .B(n53574), .Y(u_decode_u_regfile_N1194) );
  NOR2X1 U56691 ( .A(n44608), .B(n43177), .Y(n53577) );
  NOR2X1 U56692 ( .A(n44605), .B(n43180), .Y(n53576) );
  NOR2X1 U56693 ( .A(n53577), .B(n53576), .Y(n53579) );
  NOR2X1 U56694 ( .A(n24046), .B(n24045), .Y(n53578) );
  NAND2X1 U56695 ( .A(n53579), .B(n53578), .Y(u_decode_u_regfile_N1009) );
  NOR2X1 U56696 ( .A(n43176), .B(n43274), .Y(n53581) );
  NOR2X1 U56697 ( .A(n43179), .B(n43389), .Y(n53580) );
  NOR2X1 U56698 ( .A(n53581), .B(n53580), .Y(n53583) );
  NOR2X1 U56699 ( .A(n22880), .B(n22879), .Y(n53582) );
  NAND2X1 U56700 ( .A(n53583), .B(n53582), .Y(u_decode_u_regfile_N121) );
  NOR2X1 U56701 ( .A(n44461), .B(n43177), .Y(n53585) );
  NOR2X1 U56702 ( .A(n44458), .B(n43180), .Y(n53584) );
  NOR2X1 U56703 ( .A(n53585), .B(n53584), .Y(n53587) );
  NOR2X1 U56704 ( .A(n21114), .B(n21113), .Y(n53586) );
  NAND2X1 U56705 ( .A(n53587), .B(n53586), .Y(u_decode_u_regfile_N417) );
  NOR2X1 U56706 ( .A(n44551), .B(n43177), .Y(n53589) );
  NOR2X1 U56707 ( .A(n44548), .B(n43180), .Y(n53588) );
  NOR2X1 U56708 ( .A(n53589), .B(n53588), .Y(n53591) );
  NOR2X1 U56709 ( .A(n19544), .B(n19543), .Y(n53590) );
  NAND2X1 U56710 ( .A(n53591), .B(n53590), .Y(u_decode_u_regfile_N713) );
  NOR2X1 U56711 ( .A(n44566), .B(n43176), .Y(n53593) );
  NOR2X1 U56712 ( .A(n44563), .B(n43179), .Y(n53592) );
  NOR2X1 U56713 ( .A(n53593), .B(n53592), .Y(n53595) );
  NOR2X1 U56714 ( .A(n19150), .B(n19149), .Y(n53594) );
  NAND2X1 U56715 ( .A(n53595), .B(n53594), .Y(u_decode_u_regfile_N787) );
  NOR2X1 U56716 ( .A(n44317), .B(n43176), .Y(n53597) );
  NOR2X1 U56717 ( .A(n44314), .B(n43179), .Y(n53596) );
  NOR2X1 U56718 ( .A(n53597), .B(n53596), .Y(n53599) );
  NOR2X1 U56719 ( .A(n23610), .B(n23609), .Y(n53598) );
  NAND2X1 U56720 ( .A(n53599), .B(n53598), .Y(u_decode_u_regfile_N1083) );
  NOR2X1 U56721 ( .A(n44395), .B(n43176), .Y(n53601) );
  NOR2X1 U56722 ( .A(n44392), .B(n43179), .Y(n53600) );
  NOR2X1 U56723 ( .A(n53601), .B(n53600), .Y(n53603) );
  NOR2X1 U56724 ( .A(n22292), .B(n22291), .Y(n53602) );
  NAND2X1 U56725 ( .A(n53603), .B(n53602), .Y(u_decode_u_regfile_N195) );
  NOR2X1 U56726 ( .A(n44485), .B(n43177), .Y(n53605) );
  NOR2X1 U56727 ( .A(n44482), .B(n43179), .Y(n53604) );
  NOR2X1 U56728 ( .A(n53605), .B(n53604), .Y(n53607) );
  NOR2X1 U56729 ( .A(n20722), .B(n20721), .Y(n53606) );
  NAND2X1 U56730 ( .A(n53607), .B(n53606), .Y(u_decode_u_regfile_N491) );
  NOR2X1 U56731 ( .A(n44419), .B(n43176), .Y(n53609) );
  NOR2X1 U56732 ( .A(n44416), .B(n43179), .Y(n53608) );
  NOR2X1 U56733 ( .A(n53609), .B(n53608), .Y(n53611) );
  NOR2X1 U56734 ( .A(n21900), .B(n21899), .Y(n53610) );
  NAND2X1 U56735 ( .A(n53611), .B(n53610), .Y(u_decode_u_regfile_N269) );
  NOR2X1 U56736 ( .A(n44341), .B(n43176), .Y(n53613) );
  NOR2X1 U56737 ( .A(n44338), .B(n43179), .Y(n53612) );
  NOR2X1 U56738 ( .A(n53613), .B(n53612), .Y(n53615) );
  NOR2X1 U56739 ( .A(n23176), .B(n23175), .Y(n53614) );
  NAND2X1 U56740 ( .A(n53615), .B(n53614), .Y(u_decode_u_regfile_N1157) );
  NOR2X1 U56741 ( .A(n44503), .B(n43176), .Y(n53617) );
  NOR2X1 U56742 ( .A(n44500), .B(n43179), .Y(n53616) );
  NOR2X1 U56743 ( .A(n53617), .B(n53616), .Y(n53619) );
  NOR2X1 U56744 ( .A(n20330), .B(n20329), .Y(n53618) );
  NAND2X1 U56745 ( .A(n53619), .B(n53618), .Y(u_decode_u_regfile_N565) );
  NOR2X1 U56746 ( .A(n44578), .B(n43176), .Y(n53621) );
  NOR2X1 U56747 ( .A(n44575), .B(n43179), .Y(n53620) );
  NOR2X1 U56748 ( .A(n53621), .B(n53620), .Y(n53623) );
  NOR2X1 U56749 ( .A(n18758), .B(n18757), .Y(n53622) );
  NAND2X1 U56750 ( .A(n53623), .B(n53622), .Y(u_decode_u_regfile_N861) );
  NOR2X1 U56751 ( .A(n44527), .B(n43176), .Y(n53625) );
  NOR2X1 U56752 ( .A(n44524), .B(n43179), .Y(n53624) );
  NOR2X1 U56753 ( .A(n53625), .B(n53624), .Y(n53627) );
  NOR2X1 U56754 ( .A(n19938), .B(n19937), .Y(n53626) );
  NAND2X1 U56755 ( .A(n53627), .B(n53626), .Y(u_decode_u_regfile_N639) );
  NOR2X1 U56756 ( .A(n44593), .B(n43176), .Y(n53629) );
  NOR2X1 U56757 ( .A(n44590), .B(n43180), .Y(n53628) );
  NOR2X1 U56758 ( .A(n53629), .B(n53628), .Y(n53631) );
  NOR2X1 U56759 ( .A(n18368), .B(n18367), .Y(n53630) );
  NAND2X1 U56760 ( .A(n53631), .B(n53630), .Y(u_decode_u_regfile_N935) );
  NOR2X1 U56761 ( .A(n44365), .B(n43176), .Y(n53633) );
  NOR2X1 U56762 ( .A(n44362), .B(n43179), .Y(n53632) );
  NOR2X1 U56763 ( .A(n53633), .B(n53632), .Y(n53635) );
  NOR2X1 U56764 ( .A(n22736), .B(n22735), .Y(n53634) );
  NAND2X1 U56765 ( .A(n53635), .B(n53634), .Y(u_decode_u_regfile_N1231) );
  NOR2X1 U56766 ( .A(n44443), .B(n43177), .Y(n53637) );
  NOR2X1 U56767 ( .A(n44440), .B(n43180), .Y(n53636) );
  NOR2X1 U56768 ( .A(n53637), .B(n53636), .Y(n53639) );
  NOR2X1 U56769 ( .A(n21508), .B(n21507), .Y(n53638) );
  NAND2X1 U56770 ( .A(n53639), .B(n53638), .Y(u_decode_u_regfile_N343) );
  NOR2X1 U56771 ( .A(n16416), .B(n16417), .Y(n53641) );
  NOR2X1 U56772 ( .A(n16454), .B(n16455), .Y(n53640) );
  NAND2X1 U56773 ( .A(n53641), .B(n53640), .Y(u_exec_alu_p_w[22]) );
  NOR2X1 U56774 ( .A(n44538), .B(n53762), .Y(n53643) );
  NOR2X1 U56775 ( .A(n44536), .B(n37683), .Y(n53642) );
  NOR2X1 U56776 ( .A(n53643), .B(n53642), .Y(n53645) );
  NOR2X1 U56777 ( .A(n19735), .B(n19734), .Y(n53644) );
  NAND2X1 U56778 ( .A(n53645), .B(n53644), .Y(u_decode_u_regfile_N677) );
  NOR2X1 U56779 ( .A(n44602), .B(n53762), .Y(n53647) );
  NOR2X1 U56780 ( .A(n44599), .B(n37683), .Y(n53646) );
  NOR2X1 U56781 ( .A(n53647), .B(n53646), .Y(n53649) );
  NOR2X1 U56782 ( .A(n18153), .B(n18151), .Y(n53648) );
  NAND2X1 U56783 ( .A(n53649), .B(n53648), .Y(u_decode_u_regfile_N973) );
  NOR2X1 U56784 ( .A(n43182), .B(n43271), .Y(n53651) );
  NOR2X1 U56785 ( .A(n43185), .B(n43386), .Y(n53650) );
  NOR2X1 U56786 ( .A(n53651), .B(n53650), .Y(n53653) );
  NOR2X1 U56787 ( .A(n21305), .B(n21304), .Y(n53652) );
  NAND2X1 U56788 ( .A(n53653), .B(n53652), .Y(u_decode_u_regfile_N381) );
  NOR2X1 U56789 ( .A(n44473), .B(n53762), .Y(n53655) );
  NOR2X1 U56790 ( .A(n44470), .B(n37683), .Y(n53654) );
  NOR2X1 U56791 ( .A(n53655), .B(n53654), .Y(n53657) );
  NOR2X1 U56792 ( .A(n20912), .B(n20911), .Y(n53656) );
  NAND2X1 U56793 ( .A(n53657), .B(n53656), .Y(u_decode_u_regfile_N455) );
  NOR2X1 U56794 ( .A(n44560), .B(n53762), .Y(n53659) );
  NOR2X1 U56795 ( .A(n44557), .B(n37683), .Y(n53658) );
  NOR2X1 U56796 ( .A(n53659), .B(n53658), .Y(n53661) );
  NOR2X1 U56797 ( .A(n19340), .B(n19339), .Y(n53660) );
  NAND2X1 U56798 ( .A(n53661), .B(n53660), .Y(u_decode_u_regfile_N751) );
  NOR2X1 U56799 ( .A(n44383), .B(n43183), .Y(n53663) );
  NOR2X1 U56800 ( .A(n44380), .B(n43186), .Y(n53662) );
  NOR2X1 U56801 ( .A(n53663), .B(n53662), .Y(n53665) );
  NOR2X1 U56802 ( .A(n22482), .B(n22481), .Y(n53664) );
  NAND2X1 U56803 ( .A(n53665), .B(n53664), .Y(u_decode_u_regfile_N159) );
  NOR2X1 U56804 ( .A(n44305), .B(n43183), .Y(n53667) );
  NOR2X1 U56805 ( .A(n44302), .B(n43186), .Y(n53666) );
  NOR2X1 U56806 ( .A(n53667), .B(n53666), .Y(n53669) );
  NOR2X1 U56807 ( .A(n23824), .B(n23823), .Y(n53668) );
  NAND2X1 U56808 ( .A(n53669), .B(n53668), .Y(u_decode_u_regfile_N1047) );
  NOR2X1 U56809 ( .A(n44572), .B(n43183), .Y(n53671) );
  NOR2X1 U56810 ( .A(n44569), .B(n43186), .Y(n53670) );
  NOR2X1 U56811 ( .A(n53671), .B(n53670), .Y(n53673) );
  NOR2X1 U56812 ( .A(n18948), .B(n18947), .Y(n53672) );
  NAND2X1 U56813 ( .A(n53673), .B(n53672), .Y(u_decode_u_regfile_N825) );
  NOR2X1 U56814 ( .A(n43182), .B(n43277), .Y(n53675) );
  NOR2X1 U56815 ( .A(n43185), .B(n43383), .Y(n53674) );
  NOR2X1 U56816 ( .A(n53675), .B(n53674), .Y(n53677) );
  NOR2X1 U56817 ( .A(n20520), .B(n20519), .Y(n53676) );
  NAND2X1 U56818 ( .A(n53677), .B(n53676), .Y(u_decode_u_regfile_N529) );
  NOR2X1 U56819 ( .A(n44407), .B(n43183), .Y(n53679) );
  NOR2X1 U56820 ( .A(n44404), .B(n43186), .Y(n53678) );
  NOR2X1 U56821 ( .A(n53679), .B(n53678), .Y(n53681) );
  NOR2X1 U56822 ( .A(n22090), .B(n22089), .Y(n53680) );
  NAND2X1 U56823 ( .A(n53681), .B(n53680), .Y(u_decode_u_regfile_N233) );
  NOR2X1 U56824 ( .A(n44329), .B(n43183), .Y(n53683) );
  NOR2X1 U56825 ( .A(n44326), .B(n43186), .Y(n53682) );
  NOR2X1 U56826 ( .A(n53683), .B(n53682), .Y(n53685) );
  NOR2X1 U56827 ( .A(n23384), .B(n23383), .Y(n53684) );
  NAND2X1 U56828 ( .A(n53685), .B(n53684), .Y(u_decode_u_regfile_N1121) );
  NOR2X1 U56829 ( .A(n44584), .B(n43183), .Y(n53687) );
  NOR2X1 U56830 ( .A(n44581), .B(n43186), .Y(n53686) );
  NOR2X1 U56831 ( .A(n53687), .B(n53686), .Y(n53689) );
  NOR2X1 U56832 ( .A(n18556), .B(n18555), .Y(n53688) );
  NAND2X1 U56833 ( .A(n53689), .B(n53688), .Y(u_decode_u_regfile_N899) );
  NOR2X1 U56834 ( .A(n44431), .B(n43183), .Y(n53691) );
  NOR2X1 U56835 ( .A(n44428), .B(n43186), .Y(n53690) );
  NOR2X1 U56836 ( .A(n53691), .B(n53690), .Y(n53693) );
  NOR2X1 U56837 ( .A(n21698), .B(n21697), .Y(n53692) );
  NAND2X1 U56838 ( .A(n53693), .B(n53692), .Y(u_decode_u_regfile_N307) );
  NOR2X1 U56839 ( .A(n44515), .B(n43183), .Y(n53695) );
  NOR2X1 U56840 ( .A(n44512), .B(n43186), .Y(n53694) );
  NOR2X1 U56841 ( .A(n53695), .B(n53694), .Y(n53697) );
  NOR2X1 U56842 ( .A(n20128), .B(n20127), .Y(n53696) );
  NAND2X1 U56843 ( .A(n53697), .B(n53696), .Y(u_decode_u_regfile_N603) );
  NOR2X1 U56844 ( .A(n44353), .B(n43183), .Y(n53699) );
  NOR2X1 U56845 ( .A(n44350), .B(n43186), .Y(n53698) );
  NOR2X1 U56846 ( .A(n53699), .B(n53698), .Y(n53701) );
  NOR2X1 U56847 ( .A(n22950), .B(n22949), .Y(n53700) );
  NAND2X1 U56848 ( .A(n53701), .B(n53700), .Y(u_decode_u_regfile_N1195) );
  NOR2X1 U56849 ( .A(n44608), .B(n43183), .Y(n53703) );
  NOR2X1 U56850 ( .A(n44605), .B(n43186), .Y(n53702) );
  NOR2X1 U56851 ( .A(n53703), .B(n53702), .Y(n53705) );
  NOR2X1 U56852 ( .A(n24034), .B(n24033), .Y(n53704) );
  NAND2X1 U56853 ( .A(n53705), .B(n53704), .Y(u_decode_u_regfile_N1010) );
  NOR2X1 U56854 ( .A(n43182), .B(n43274), .Y(n53707) );
  NOR2X1 U56855 ( .A(n43185), .B(n43389), .Y(n53706) );
  NOR2X1 U56856 ( .A(n53707), .B(n53706), .Y(n53709) );
  NOR2X1 U56857 ( .A(n22814), .B(n22813), .Y(n53708) );
  NAND2X1 U56858 ( .A(n53709), .B(n53708), .Y(u_decode_u_regfile_N122) );
  NOR2X1 U56859 ( .A(n44461), .B(n43183), .Y(n53711) );
  NOR2X1 U56860 ( .A(n44458), .B(n43186), .Y(n53710) );
  NOR2X1 U56861 ( .A(n53711), .B(n53710), .Y(n53713) );
  NOR2X1 U56862 ( .A(n21108), .B(n21107), .Y(n53712) );
  NAND2X1 U56863 ( .A(n53713), .B(n53712), .Y(u_decode_u_regfile_N418) );
  NOR2X1 U56864 ( .A(n44551), .B(n43183), .Y(n53715) );
  NOR2X1 U56865 ( .A(n44548), .B(n43186), .Y(n53714) );
  NOR2X1 U56866 ( .A(n53715), .B(n53714), .Y(n53717) );
  NOR2X1 U56867 ( .A(n19538), .B(n19537), .Y(n53716) );
  NAND2X1 U56868 ( .A(n53717), .B(n53716), .Y(u_decode_u_regfile_N714) );
  NOR2X1 U56869 ( .A(n44566), .B(n43182), .Y(n53719) );
  NOR2X1 U56870 ( .A(n44563), .B(n43185), .Y(n53718) );
  NOR2X1 U56871 ( .A(n53719), .B(n53718), .Y(n53721) );
  NOR2X1 U56872 ( .A(n19144), .B(n19143), .Y(n53720) );
  NAND2X1 U56873 ( .A(n53721), .B(n53720), .Y(u_decode_u_regfile_N788) );
  NOR2X1 U56874 ( .A(n44317), .B(n43182), .Y(n53723) );
  NOR2X1 U56875 ( .A(n44314), .B(n43185), .Y(n53722) );
  NOR2X1 U56876 ( .A(n53723), .B(n53722), .Y(n53725) );
  NOR2X1 U56877 ( .A(n23604), .B(n23603), .Y(n53724) );
  NAND2X1 U56878 ( .A(n53725), .B(n53724), .Y(u_decode_u_regfile_N1084) );
  NOR2X1 U56879 ( .A(n44395), .B(n43182), .Y(n53727) );
  NOR2X1 U56880 ( .A(n44392), .B(n43185), .Y(n53726) );
  NOR2X1 U56881 ( .A(n53727), .B(n53726), .Y(n53729) );
  NOR2X1 U56882 ( .A(n22286), .B(n22285), .Y(n53728) );
  NAND2X1 U56883 ( .A(n53729), .B(n53728), .Y(u_decode_u_regfile_N196) );
  NOR2X1 U56884 ( .A(n44485), .B(n43182), .Y(n53731) );
  NOR2X1 U56885 ( .A(n44482), .B(n43185), .Y(n53730) );
  NOR2X1 U56886 ( .A(n53731), .B(n53730), .Y(n53733) );
  NOR2X1 U56887 ( .A(n20716), .B(n20715), .Y(n53732) );
  NAND2X1 U56888 ( .A(n53733), .B(n53732), .Y(u_decode_u_regfile_N492) );
  NOR2X1 U56889 ( .A(n44419), .B(n43182), .Y(n53735) );
  NOR2X1 U56890 ( .A(n44416), .B(n43185), .Y(n53734) );
  NOR2X1 U56891 ( .A(n53735), .B(n53734), .Y(n53737) );
  NOR2X1 U56892 ( .A(n21894), .B(n21893), .Y(n53736) );
  NAND2X1 U56893 ( .A(n53737), .B(n53736), .Y(u_decode_u_regfile_N270) );
  NOR2X1 U56894 ( .A(n44341), .B(n43182), .Y(n53739) );
  NOR2X1 U56895 ( .A(n44338), .B(n43185), .Y(n53738) );
  NOR2X1 U56896 ( .A(n53739), .B(n53738), .Y(n53741) );
  NOR2X1 U56897 ( .A(n23170), .B(n23169), .Y(n53740) );
  NAND2X1 U56898 ( .A(n53741), .B(n53740), .Y(u_decode_u_regfile_N1158) );
  NOR2X1 U56899 ( .A(n44503), .B(n43182), .Y(n53743) );
  NOR2X1 U56900 ( .A(n44500), .B(n43185), .Y(n53742) );
  NOR2X1 U56901 ( .A(n53743), .B(n53742), .Y(n53745) );
  NOR2X1 U56902 ( .A(n20324), .B(n20323), .Y(n53744) );
  NAND2X1 U56903 ( .A(n53745), .B(n53744), .Y(u_decode_u_regfile_N566) );
  NOR2X1 U56904 ( .A(n44578), .B(n43182), .Y(n53747) );
  NOR2X1 U56905 ( .A(n44575), .B(n43185), .Y(n53746) );
  NOR2X1 U56906 ( .A(n53747), .B(n53746), .Y(n53749) );
  NOR2X1 U56907 ( .A(n18752), .B(n18751), .Y(n53748) );
  NAND2X1 U56908 ( .A(n53749), .B(n53748), .Y(u_decode_u_regfile_N862) );
  NOR2X1 U56909 ( .A(n44527), .B(n43182), .Y(n53751) );
  NOR2X1 U56910 ( .A(n44524), .B(n43185), .Y(n53750) );
  NOR2X1 U56911 ( .A(n53751), .B(n53750), .Y(n53753) );
  NOR2X1 U56912 ( .A(n19932), .B(n19931), .Y(n53752) );
  NAND2X1 U56913 ( .A(n53753), .B(n53752), .Y(u_decode_u_regfile_N640) );
  NOR2X1 U56914 ( .A(n44593), .B(n43183), .Y(n53755) );
  NOR2X1 U56915 ( .A(n44590), .B(n43186), .Y(n53754) );
  NOR2X1 U56916 ( .A(n53755), .B(n53754), .Y(n53757) );
  NOR2X1 U56917 ( .A(n18362), .B(n18361), .Y(n53756) );
  NAND2X1 U56918 ( .A(n53757), .B(n53756), .Y(u_decode_u_regfile_N936) );
  NOR2X1 U56919 ( .A(n44365), .B(n43182), .Y(n53759) );
  NOR2X1 U56920 ( .A(n44362), .B(n43185), .Y(n53758) );
  NOR2X1 U56921 ( .A(n53759), .B(n53758), .Y(n53761) );
  NOR2X1 U56922 ( .A(n22730), .B(n22729), .Y(n53760) );
  NAND2X1 U56923 ( .A(n53761), .B(n53760), .Y(u_decode_u_regfile_N1232) );
  NOR2X1 U56924 ( .A(n44443), .B(n43183), .Y(n53764) );
  NOR2X1 U56925 ( .A(n44440), .B(n43186), .Y(n53763) );
  NOR2X1 U56926 ( .A(n53764), .B(n53763), .Y(n53766) );
  NOR2X1 U56927 ( .A(n21502), .B(n21501), .Y(n53765) );
  NAND2X1 U56928 ( .A(n53766), .B(n53765), .Y(u_decode_u_regfile_N344) );
  NOR2X1 U56929 ( .A(n16363), .B(n16364), .Y(n53768) );
  NOR2X1 U56930 ( .A(n16400), .B(n16401), .Y(n53767) );
  NAND2X1 U56931 ( .A(n53768), .B(n53767), .Y(u_exec_alu_p_w[23]) );
  NOR2X1 U56932 ( .A(n44538), .B(n53889), .Y(n53770) );
  NOR2X1 U56933 ( .A(n44536), .B(n37684), .Y(n53769) );
  NOR2X1 U56934 ( .A(n53770), .B(n53769), .Y(n53772) );
  NOR2X1 U56935 ( .A(n19729), .B(n19728), .Y(n53771) );
  NAND2X1 U56936 ( .A(n53772), .B(n53771), .Y(u_decode_u_regfile_N678) );
  NOR2X1 U56937 ( .A(n44602), .B(n53889), .Y(n53774) );
  NOR2X1 U56938 ( .A(n44599), .B(n37684), .Y(n53773) );
  NOR2X1 U56939 ( .A(n53774), .B(n53773), .Y(n53776) );
  NOR2X1 U56940 ( .A(n18146), .B(n18144), .Y(n53775) );
  NAND2X1 U56941 ( .A(n53776), .B(n53775), .Y(u_decode_u_regfile_N974) );
  NOR2X1 U56942 ( .A(n43188), .B(n43271), .Y(n53778) );
  NOR2X1 U56943 ( .A(n43191), .B(n43386), .Y(n53777) );
  NOR2X1 U56944 ( .A(n53778), .B(n53777), .Y(n53780) );
  NOR2X1 U56945 ( .A(n21299), .B(n21298), .Y(n53779) );
  NAND2X1 U56946 ( .A(n53780), .B(n53779), .Y(u_decode_u_regfile_N382) );
  NOR2X1 U56947 ( .A(n44473), .B(n53889), .Y(n53782) );
  NOR2X1 U56948 ( .A(n44470), .B(n37684), .Y(n53781) );
  NOR2X1 U56949 ( .A(n53782), .B(n53781), .Y(n53784) );
  NOR2X1 U56950 ( .A(n20906), .B(n20905), .Y(n53783) );
  NAND2X1 U56951 ( .A(n53784), .B(n53783), .Y(u_decode_u_regfile_N456) );
  NOR2X1 U56952 ( .A(n44560), .B(n53889), .Y(n53786) );
  NOR2X1 U56953 ( .A(n44557), .B(n37684), .Y(n53785) );
  NOR2X1 U56954 ( .A(n53786), .B(n53785), .Y(n53788) );
  NOR2X1 U56955 ( .A(n19334), .B(n19333), .Y(n53787) );
  NAND2X1 U56956 ( .A(n53788), .B(n53787), .Y(u_decode_u_regfile_N752) );
  NOR2X1 U56957 ( .A(n44383), .B(n43189), .Y(n53790) );
  NOR2X1 U56958 ( .A(n44380), .B(n43192), .Y(n53789) );
  NOR2X1 U56959 ( .A(n53790), .B(n53789), .Y(n53792) );
  NOR2X1 U56960 ( .A(n22476), .B(n22475), .Y(n53791) );
  NAND2X1 U56961 ( .A(n53792), .B(n53791), .Y(u_decode_u_regfile_N160) );
  NOR2X1 U56962 ( .A(n44305), .B(n43189), .Y(n53794) );
  NOR2X1 U56963 ( .A(n44302), .B(n43192), .Y(n53793) );
  NOR2X1 U56964 ( .A(n53794), .B(n53793), .Y(n53796) );
  NOR2X1 U56965 ( .A(n23818), .B(n23817), .Y(n53795) );
  NAND2X1 U56966 ( .A(n53796), .B(n53795), .Y(u_decode_u_regfile_N1048) );
  NOR2X1 U56967 ( .A(n44572), .B(n43189), .Y(n53798) );
  NOR2X1 U56968 ( .A(n44569), .B(n43192), .Y(n53797) );
  NOR2X1 U56969 ( .A(n53798), .B(n53797), .Y(n53800) );
  NOR2X1 U56970 ( .A(n18942), .B(n18941), .Y(n53799) );
  NAND2X1 U56971 ( .A(n53800), .B(n53799), .Y(u_decode_u_regfile_N826) );
  NOR2X1 U56972 ( .A(n43188), .B(n43277), .Y(n53802) );
  NOR2X1 U56973 ( .A(n43191), .B(n43383), .Y(n53801) );
  NOR2X1 U56974 ( .A(n53802), .B(n53801), .Y(n53804) );
  NOR2X1 U56975 ( .A(n20514), .B(n20513), .Y(n53803) );
  NAND2X1 U56976 ( .A(n53804), .B(n53803), .Y(u_decode_u_regfile_N530) );
  NOR2X1 U56977 ( .A(n44407), .B(n43189), .Y(n53806) );
  NOR2X1 U56978 ( .A(n44404), .B(n43192), .Y(n53805) );
  NOR2X1 U56979 ( .A(n53806), .B(n53805), .Y(n53808) );
  NOR2X1 U56980 ( .A(n22084), .B(n22083), .Y(n53807) );
  NAND2X1 U56981 ( .A(n53808), .B(n53807), .Y(u_decode_u_regfile_N234) );
  NOR2X1 U56982 ( .A(n44329), .B(n43189), .Y(n53810) );
  NOR2X1 U56983 ( .A(n44326), .B(n43192), .Y(n53809) );
  NOR2X1 U56984 ( .A(n53810), .B(n53809), .Y(n53812) );
  NOR2X1 U56985 ( .A(n23378), .B(n23377), .Y(n53811) );
  NAND2X1 U56986 ( .A(n53812), .B(n53811), .Y(u_decode_u_regfile_N1122) );
  NOR2X1 U56987 ( .A(n44584), .B(n43189), .Y(n53814) );
  NOR2X1 U56988 ( .A(n44581), .B(n43192), .Y(n53813) );
  NOR2X1 U56989 ( .A(n53814), .B(n53813), .Y(n53816) );
  NOR2X1 U56990 ( .A(n18550), .B(n18549), .Y(n53815) );
  NAND2X1 U56991 ( .A(n53816), .B(n53815), .Y(u_decode_u_regfile_N900) );
  NOR2X1 U56992 ( .A(n44431), .B(n43189), .Y(n53818) );
  NOR2X1 U56993 ( .A(n44428), .B(n43192), .Y(n53817) );
  NOR2X1 U56994 ( .A(n53818), .B(n53817), .Y(n53820) );
  NOR2X1 U56995 ( .A(n21692), .B(n21691), .Y(n53819) );
  NAND2X1 U56996 ( .A(n53820), .B(n53819), .Y(u_decode_u_regfile_N308) );
  NOR2X1 U56997 ( .A(n44515), .B(n43189), .Y(n53822) );
  NOR2X1 U56998 ( .A(n44512), .B(n43192), .Y(n53821) );
  NOR2X1 U56999 ( .A(n53822), .B(n53821), .Y(n53824) );
  NOR2X1 U57000 ( .A(n20122), .B(n20121), .Y(n53823) );
  NAND2X1 U57001 ( .A(n53824), .B(n53823), .Y(u_decode_u_regfile_N604) );
  NOR2X1 U57002 ( .A(n44353), .B(n43189), .Y(n53826) );
  NOR2X1 U57003 ( .A(n44350), .B(n43192), .Y(n53825) );
  NOR2X1 U57004 ( .A(n53826), .B(n53825), .Y(n53828) );
  NOR2X1 U57005 ( .A(n22944), .B(n22943), .Y(n53827) );
  NAND2X1 U57006 ( .A(n53828), .B(n53827), .Y(u_decode_u_regfile_N1196) );
  NOR2X1 U57007 ( .A(n44608), .B(n43189), .Y(n53830) );
  NOR2X1 U57008 ( .A(n44605), .B(n43192), .Y(n53829) );
  NOR2X1 U57009 ( .A(n53830), .B(n53829), .Y(n53832) );
  NOR2X1 U57010 ( .A(n24028), .B(n24027), .Y(n53831) );
  NAND2X1 U57011 ( .A(n53832), .B(n53831), .Y(u_decode_u_regfile_N1011) );
  NOR2X1 U57012 ( .A(n43188), .B(n43274), .Y(n53834) );
  NOR2X1 U57013 ( .A(n43191), .B(n43389), .Y(n53833) );
  NOR2X1 U57014 ( .A(n53834), .B(n53833), .Y(n53836) );
  NOR2X1 U57015 ( .A(n22748), .B(n22747), .Y(n53835) );
  NAND2X1 U57016 ( .A(n53836), .B(n53835), .Y(u_decode_u_regfile_N123) );
  NOR2X1 U57017 ( .A(n44461), .B(n43189), .Y(n53838) );
  NOR2X1 U57018 ( .A(n44458), .B(n43192), .Y(n53837) );
  NOR2X1 U57019 ( .A(n53838), .B(n53837), .Y(n53840) );
  NOR2X1 U57020 ( .A(n21102), .B(n21101), .Y(n53839) );
  NAND2X1 U57021 ( .A(n53840), .B(n53839), .Y(u_decode_u_regfile_N419) );
  NOR2X1 U57022 ( .A(n44551), .B(n43189), .Y(n53842) );
  NOR2X1 U57023 ( .A(n44548), .B(n43192), .Y(n53841) );
  NOR2X1 U57024 ( .A(n53842), .B(n53841), .Y(n53844) );
  NOR2X1 U57025 ( .A(n19532), .B(n19531), .Y(n53843) );
  NAND2X1 U57026 ( .A(n53844), .B(n53843), .Y(u_decode_u_regfile_N715) );
  NOR2X1 U57027 ( .A(n44566), .B(n43188), .Y(n53846) );
  NOR2X1 U57028 ( .A(n44563), .B(n43191), .Y(n53845) );
  NOR2X1 U57029 ( .A(n53846), .B(n53845), .Y(n53848) );
  NOR2X1 U57030 ( .A(n19138), .B(n19137), .Y(n53847) );
  NAND2X1 U57031 ( .A(n53848), .B(n53847), .Y(u_decode_u_regfile_N789) );
  NOR2X1 U57032 ( .A(n44317), .B(n43188), .Y(n53850) );
  NOR2X1 U57033 ( .A(n44314), .B(n43191), .Y(n53849) );
  NOR2X1 U57034 ( .A(n53850), .B(n53849), .Y(n53852) );
  NOR2X1 U57035 ( .A(n23598), .B(n23597), .Y(n53851) );
  NAND2X1 U57036 ( .A(n53852), .B(n53851), .Y(u_decode_u_regfile_N1085) );
  NOR2X1 U57037 ( .A(n44395), .B(n43188), .Y(n53854) );
  NOR2X1 U57038 ( .A(n44392), .B(n43191), .Y(n53853) );
  NOR2X1 U57039 ( .A(n53854), .B(n53853), .Y(n53856) );
  NOR2X1 U57040 ( .A(n22280), .B(n22279), .Y(n53855) );
  NAND2X1 U57041 ( .A(n53856), .B(n53855), .Y(u_decode_u_regfile_N197) );
  NOR2X1 U57042 ( .A(n44485), .B(n43188), .Y(n53858) );
  NOR2X1 U57043 ( .A(n44482), .B(n43191), .Y(n53857) );
  NOR2X1 U57044 ( .A(n53858), .B(n53857), .Y(n53860) );
  NOR2X1 U57045 ( .A(n20710), .B(n20709), .Y(n53859) );
  NAND2X1 U57046 ( .A(n53860), .B(n53859), .Y(u_decode_u_regfile_N493) );
  NOR2X1 U57047 ( .A(n44419), .B(n43188), .Y(n53862) );
  NOR2X1 U57048 ( .A(n44416), .B(n43191), .Y(n53861) );
  NOR2X1 U57049 ( .A(n53862), .B(n53861), .Y(n53864) );
  NOR2X1 U57050 ( .A(n21888), .B(n21887), .Y(n53863) );
  NAND2X1 U57051 ( .A(n53864), .B(n53863), .Y(u_decode_u_regfile_N271) );
  NOR2X1 U57052 ( .A(n44341), .B(n43188), .Y(n53866) );
  NOR2X1 U57053 ( .A(n44338), .B(n43191), .Y(n53865) );
  NOR2X1 U57054 ( .A(n53866), .B(n53865), .Y(n53868) );
  NOR2X1 U57055 ( .A(n23164), .B(n23163), .Y(n53867) );
  NAND2X1 U57056 ( .A(n53868), .B(n53867), .Y(u_decode_u_regfile_N1159) );
  NOR2X1 U57057 ( .A(n44503), .B(n43188), .Y(n53870) );
  NOR2X1 U57058 ( .A(n44500), .B(n43191), .Y(n53869) );
  NOR2X1 U57059 ( .A(n53870), .B(n53869), .Y(n53872) );
  NOR2X1 U57060 ( .A(n20318), .B(n20317), .Y(n53871) );
  NAND2X1 U57061 ( .A(n53872), .B(n53871), .Y(u_decode_u_regfile_N567) );
  NOR2X1 U57062 ( .A(n44578), .B(n43188), .Y(n53874) );
  NOR2X1 U57063 ( .A(n44575), .B(n43191), .Y(n53873) );
  NOR2X1 U57064 ( .A(n53874), .B(n53873), .Y(n53876) );
  NOR2X1 U57065 ( .A(n18746), .B(n18745), .Y(n53875) );
  NAND2X1 U57066 ( .A(n53876), .B(n53875), .Y(u_decode_u_regfile_N863) );
  NOR2X1 U57067 ( .A(n44527), .B(n43188), .Y(n53878) );
  NOR2X1 U57068 ( .A(n44524), .B(n43191), .Y(n53877) );
  NOR2X1 U57069 ( .A(n53878), .B(n53877), .Y(n53880) );
  NOR2X1 U57070 ( .A(n19926), .B(n19925), .Y(n53879) );
  NAND2X1 U57071 ( .A(n53880), .B(n53879), .Y(u_decode_u_regfile_N641) );
  NOR2X1 U57072 ( .A(n44593), .B(n43189), .Y(n53882) );
  NOR2X1 U57073 ( .A(n44590), .B(n43192), .Y(n53881) );
  NOR2X1 U57074 ( .A(n53882), .B(n53881), .Y(n53884) );
  NOR2X1 U57075 ( .A(n18356), .B(n18355), .Y(n53883) );
  NAND2X1 U57076 ( .A(n53884), .B(n53883), .Y(u_decode_u_regfile_N937) );
  NOR2X1 U57077 ( .A(n44365), .B(n43188), .Y(n53886) );
  NOR2X1 U57078 ( .A(n44362), .B(n43191), .Y(n53885) );
  NOR2X1 U57079 ( .A(n53886), .B(n53885), .Y(n53888) );
  NOR2X1 U57080 ( .A(n22724), .B(n22723), .Y(n53887) );
  NAND2X1 U57081 ( .A(n53888), .B(n53887), .Y(u_decode_u_regfile_N1233) );
  NOR2X1 U57082 ( .A(n44443), .B(n43189), .Y(n53891) );
  NOR2X1 U57083 ( .A(n44440), .B(n43192), .Y(n53890) );
  NOR2X1 U57084 ( .A(n53891), .B(n53890), .Y(n53893) );
  NOR2X1 U57085 ( .A(n21496), .B(n21495), .Y(n53892) );
  NAND2X1 U57086 ( .A(n53893), .B(n53892), .Y(u_decode_u_regfile_N345) );
  NOR2X1 U57087 ( .A(n16304), .B(n16305), .Y(n53895) );
  NOR2X1 U57088 ( .A(n16344), .B(n16345), .Y(n53894) );
  NAND2X1 U57089 ( .A(n53895), .B(n53894), .Y(u_exec_alu_p_w[24]) );
  NOR2X1 U57090 ( .A(n44539), .B(n43196), .Y(n53897) );
  NOR2X1 U57091 ( .A(n44537), .B(n43198), .Y(n53896) );
  NOR2X1 U57092 ( .A(n53897), .B(n53896), .Y(n53899) );
  NOR2X1 U57093 ( .A(n19723), .B(n19722), .Y(n53898) );
  NAND2X1 U57094 ( .A(n53899), .B(n53898), .Y(u_decode_u_regfile_N679) );
  NOR2X1 U57095 ( .A(n44603), .B(n43196), .Y(n53901) );
  NOR2X1 U57096 ( .A(n44600), .B(n43198), .Y(n53900) );
  NOR2X1 U57097 ( .A(n53901), .B(n53900), .Y(n53903) );
  NOR2X1 U57098 ( .A(n18139), .B(n18137), .Y(n53902) );
  NAND2X1 U57099 ( .A(n53903), .B(n53902), .Y(u_decode_u_regfile_N975) );
  NOR2X1 U57100 ( .A(n43194), .B(n57131), .Y(n53905) );
  NOR2X1 U57101 ( .A(n43197), .B(n43387), .Y(n53904) );
  NOR2X1 U57102 ( .A(n53905), .B(n53904), .Y(n53907) );
  NOR2X1 U57103 ( .A(n21293), .B(n21292), .Y(n53906) );
  NAND2X1 U57104 ( .A(n53907), .B(n53906), .Y(u_decode_u_regfile_N383) );
  NOR2X1 U57105 ( .A(n44474), .B(n43196), .Y(n53909) );
  NOR2X1 U57106 ( .A(n44471), .B(n43198), .Y(n53908) );
  NOR2X1 U57107 ( .A(n53909), .B(n53908), .Y(n53911) );
  NOR2X1 U57108 ( .A(n20900), .B(n20899), .Y(n53910) );
  NAND2X1 U57109 ( .A(n53911), .B(n53910), .Y(u_decode_u_regfile_N457) );
  NOR2X1 U57110 ( .A(n44561), .B(n43196), .Y(n53913) );
  NOR2X1 U57111 ( .A(n44558), .B(n43198), .Y(n53912) );
  NOR2X1 U57112 ( .A(n53913), .B(n53912), .Y(n53915) );
  NOR2X1 U57113 ( .A(n19328), .B(n19327), .Y(n53914) );
  NAND2X1 U57114 ( .A(n53915), .B(n53914), .Y(u_decode_u_regfile_N753) );
  NOR2X1 U57115 ( .A(n22425), .B(n43196), .Y(n53917) );
  NOR2X1 U57116 ( .A(n44381), .B(n37595), .Y(n53916) );
  NOR2X1 U57117 ( .A(n53917), .B(n53916), .Y(n53919) );
  NOR2X1 U57118 ( .A(n22470), .B(n22469), .Y(n53918) );
  NAND2X1 U57119 ( .A(n53919), .B(n53918), .Y(u_decode_u_regfile_N161) );
  NOR2X1 U57120 ( .A(n23761), .B(n43195), .Y(n53921) );
  NOR2X1 U57121 ( .A(n44303), .B(n37595), .Y(n53920) );
  NOR2X1 U57122 ( .A(n53921), .B(n53920), .Y(n53923) );
  NOR2X1 U57123 ( .A(n23812), .B(n23811), .Y(n53922) );
  NAND2X1 U57124 ( .A(n53923), .B(n53922), .Y(u_decode_u_regfile_N1049) );
  NOR2X1 U57125 ( .A(n44573), .B(n43195), .Y(n53925) );
  NOR2X1 U57126 ( .A(n44570), .B(n37595), .Y(n53924) );
  NOR2X1 U57127 ( .A(n53925), .B(n53924), .Y(n53927) );
  NOR2X1 U57128 ( .A(n18936), .B(n18935), .Y(n53926) );
  NAND2X1 U57129 ( .A(n53927), .B(n53926), .Y(u_decode_u_regfile_N827) );
  NOR2X1 U57130 ( .A(n43194), .B(n57209), .Y(n53929) );
  NOR2X1 U57131 ( .A(n43197), .B(n43384), .Y(n53928) );
  NOR2X1 U57132 ( .A(n53929), .B(n53928), .Y(n53931) );
  NOR2X1 U57133 ( .A(n20508), .B(n20507), .Y(n53930) );
  NAND2X1 U57134 ( .A(n53931), .B(n53930), .Y(u_decode_u_regfile_N531) );
  NOR2X1 U57135 ( .A(n22033), .B(n43195), .Y(n53933) );
  NOR2X1 U57136 ( .A(n44405), .B(n37595), .Y(n53932) );
  NOR2X1 U57137 ( .A(n53933), .B(n53932), .Y(n53935) );
  NOR2X1 U57138 ( .A(n22078), .B(n22077), .Y(n53934) );
  NAND2X1 U57139 ( .A(n53935), .B(n53934), .Y(u_decode_u_regfile_N235) );
  NOR2X1 U57140 ( .A(n23321), .B(n43195), .Y(n53937) );
  NOR2X1 U57141 ( .A(n44327), .B(n37595), .Y(n53936) );
  NOR2X1 U57142 ( .A(n53937), .B(n53936), .Y(n53939) );
  NOR2X1 U57143 ( .A(n23372), .B(n23371), .Y(n53938) );
  NAND2X1 U57144 ( .A(n53939), .B(n53938), .Y(u_decode_u_regfile_N1123) );
  NOR2X1 U57145 ( .A(n44585), .B(n43195), .Y(n53941) );
  NOR2X1 U57146 ( .A(n44582), .B(n37595), .Y(n53940) );
  NOR2X1 U57147 ( .A(n53941), .B(n53940), .Y(n53943) );
  NOR2X1 U57148 ( .A(n18544), .B(n18543), .Y(n53942) );
  NAND2X1 U57149 ( .A(n53943), .B(n53942), .Y(u_decode_u_regfile_N901) );
  NOR2X1 U57150 ( .A(n21641), .B(n43195), .Y(n53945) );
  NOR2X1 U57151 ( .A(n44429), .B(n37595), .Y(n53944) );
  NOR2X1 U57152 ( .A(n53945), .B(n53944), .Y(n53947) );
  NOR2X1 U57153 ( .A(n21686), .B(n21685), .Y(n53946) );
  NAND2X1 U57154 ( .A(n53947), .B(n53946), .Y(u_decode_u_regfile_N309) );
  NOR2X1 U57155 ( .A(n20071), .B(n43195), .Y(n53949) );
  NOR2X1 U57156 ( .A(n44513), .B(n37595), .Y(n53948) );
  NOR2X1 U57157 ( .A(n53949), .B(n53948), .Y(n53951) );
  NOR2X1 U57158 ( .A(n20116), .B(n20115), .Y(n53950) );
  NAND2X1 U57159 ( .A(n53951), .B(n53950), .Y(u_decode_u_regfile_N605) );
  NOR2X1 U57160 ( .A(n22887), .B(n43195), .Y(n53953) );
  NOR2X1 U57161 ( .A(n44351), .B(n37595), .Y(n53952) );
  NOR2X1 U57162 ( .A(n53953), .B(n53952), .Y(n53955) );
  NOR2X1 U57163 ( .A(n22938), .B(n22937), .Y(n53954) );
  NAND2X1 U57164 ( .A(n53955), .B(n53954), .Y(u_decode_u_regfile_N1197) );
  NOR2X1 U57165 ( .A(n44608), .B(n43195), .Y(n53957) );
  NOR2X1 U57166 ( .A(n44605), .B(n37595), .Y(n53956) );
  NOR2X1 U57167 ( .A(n53957), .B(n53956), .Y(n53959) );
  NOR2X1 U57168 ( .A(n24022), .B(n24021), .Y(n53958) );
  NAND2X1 U57169 ( .A(n53959), .B(n53958), .Y(u_decode_u_regfile_N1012) );
  NOR2X1 U57170 ( .A(n43194), .B(n57144), .Y(n53961) );
  NOR2X1 U57171 ( .A(n43197), .B(n43390), .Y(n53960) );
  NOR2X1 U57172 ( .A(n53961), .B(n53960), .Y(n53963) );
  NOR2X1 U57173 ( .A(n22682), .B(n22681), .Y(n53962) );
  NAND2X1 U57174 ( .A(n53963), .B(n53962), .Y(u_decode_u_regfile_N124) );
  NOR2X1 U57175 ( .A(n21051), .B(n43195), .Y(n53965) );
  NOR2X1 U57176 ( .A(n44459), .B(n37595), .Y(n53964) );
  NOR2X1 U57177 ( .A(n53965), .B(n53964), .Y(n53967) );
  NOR2X1 U57178 ( .A(n21096), .B(n21095), .Y(n53966) );
  NAND2X1 U57179 ( .A(n53967), .B(n53966), .Y(u_decode_u_regfile_N420) );
  NOR2X1 U57180 ( .A(n19481), .B(n43195), .Y(n53969) );
  NOR2X1 U57181 ( .A(n44549), .B(n37595), .Y(n53968) );
  NOR2X1 U57182 ( .A(n53969), .B(n53968), .Y(n53971) );
  NOR2X1 U57183 ( .A(n19526), .B(n19525), .Y(n53970) );
  NAND2X1 U57184 ( .A(n53971), .B(n53970), .Y(u_decode_u_regfile_N716) );
  NOR2X1 U57185 ( .A(n19088), .B(n43195), .Y(n53973) );
  NOR2X1 U57186 ( .A(n44564), .B(n43197), .Y(n53972) );
  NOR2X1 U57187 ( .A(n53973), .B(n53972), .Y(n53975) );
  NOR2X1 U57188 ( .A(n19132), .B(n19131), .Y(n53974) );
  NAND2X1 U57189 ( .A(n53975), .B(n53974), .Y(u_decode_u_regfile_N790) );
  NOR2X1 U57190 ( .A(n23541), .B(n43194), .Y(n53977) );
  NOR2X1 U57191 ( .A(n44315), .B(n43197), .Y(n53976) );
  NOR2X1 U57192 ( .A(n53977), .B(n53976), .Y(n53979) );
  NOR2X1 U57193 ( .A(n23592), .B(n23591), .Y(n53978) );
  NAND2X1 U57194 ( .A(n53979), .B(n53978), .Y(u_decode_u_regfile_N1086) );
  NOR2X1 U57195 ( .A(n22229), .B(n43194), .Y(n53981) );
  NOR2X1 U57196 ( .A(n44393), .B(n43197), .Y(n53980) );
  NOR2X1 U57197 ( .A(n53981), .B(n53980), .Y(n53983) );
  NOR2X1 U57198 ( .A(n22274), .B(n22273), .Y(n53982) );
  NAND2X1 U57199 ( .A(n53983), .B(n53982), .Y(u_decode_u_regfile_N198) );
  NOR2X1 U57200 ( .A(n20659), .B(n43194), .Y(n53985) );
  NOR2X1 U57201 ( .A(n44483), .B(n37595), .Y(n53984) );
  NOR2X1 U57202 ( .A(n53985), .B(n53984), .Y(n53987) );
  NOR2X1 U57203 ( .A(n20704), .B(n20703), .Y(n53986) );
  NAND2X1 U57204 ( .A(n53987), .B(n53986), .Y(u_decode_u_regfile_N494) );
  NOR2X1 U57205 ( .A(n21837), .B(n43194), .Y(n53989) );
  NOR2X1 U57206 ( .A(n44417), .B(n43197), .Y(n53988) );
  NOR2X1 U57207 ( .A(n53989), .B(n53988), .Y(n53991) );
  NOR2X1 U57208 ( .A(n21882), .B(n21881), .Y(n53990) );
  NAND2X1 U57209 ( .A(n53991), .B(n53990), .Y(u_decode_u_regfile_N272) );
  NOR2X1 U57210 ( .A(n23107), .B(n43194), .Y(n53993) );
  NOR2X1 U57211 ( .A(n44339), .B(n43197), .Y(n53992) );
  NOR2X1 U57212 ( .A(n53993), .B(n53992), .Y(n53995) );
  NOR2X1 U57213 ( .A(n23152), .B(n23151), .Y(n53994) );
  NAND2X1 U57214 ( .A(n53995), .B(n53994), .Y(u_decode_u_regfile_N1160) );
  NOR2X1 U57215 ( .A(n20267), .B(n43194), .Y(n53997) );
  NOR2X1 U57216 ( .A(n44501), .B(n43197), .Y(n53996) );
  NOR2X1 U57217 ( .A(n53997), .B(n53996), .Y(n53999) );
  NOR2X1 U57218 ( .A(n20312), .B(n20311), .Y(n53998) );
  NAND2X1 U57219 ( .A(n53999), .B(n53998), .Y(u_decode_u_regfile_N568) );
  NOR2X1 U57220 ( .A(n18696), .B(n43194), .Y(n54001) );
  NOR2X1 U57221 ( .A(n44576), .B(n43197), .Y(n54000) );
  NOR2X1 U57222 ( .A(n54001), .B(n54000), .Y(n54003) );
  NOR2X1 U57223 ( .A(n18740), .B(n18739), .Y(n54002) );
  NAND2X1 U57224 ( .A(n54003), .B(n54002), .Y(u_decode_u_regfile_N864) );
  NOR2X1 U57225 ( .A(n19875), .B(n43194), .Y(n54005) );
  NOR2X1 U57226 ( .A(n44525), .B(n43197), .Y(n54004) );
  NOR2X1 U57227 ( .A(n54005), .B(n54004), .Y(n54007) );
  NOR2X1 U57228 ( .A(n19920), .B(n19919), .Y(n54006) );
  NAND2X1 U57229 ( .A(n54007), .B(n54006), .Y(u_decode_u_regfile_N642) );
  NOR2X1 U57230 ( .A(n18305), .B(n43195), .Y(n54009) );
  NOR2X1 U57231 ( .A(n44591), .B(n43197), .Y(n54008) );
  NOR2X1 U57232 ( .A(n54009), .B(n54008), .Y(n54011) );
  NOR2X1 U57233 ( .A(n18350), .B(n18349), .Y(n54010) );
  NAND2X1 U57234 ( .A(n54011), .B(n54010), .Y(u_decode_u_regfile_N938) );
  NOR2X1 U57235 ( .A(n44365), .B(n43194), .Y(n54013) );
  NOR2X1 U57236 ( .A(n44362), .B(n43197), .Y(n54012) );
  NOR2X1 U57237 ( .A(n54013), .B(n54012), .Y(n54015) );
  NOR2X1 U57238 ( .A(n22718), .B(n22717), .Y(n54014) );
  NAND2X1 U57239 ( .A(n54015), .B(n54014), .Y(u_decode_u_regfile_N1234) );
  NOR2X1 U57240 ( .A(n21445), .B(n43195), .Y(n54017) );
  NOR2X1 U57241 ( .A(n44441), .B(n37595), .Y(n54016) );
  NOR2X1 U57242 ( .A(n54017), .B(n54016), .Y(n54019) );
  NOR2X1 U57243 ( .A(n21490), .B(n21489), .Y(n54018) );
  NAND2X1 U57244 ( .A(n54019), .B(n54018), .Y(u_decode_u_regfile_N346) );
  NOR2X1 U57245 ( .A(n16240), .B(n16241), .Y(n54021) );
  NOR2X1 U57246 ( .A(n16282), .B(n16283), .Y(n54020) );
  NAND2X1 U57247 ( .A(n54021), .B(n54020), .Y(u_exec_alu_p_w[25]) );
  NOR2X1 U57248 ( .A(n44539), .B(n43201), .Y(n54023) );
  NOR2X1 U57249 ( .A(n44537), .B(n43203), .Y(n54022) );
  NOR2X1 U57250 ( .A(n54023), .B(n54022), .Y(n54025) );
  NOR2X1 U57251 ( .A(n19717), .B(n19716), .Y(n54024) );
  NAND2X1 U57252 ( .A(n54025), .B(n54024), .Y(u_decode_u_regfile_N680) );
  NOR2X1 U57253 ( .A(n44603), .B(n43201), .Y(n54027) );
  NOR2X1 U57254 ( .A(n44600), .B(n43203), .Y(n54026) );
  NOR2X1 U57255 ( .A(n54027), .B(n54026), .Y(n54029) );
  NOR2X1 U57256 ( .A(n18132), .B(n18130), .Y(n54028) );
  NAND2X1 U57257 ( .A(n54029), .B(n54028), .Y(u_decode_u_regfile_N976) );
  NOR2X1 U57258 ( .A(n43199), .B(n57131), .Y(n54031) );
  NOR2X1 U57259 ( .A(n43202), .B(n43386), .Y(n54030) );
  NOR2X1 U57260 ( .A(n54031), .B(n54030), .Y(n54033) );
  NOR2X1 U57261 ( .A(n21287), .B(n21286), .Y(n54032) );
  NAND2X1 U57262 ( .A(n54033), .B(n54032), .Y(u_decode_u_regfile_N384) );
  NOR2X1 U57263 ( .A(n44474), .B(n43201), .Y(n54035) );
  NOR2X1 U57264 ( .A(n44471), .B(n43203), .Y(n54034) );
  NOR2X1 U57265 ( .A(n54035), .B(n54034), .Y(n54037) );
  NOR2X1 U57266 ( .A(n20894), .B(n20893), .Y(n54036) );
  NAND2X1 U57267 ( .A(n54037), .B(n54036), .Y(u_decode_u_regfile_N458) );
  NOR2X1 U57268 ( .A(n44561), .B(n43201), .Y(n54039) );
  NOR2X1 U57269 ( .A(n44558), .B(n43203), .Y(n54038) );
  NOR2X1 U57270 ( .A(n54039), .B(n54038), .Y(n54041) );
  NOR2X1 U57271 ( .A(n19322), .B(n19321), .Y(n54040) );
  NAND2X1 U57272 ( .A(n54041), .B(n54040), .Y(u_decode_u_regfile_N754) );
  NOR2X1 U57273 ( .A(n22425), .B(n43201), .Y(n54043) );
  NOR2X1 U57274 ( .A(n44381), .B(n37596), .Y(n54042) );
  NOR2X1 U57275 ( .A(n54043), .B(n54042), .Y(n54045) );
  NOR2X1 U57276 ( .A(n22464), .B(n22463), .Y(n54044) );
  NAND2X1 U57277 ( .A(n54045), .B(n54044), .Y(u_decode_u_regfile_N162) );
  NOR2X1 U57278 ( .A(n23761), .B(n43200), .Y(n54047) );
  NOR2X1 U57279 ( .A(n44303), .B(n37596), .Y(n54046) );
  NOR2X1 U57280 ( .A(n54047), .B(n54046), .Y(n54049) );
  NOR2X1 U57281 ( .A(n23800), .B(n23799), .Y(n54048) );
  NAND2X1 U57282 ( .A(n54049), .B(n54048), .Y(u_decode_u_regfile_N1050) );
  NOR2X1 U57283 ( .A(n44573), .B(n43200), .Y(n54051) );
  NOR2X1 U57284 ( .A(n44570), .B(n37596), .Y(n54050) );
  NOR2X1 U57285 ( .A(n54051), .B(n54050), .Y(n54053) );
  NOR2X1 U57286 ( .A(n18930), .B(n18929), .Y(n54052) );
  NAND2X1 U57287 ( .A(n54053), .B(n54052), .Y(u_decode_u_regfile_N828) );
  NOR2X1 U57288 ( .A(n43199), .B(n57209), .Y(n54055) );
  NOR2X1 U57289 ( .A(n43202), .B(n43383), .Y(n54054) );
  NOR2X1 U57290 ( .A(n54055), .B(n54054), .Y(n54057) );
  NOR2X1 U57291 ( .A(n20502), .B(n20501), .Y(n54056) );
  NAND2X1 U57292 ( .A(n54057), .B(n54056), .Y(u_decode_u_regfile_N532) );
  NOR2X1 U57293 ( .A(n22033), .B(n43200), .Y(n54059) );
  NOR2X1 U57294 ( .A(n44405), .B(n37596), .Y(n54058) );
  NOR2X1 U57295 ( .A(n54059), .B(n54058), .Y(n54061) );
  NOR2X1 U57296 ( .A(n22072), .B(n22071), .Y(n54060) );
  NAND2X1 U57297 ( .A(n54061), .B(n54060), .Y(u_decode_u_regfile_N236) );
  NOR2X1 U57298 ( .A(n23321), .B(n43200), .Y(n54063) );
  NOR2X1 U57299 ( .A(n44327), .B(n37596), .Y(n54062) );
  NOR2X1 U57300 ( .A(n54063), .B(n54062), .Y(n54065) );
  NOR2X1 U57301 ( .A(n23366), .B(n23365), .Y(n54064) );
  NAND2X1 U57302 ( .A(n54065), .B(n54064), .Y(u_decode_u_regfile_N1124) );
  NOR2X1 U57303 ( .A(n44585), .B(n43200), .Y(n54067) );
  NOR2X1 U57304 ( .A(n44582), .B(n37596), .Y(n54066) );
  NOR2X1 U57305 ( .A(n54067), .B(n54066), .Y(n54069) );
  NOR2X1 U57306 ( .A(n18538), .B(n18537), .Y(n54068) );
  NAND2X1 U57307 ( .A(n54069), .B(n54068), .Y(u_decode_u_regfile_N902) );
  NOR2X1 U57308 ( .A(n21641), .B(n43200), .Y(n54071) );
  NOR2X1 U57309 ( .A(n44429), .B(n37596), .Y(n54070) );
  NOR2X1 U57310 ( .A(n54071), .B(n54070), .Y(n54073) );
  NOR2X1 U57311 ( .A(n21680), .B(n21679), .Y(n54072) );
  NAND2X1 U57312 ( .A(n54073), .B(n54072), .Y(u_decode_u_regfile_N310) );
  NOR2X1 U57313 ( .A(n20071), .B(n43200), .Y(n54075) );
  NOR2X1 U57314 ( .A(n44513), .B(n37596), .Y(n54074) );
  NOR2X1 U57315 ( .A(n54075), .B(n54074), .Y(n54077) );
  NOR2X1 U57316 ( .A(n20110), .B(n20109), .Y(n54076) );
  NAND2X1 U57317 ( .A(n54077), .B(n54076), .Y(u_decode_u_regfile_N606) );
  NOR2X1 U57318 ( .A(n22887), .B(n43200), .Y(n54079) );
  NOR2X1 U57319 ( .A(n44351), .B(n37596), .Y(n54078) );
  NOR2X1 U57320 ( .A(n54079), .B(n54078), .Y(n54081) );
  NOR2X1 U57321 ( .A(n22932), .B(n22931), .Y(n54080) );
  NAND2X1 U57322 ( .A(n54081), .B(n54080), .Y(u_decode_u_regfile_N1198) );
  NOR2X1 U57323 ( .A(n18002), .B(n43200), .Y(n54083) );
  NOR2X1 U57324 ( .A(n44606), .B(n37596), .Y(n54082) );
  NOR2X1 U57325 ( .A(n54083), .B(n54082), .Y(n54085) );
  NOR2X1 U57326 ( .A(n24016), .B(n24015), .Y(n54084) );
  NAND2X1 U57327 ( .A(n54085), .B(n54084), .Y(u_decode_u_regfile_N1013) );
  NOR2X1 U57328 ( .A(n43199), .B(n57144), .Y(n54087) );
  NOR2X1 U57329 ( .A(n43202), .B(n43389), .Y(n54086) );
  NOR2X1 U57330 ( .A(n54087), .B(n54086), .Y(n54089) );
  NOR2X1 U57331 ( .A(n22660), .B(n22659), .Y(n54088) );
  NAND2X1 U57332 ( .A(n54089), .B(n54088), .Y(u_decode_u_regfile_N125) );
  NOR2X1 U57333 ( .A(n21051), .B(n43200), .Y(n54091) );
  NOR2X1 U57334 ( .A(n44459), .B(n37596), .Y(n54090) );
  NOR2X1 U57335 ( .A(n54091), .B(n54090), .Y(n54093) );
  NOR2X1 U57336 ( .A(n21090), .B(n21089), .Y(n54092) );
  NAND2X1 U57337 ( .A(n54093), .B(n54092), .Y(u_decode_u_regfile_N421) );
  NOR2X1 U57338 ( .A(n19481), .B(n43200), .Y(n54095) );
  NOR2X1 U57339 ( .A(n44549), .B(n37596), .Y(n54094) );
  NOR2X1 U57340 ( .A(n54095), .B(n54094), .Y(n54097) );
  NOR2X1 U57341 ( .A(n19520), .B(n19519), .Y(n54096) );
  NAND2X1 U57342 ( .A(n54097), .B(n54096), .Y(u_decode_u_regfile_N717) );
  NOR2X1 U57343 ( .A(n19088), .B(n43200), .Y(n54099) );
  NOR2X1 U57344 ( .A(n44564), .B(n43202), .Y(n54098) );
  NOR2X1 U57345 ( .A(n54099), .B(n54098), .Y(n54101) );
  NOR2X1 U57346 ( .A(n19126), .B(n19125), .Y(n54100) );
  NAND2X1 U57347 ( .A(n54101), .B(n54100), .Y(u_decode_u_regfile_N791) );
  NOR2X1 U57348 ( .A(n23541), .B(n43199), .Y(n54103) );
  NOR2X1 U57349 ( .A(n44315), .B(n43202), .Y(n54102) );
  NOR2X1 U57350 ( .A(n54103), .B(n54102), .Y(n54105) );
  NOR2X1 U57351 ( .A(n23586), .B(n23585), .Y(n54104) );
  NAND2X1 U57352 ( .A(n54105), .B(n54104), .Y(u_decode_u_regfile_N1087) );
  NOR2X1 U57353 ( .A(n22229), .B(n43199), .Y(n54107) );
  NOR2X1 U57354 ( .A(n44393), .B(n43202), .Y(n54106) );
  NOR2X1 U57355 ( .A(n54107), .B(n54106), .Y(n54109) );
  NOR2X1 U57356 ( .A(n22268), .B(n22267), .Y(n54108) );
  NAND2X1 U57357 ( .A(n54109), .B(n54108), .Y(u_decode_u_regfile_N199) );
  NOR2X1 U57358 ( .A(n20659), .B(n43199), .Y(n54111) );
  NOR2X1 U57359 ( .A(n44483), .B(n37596), .Y(n54110) );
  NOR2X1 U57360 ( .A(n54111), .B(n54110), .Y(n54113) );
  NOR2X1 U57361 ( .A(n20698), .B(n20697), .Y(n54112) );
  NAND2X1 U57362 ( .A(n54113), .B(n54112), .Y(u_decode_u_regfile_N495) );
  NOR2X1 U57363 ( .A(n21837), .B(n43199), .Y(n54115) );
  NOR2X1 U57364 ( .A(n44417), .B(n43202), .Y(n54114) );
  NOR2X1 U57365 ( .A(n54115), .B(n54114), .Y(n54117) );
  NOR2X1 U57366 ( .A(n21876), .B(n21875), .Y(n54116) );
  NAND2X1 U57367 ( .A(n54117), .B(n54116), .Y(u_decode_u_regfile_N273) );
  NOR2X1 U57368 ( .A(n23107), .B(n43199), .Y(n54119) );
  NOR2X1 U57369 ( .A(n44339), .B(n43202), .Y(n54118) );
  NOR2X1 U57370 ( .A(n54119), .B(n54118), .Y(n54121) );
  NOR2X1 U57371 ( .A(n23146), .B(n23145), .Y(n54120) );
  NAND2X1 U57372 ( .A(n54121), .B(n54120), .Y(u_decode_u_regfile_N1161) );
  NOR2X1 U57373 ( .A(n20267), .B(n43199), .Y(n54123) );
  NOR2X1 U57374 ( .A(n44501), .B(n43202), .Y(n54122) );
  NOR2X1 U57375 ( .A(n54123), .B(n54122), .Y(n54125) );
  NOR2X1 U57376 ( .A(n20306), .B(n20305), .Y(n54124) );
  NAND2X1 U57377 ( .A(n54125), .B(n54124), .Y(u_decode_u_regfile_N569) );
  NOR2X1 U57378 ( .A(n18696), .B(n43199), .Y(n54127) );
  NOR2X1 U57379 ( .A(n44576), .B(n43202), .Y(n54126) );
  NOR2X1 U57380 ( .A(n54127), .B(n54126), .Y(n54129) );
  NOR2X1 U57381 ( .A(n18734), .B(n18733), .Y(n54128) );
  NAND2X1 U57382 ( .A(n54129), .B(n54128), .Y(u_decode_u_regfile_N865) );
  NOR2X1 U57383 ( .A(n19875), .B(n43199), .Y(n54131) );
  NOR2X1 U57384 ( .A(n44525), .B(n43202), .Y(n54130) );
  NOR2X1 U57385 ( .A(n54131), .B(n54130), .Y(n54133) );
  NOR2X1 U57386 ( .A(n19914), .B(n19913), .Y(n54132) );
  NAND2X1 U57387 ( .A(n54133), .B(n54132), .Y(u_decode_u_regfile_N643) );
  NOR2X1 U57388 ( .A(n18305), .B(n43200), .Y(n54135) );
  NOR2X1 U57389 ( .A(n44591), .B(n43202), .Y(n54134) );
  NOR2X1 U57390 ( .A(n54135), .B(n54134), .Y(n54137) );
  NOR2X1 U57391 ( .A(n18344), .B(n18343), .Y(n54136) );
  NAND2X1 U57392 ( .A(n54137), .B(n54136), .Y(u_decode_u_regfile_N939) );
  NOR2X1 U57393 ( .A(n44365), .B(n43199), .Y(n54139) );
  NOR2X1 U57394 ( .A(n44362), .B(n43202), .Y(n54138) );
  NOR2X1 U57395 ( .A(n54139), .B(n54138), .Y(n54141) );
  NOR2X1 U57396 ( .A(n22712), .B(n22711), .Y(n54140) );
  NAND2X1 U57397 ( .A(n54141), .B(n54140), .Y(u_decode_u_regfile_N1235) );
  NOR2X1 U57398 ( .A(n21445), .B(n43200), .Y(n54143) );
  NOR2X1 U57399 ( .A(n44441), .B(n37596), .Y(n54142) );
  NOR2X1 U57400 ( .A(n54143), .B(n54142), .Y(n54145) );
  NOR2X1 U57401 ( .A(n21484), .B(n21483), .Y(n54144) );
  NAND2X1 U57402 ( .A(n54145), .B(n54144), .Y(u_decode_u_regfile_N347) );
  NOR2X1 U57403 ( .A(n16171), .B(n16172), .Y(n54147) );
  NOR2X1 U57404 ( .A(n16218), .B(n16219), .Y(n54146) );
  NAND2X1 U57405 ( .A(n54147), .B(n54146), .Y(u_exec_alu_p_w[26]) );
  NOR2X1 U57406 ( .A(n44539), .B(n43206), .Y(n54149) );
  NOR2X1 U57407 ( .A(n44537), .B(n43209), .Y(n54148) );
  NOR2X1 U57408 ( .A(n54149), .B(n54148), .Y(n54151) );
  NOR2X1 U57409 ( .A(n19711), .B(n19710), .Y(n54150) );
  NAND2X1 U57410 ( .A(n54151), .B(n54150), .Y(u_decode_u_regfile_N681) );
  NOR2X1 U57411 ( .A(n44603), .B(n43206), .Y(n54153) );
  NOR2X1 U57412 ( .A(n44600), .B(n43209), .Y(n54152) );
  NOR2X1 U57413 ( .A(n54153), .B(n54152), .Y(n54155) );
  NOR2X1 U57414 ( .A(n18125), .B(n18123), .Y(n54154) );
  NAND2X1 U57415 ( .A(n54155), .B(n54154), .Y(u_decode_u_regfile_N977) );
  NOR2X1 U57416 ( .A(n43204), .B(n57131), .Y(n54157) );
  NOR2X1 U57417 ( .A(n43207), .B(n43386), .Y(n54156) );
  NOR2X1 U57418 ( .A(n54157), .B(n54156), .Y(n54159) );
  NOR2X1 U57419 ( .A(n21281), .B(n21280), .Y(n54158) );
  NAND2X1 U57420 ( .A(n54159), .B(n54158), .Y(u_decode_u_regfile_N385) );
  NOR2X1 U57421 ( .A(n44474), .B(n43206), .Y(n54161) );
  NOR2X1 U57422 ( .A(n44471), .B(n43209), .Y(n54160) );
  NOR2X1 U57423 ( .A(n54161), .B(n54160), .Y(n54163) );
  NOR2X1 U57424 ( .A(n20888), .B(n20887), .Y(n54162) );
  NAND2X1 U57425 ( .A(n54163), .B(n54162), .Y(u_decode_u_regfile_N459) );
  NOR2X1 U57426 ( .A(n44561), .B(n43206), .Y(n54165) );
  NOR2X1 U57427 ( .A(n44558), .B(n43209), .Y(n54164) );
  NOR2X1 U57428 ( .A(n54165), .B(n54164), .Y(n54167) );
  NOR2X1 U57429 ( .A(n19316), .B(n19315), .Y(n54166) );
  NAND2X1 U57430 ( .A(n54167), .B(n54166), .Y(u_decode_u_regfile_N755) );
  NOR2X1 U57431 ( .A(n22425), .B(n43206), .Y(n54169) );
  NOR2X1 U57432 ( .A(n44381), .B(n43208), .Y(n54168) );
  NOR2X1 U57433 ( .A(n54169), .B(n54168), .Y(n54171) );
  NOR2X1 U57434 ( .A(n22458), .B(n22457), .Y(n54170) );
  NAND2X1 U57435 ( .A(n54171), .B(n54170), .Y(u_decode_u_regfile_N163) );
  NOR2X1 U57436 ( .A(n23761), .B(n43205), .Y(n54173) );
  NOR2X1 U57437 ( .A(n44303), .B(n43208), .Y(n54172) );
  NOR2X1 U57438 ( .A(n54173), .B(n54172), .Y(n54175) );
  NOR2X1 U57439 ( .A(n23794), .B(n23793), .Y(n54174) );
  NAND2X1 U57440 ( .A(n54175), .B(n54174), .Y(u_decode_u_regfile_N1051) );
  NOR2X1 U57441 ( .A(n44573), .B(n43205), .Y(n54177) );
  NOR2X1 U57442 ( .A(n44570), .B(n43208), .Y(n54176) );
  NOR2X1 U57443 ( .A(n54177), .B(n54176), .Y(n54179) );
  NOR2X1 U57444 ( .A(n18924), .B(n18923), .Y(n54178) );
  NAND2X1 U57445 ( .A(n54179), .B(n54178), .Y(u_decode_u_regfile_N829) );
  NOR2X1 U57446 ( .A(n43204), .B(n57209), .Y(n54181) );
  NOR2X1 U57447 ( .A(n43207), .B(n43383), .Y(n54180) );
  NOR2X1 U57448 ( .A(n54181), .B(n54180), .Y(n54183) );
  NOR2X1 U57449 ( .A(n20496), .B(n20495), .Y(n54182) );
  NAND2X1 U57450 ( .A(n54183), .B(n54182), .Y(u_decode_u_regfile_N533) );
  NOR2X1 U57451 ( .A(n22033), .B(n43205), .Y(n54185) );
  NOR2X1 U57452 ( .A(n44405), .B(n43208), .Y(n54184) );
  NOR2X1 U57453 ( .A(n54185), .B(n54184), .Y(n54187) );
  NOR2X1 U57454 ( .A(n22066), .B(n22065), .Y(n54186) );
  NAND2X1 U57455 ( .A(n54187), .B(n54186), .Y(u_decode_u_regfile_N237) );
  NOR2X1 U57456 ( .A(n23321), .B(n43205), .Y(n54189) );
  NOR2X1 U57457 ( .A(n44327), .B(n43208), .Y(n54188) );
  NOR2X1 U57458 ( .A(n54189), .B(n54188), .Y(n54191) );
  NOR2X1 U57459 ( .A(n23360), .B(n23359), .Y(n54190) );
  NAND2X1 U57460 ( .A(n54191), .B(n54190), .Y(u_decode_u_regfile_N1125) );
  NOR2X1 U57461 ( .A(n44585), .B(n43205), .Y(n54193) );
  NOR2X1 U57462 ( .A(n44582), .B(n43208), .Y(n54192) );
  NOR2X1 U57463 ( .A(n54193), .B(n54192), .Y(n54195) );
  NOR2X1 U57464 ( .A(n18532), .B(n18531), .Y(n54194) );
  NAND2X1 U57465 ( .A(n54195), .B(n54194), .Y(u_decode_u_regfile_N903) );
  NOR2X1 U57466 ( .A(n21641), .B(n43205), .Y(n54197) );
  NOR2X1 U57467 ( .A(n44429), .B(n43208), .Y(n54196) );
  NOR2X1 U57468 ( .A(n54197), .B(n54196), .Y(n54199) );
  NOR2X1 U57469 ( .A(n21674), .B(n21673), .Y(n54198) );
  NAND2X1 U57470 ( .A(n54199), .B(n54198), .Y(u_decode_u_regfile_N311) );
  NOR2X1 U57471 ( .A(n20071), .B(n43205), .Y(n54201) );
  NOR2X1 U57472 ( .A(n44513), .B(n43208), .Y(n54200) );
  NOR2X1 U57473 ( .A(n54201), .B(n54200), .Y(n54203) );
  NOR2X1 U57474 ( .A(n20104), .B(n20103), .Y(n54202) );
  NAND2X1 U57475 ( .A(n54203), .B(n54202), .Y(u_decode_u_regfile_N607) );
  NOR2X1 U57476 ( .A(n22887), .B(n43205), .Y(n54205) );
  NOR2X1 U57477 ( .A(n44351), .B(n43208), .Y(n54204) );
  NOR2X1 U57478 ( .A(n54205), .B(n54204), .Y(n54207) );
  NOR2X1 U57479 ( .A(n22926), .B(n22925), .Y(n54206) );
  NAND2X1 U57480 ( .A(n54207), .B(n54206), .Y(u_decode_u_regfile_N1199) );
  NOR2X1 U57481 ( .A(n18002), .B(n43205), .Y(n54209) );
  NOR2X1 U57482 ( .A(n44606), .B(n43208), .Y(n54208) );
  NOR2X1 U57483 ( .A(n54209), .B(n54208), .Y(n54211) );
  NOR2X1 U57484 ( .A(n24010), .B(n24009), .Y(n54210) );
  NAND2X1 U57485 ( .A(n54211), .B(n54210), .Y(u_decode_u_regfile_N1014) );
  NOR2X1 U57486 ( .A(n43204), .B(n57144), .Y(n54213) );
  NOR2X1 U57487 ( .A(n43207), .B(n43389), .Y(n54212) );
  NOR2X1 U57488 ( .A(n54213), .B(n54212), .Y(n54215) );
  NOR2X1 U57489 ( .A(n22654), .B(n22653), .Y(n54214) );
  NAND2X1 U57490 ( .A(n54215), .B(n54214), .Y(u_decode_u_regfile_N126) );
  NOR2X1 U57491 ( .A(n21051), .B(n43205), .Y(n54217) );
  NOR2X1 U57492 ( .A(n44459), .B(n43208), .Y(n54216) );
  NOR2X1 U57493 ( .A(n54217), .B(n54216), .Y(n54219) );
  NOR2X1 U57494 ( .A(n21084), .B(n21083), .Y(n54218) );
  NAND2X1 U57495 ( .A(n54219), .B(n54218), .Y(u_decode_u_regfile_N422) );
  NOR2X1 U57496 ( .A(n19481), .B(n43205), .Y(n54221) );
  NOR2X1 U57497 ( .A(n44549), .B(n43208), .Y(n54220) );
  NOR2X1 U57498 ( .A(n54221), .B(n54220), .Y(n54223) );
  NOR2X1 U57499 ( .A(n19514), .B(n19513), .Y(n54222) );
  NAND2X1 U57500 ( .A(n54223), .B(n54222), .Y(u_decode_u_regfile_N718) );
  NOR2X1 U57501 ( .A(n19088), .B(n43205), .Y(n54225) );
  NOR2X1 U57502 ( .A(n44564), .B(n43207), .Y(n54224) );
  NOR2X1 U57503 ( .A(n54225), .B(n54224), .Y(n54227) );
  NOR2X1 U57504 ( .A(n19120), .B(n19119), .Y(n54226) );
  NAND2X1 U57505 ( .A(n54227), .B(n54226), .Y(u_decode_u_regfile_N792) );
  NOR2X1 U57506 ( .A(n23541), .B(n43204), .Y(n54229) );
  NOR2X1 U57507 ( .A(n44315), .B(n43207), .Y(n54228) );
  NOR2X1 U57508 ( .A(n54229), .B(n54228), .Y(n54231) );
  NOR2X1 U57509 ( .A(n23580), .B(n23579), .Y(n54230) );
  NAND2X1 U57510 ( .A(n54231), .B(n54230), .Y(u_decode_u_regfile_N1088) );
  NOR2X1 U57511 ( .A(n22229), .B(n43204), .Y(n54233) );
  NOR2X1 U57512 ( .A(n44393), .B(n43207), .Y(n54232) );
  NOR2X1 U57513 ( .A(n54233), .B(n54232), .Y(n54235) );
  NOR2X1 U57514 ( .A(n22262), .B(n22261), .Y(n54234) );
  NAND2X1 U57515 ( .A(n54235), .B(n54234), .Y(u_decode_u_regfile_N200) );
  NOR2X1 U57516 ( .A(n20659), .B(n43204), .Y(n54237) );
  NOR2X1 U57517 ( .A(n44483), .B(n43208), .Y(n54236) );
  NOR2X1 U57518 ( .A(n54237), .B(n54236), .Y(n54239) );
  NOR2X1 U57519 ( .A(n20692), .B(n20691), .Y(n54238) );
  NAND2X1 U57520 ( .A(n54239), .B(n54238), .Y(u_decode_u_regfile_N496) );
  NOR2X1 U57521 ( .A(n21837), .B(n43204), .Y(n54241) );
  NOR2X1 U57522 ( .A(n44417), .B(n43207), .Y(n54240) );
  NOR2X1 U57523 ( .A(n54241), .B(n54240), .Y(n54243) );
  NOR2X1 U57524 ( .A(n21870), .B(n21869), .Y(n54242) );
  NAND2X1 U57525 ( .A(n54243), .B(n54242), .Y(u_decode_u_regfile_N274) );
  NOR2X1 U57526 ( .A(n23107), .B(n43204), .Y(n54245) );
  NOR2X1 U57527 ( .A(n44339), .B(n43207), .Y(n54244) );
  NOR2X1 U57528 ( .A(n54245), .B(n54244), .Y(n54247) );
  NOR2X1 U57529 ( .A(n23140), .B(n23139), .Y(n54246) );
  NAND2X1 U57530 ( .A(n54247), .B(n54246), .Y(u_decode_u_regfile_N1162) );
  NOR2X1 U57531 ( .A(n20267), .B(n43204), .Y(n54249) );
  NOR2X1 U57532 ( .A(n44501), .B(n43207), .Y(n54248) );
  NOR2X1 U57533 ( .A(n54249), .B(n54248), .Y(n54251) );
  NOR2X1 U57534 ( .A(n20300), .B(n20299), .Y(n54250) );
  NAND2X1 U57535 ( .A(n54251), .B(n54250), .Y(u_decode_u_regfile_N570) );
  NOR2X1 U57536 ( .A(n18696), .B(n43204), .Y(n54253) );
  NOR2X1 U57537 ( .A(n44576), .B(n43207), .Y(n54252) );
  NOR2X1 U57538 ( .A(n54253), .B(n54252), .Y(n54255) );
  NOR2X1 U57539 ( .A(n18728), .B(n18727), .Y(n54254) );
  NAND2X1 U57540 ( .A(n54255), .B(n54254), .Y(u_decode_u_regfile_N866) );
  NOR2X1 U57541 ( .A(n19875), .B(n43204), .Y(n54257) );
  NOR2X1 U57542 ( .A(n44525), .B(n43207), .Y(n54256) );
  NOR2X1 U57543 ( .A(n54257), .B(n54256), .Y(n54259) );
  NOR2X1 U57544 ( .A(n19908), .B(n19907), .Y(n54258) );
  NAND2X1 U57545 ( .A(n54259), .B(n54258), .Y(u_decode_u_regfile_N644) );
  NOR2X1 U57546 ( .A(n18305), .B(n43205), .Y(n54261) );
  NOR2X1 U57547 ( .A(n44591), .B(n43207), .Y(n54260) );
  NOR2X1 U57548 ( .A(n54261), .B(n54260), .Y(n54263) );
  NOR2X1 U57549 ( .A(n18338), .B(n18337), .Y(n54262) );
  NAND2X1 U57550 ( .A(n54263), .B(n54262), .Y(u_decode_u_regfile_N940) );
  NOR2X1 U57551 ( .A(n22667), .B(n43204), .Y(n54265) );
  NOR2X1 U57552 ( .A(n44363), .B(n43207), .Y(n54264) );
  NOR2X1 U57553 ( .A(n54265), .B(n54264), .Y(n54267) );
  NOR2X1 U57554 ( .A(n22706), .B(n22705), .Y(n54266) );
  NAND2X1 U57555 ( .A(n54267), .B(n54266), .Y(u_decode_u_regfile_N1236) );
  NOR2X1 U57556 ( .A(n21445), .B(n43205), .Y(n54269) );
  NOR2X1 U57557 ( .A(n44441), .B(n43208), .Y(n54268) );
  NOR2X1 U57558 ( .A(n54269), .B(n54268), .Y(n54271) );
  NOR2X1 U57559 ( .A(n21478), .B(n21477), .Y(n54270) );
  NAND2X1 U57560 ( .A(n54271), .B(n54270), .Y(u_decode_u_regfile_N348) );
  NAND2X1 U57561 ( .A(n44834), .B(n43991), .Y(n54352) );
  NAND2X1 U57562 ( .A(n43996), .B(n44845), .Y(n54350) );
  NAND2X1 U57563 ( .A(n44834), .B(n43983), .Y(n54349) );
  NAND2X1 U57564 ( .A(n43988), .B(n44845), .Y(n54347) );
  NAND2X1 U57565 ( .A(n44834), .B(n43972), .Y(n54346) );
  NAND2X1 U57566 ( .A(n43978), .B(n44845), .Y(n54344) );
  NAND2X1 U57567 ( .A(n44834), .B(n43945), .Y(n54343) );
  NAND2X1 U57568 ( .A(n43947), .B(n44845), .Y(n54341) );
  NAND2X1 U57569 ( .A(n44834), .B(n43933), .Y(n54340) );
  NAND2X1 U57570 ( .A(n43938), .B(n44845), .Y(n54338) );
  NAND2X1 U57571 ( .A(n44834), .B(n43928), .Y(n54337) );
  NAND2X1 U57572 ( .A(n43931), .B(n42850), .Y(n54335) );
  NAND2X1 U57573 ( .A(n44834), .B(n43921), .Y(n54334) );
  NAND2X1 U57574 ( .A(n43923), .B(n42850), .Y(n54332) );
  NAND2X1 U57575 ( .A(n44834), .B(n43912), .Y(n54331) );
  NAND2X1 U57576 ( .A(n43914), .B(n44845), .Y(n54329) );
  NAND2X1 U57577 ( .A(n44834), .B(n43906), .Y(n54328) );
  NAND2X1 U57578 ( .A(n43908), .B(n44845), .Y(n54326) );
  NAND2X1 U57579 ( .A(n44834), .B(n43898), .Y(n54325) );
  NAND2X1 U57580 ( .A(n43901), .B(n42850), .Y(n54323) );
  NAND2X1 U57581 ( .A(n44834), .B(n43892), .Y(n54322) );
  NAND2X1 U57582 ( .A(n43895), .B(n42850), .Y(n54320) );
  NAND2X1 U57583 ( .A(n44834), .B(n43882), .Y(n54319) );
  NAND2X1 U57584 ( .A(n43885), .B(n42850), .Y(n54317) );
  NAND2X1 U57585 ( .A(n44833), .B(n43872), .Y(n54316) );
  NAND2X1 U57586 ( .A(n43875), .B(n44843), .Y(n54314) );
  NAND2X1 U57587 ( .A(n44833), .B(n43953), .Y(n54313) );
  NAND2X1 U57588 ( .A(n43958), .B(n44843), .Y(n54311) );
  NAND2X1 U57589 ( .A(n44833), .B(n43965), .Y(n54310) );
  NAND2X1 U57590 ( .A(n43967), .B(n44844), .Y(n54308) );
  NAND2X1 U57591 ( .A(opcode_opcode_w[30]), .B(n43861), .Y(n54307) );
  NAND2X1 U57592 ( .A(n43866), .B(n57889), .Y(n54305) );
  NAND2X1 U57593 ( .A(opcode_opcode_w[29]), .B(n43853), .Y(n54304) );
  NAND2X1 U57594 ( .A(n43855), .B(n73367), .Y(n54302) );
  NAND2X1 U57595 ( .A(opcode_opcode_w[28]), .B(n44038), .Y(n54301) );
  NAND2X1 U57596 ( .A(n44040), .B(n58457), .Y(n54299) );
  NAND2X1 U57597 ( .A(opcode_opcode_w[27]), .B(n38379), .Y(n54298) );
  NAND2X1 U57598 ( .A(n38387), .B(n58818), .Y(n54296) );
  NAND2X1 U57599 ( .A(opcode_opcode_w[26]), .B(n43842), .Y(n54295) );
  NAND2X1 U57600 ( .A(n43847), .B(n73364), .Y(n54293) );
  NAND2X1 U57601 ( .A(opcode_opcode_w[25]), .B(n39937), .Y(n54292) );
  NAND2X1 U57602 ( .A(n39946), .B(n58817), .Y(n54290) );
  MX2X1 U57603 ( .A(n57436), .B(n39640), .S0(n54286), .Y(n58066) );
  INVX1 U57604 ( .A(n58066), .Y(n54272) );
  NAND2X1 U57605 ( .A(n54272), .B(n43456), .Y(n54280) );
  NAND2X1 U57606 ( .A(n58066), .B(n40627), .Y(n54278) );
  NAND2X1 U57607 ( .A(n54273), .B(n42717), .Y(n54277) );
  NAND2X1 U57608 ( .A(n38518), .B(n54274), .Y(n54275) );
  NAND2X1 U57609 ( .A(n42296), .B(n54275), .Y(n54276) );
  NAND2X1 U57610 ( .A(n54277), .B(n54276), .Y(n58065) );
  NAND2X1 U57611 ( .A(n54278), .B(n58065), .Y(n54279) );
  NAND2X1 U57612 ( .A(n54280), .B(n54279), .Y(n58088) );
  NAND2X1 U57613 ( .A(n58088), .B(n43471), .Y(n54285) );
  INVX1 U57614 ( .A(n58088), .Y(n54281) );
  NAND2X1 U57615 ( .A(n54281), .B(n43474), .Y(n54283) );
  MX2X1 U57616 ( .A(n54447), .B(n42760), .S0(n54286), .Y(n54282) );
  INVX1 U57617 ( .A(n54282), .Y(n58087) );
  NAND2X1 U57618 ( .A(n54283), .B(n58087), .Y(n54284) );
  NAND2X1 U57619 ( .A(n54285), .B(n54284), .Y(n58094) );
  NAND2X1 U57620 ( .A(n58094), .B(n43466), .Y(n54289) );
  MX2X1 U57621 ( .A(n54586), .B(n42749), .S0(n54286), .Y(n58093) );
  NOR2X1 U57622 ( .A(n43465), .B(n58094), .Y(n54287) );
  OR2X1 U57623 ( .A(n58093), .B(n54287), .Y(n54288) );
  NAND2X1 U57624 ( .A(n54289), .B(n54288), .Y(n58099) );
  NAND2X1 U57625 ( .A(n54290), .B(n58099), .Y(n54291) );
  NAND2X1 U57626 ( .A(n54292), .B(n54291), .Y(n58104) );
  NAND2X1 U57627 ( .A(n54293), .B(n58104), .Y(n54294) );
  NAND2X1 U57628 ( .A(n54295), .B(n54294), .Y(n58109) );
  NAND2X1 U57629 ( .A(n54296), .B(n58109), .Y(n54297) );
  NAND2X1 U57630 ( .A(n54298), .B(n54297), .Y(n58114) );
  NAND2X1 U57631 ( .A(n54299), .B(n58114), .Y(n54300) );
  NAND2X1 U57632 ( .A(n54301), .B(n54300), .Y(n58118) );
  NAND2X1 U57633 ( .A(n54302), .B(n58118), .Y(n54303) );
  NAND2X1 U57634 ( .A(n54304), .B(n54303), .Y(n57896) );
  NAND2X1 U57635 ( .A(n54305), .B(n57896), .Y(n54306) );
  NAND2X1 U57636 ( .A(n54307), .B(n54306), .Y(n57901) );
  NAND2X1 U57637 ( .A(n54308), .B(n57901), .Y(n54309) );
  NAND2X1 U57638 ( .A(n54310), .B(n54309), .Y(n56721) );
  NAND2X1 U57639 ( .A(n54311), .B(n56721), .Y(n54312) );
  NAND2X1 U57640 ( .A(n54313), .B(n54312), .Y(n56758) );
  NAND2X1 U57641 ( .A(n54314), .B(n56758), .Y(n54315) );
  NAND2X1 U57642 ( .A(n54316), .B(n54315), .Y(n56740) );
  NAND2X1 U57643 ( .A(n54317), .B(n56740), .Y(n54318) );
  NAND2X1 U57644 ( .A(n54319), .B(n54318), .Y(n56731) );
  NAND2X1 U57645 ( .A(n54320), .B(n56731), .Y(n54321) );
  NAND2X1 U57646 ( .A(n54322), .B(n54321), .Y(n56667) );
  NAND2X1 U57647 ( .A(n54323), .B(n56667), .Y(n54324) );
  NAND2X1 U57648 ( .A(n54325), .B(n54324), .Y(n56649) );
  NAND2X1 U57649 ( .A(n54326), .B(n56649), .Y(n54327) );
  NAND2X1 U57650 ( .A(n54328), .B(n54327), .Y(n56749) );
  NAND2X1 U57651 ( .A(n54329), .B(n56749), .Y(n54330) );
  NAND2X1 U57652 ( .A(n54331), .B(n54330), .Y(n56712) );
  NAND2X1 U57653 ( .A(n54332), .B(n56712), .Y(n54333) );
  NAND2X1 U57654 ( .A(n54334), .B(n54333), .Y(n56658) );
  NAND2X1 U57655 ( .A(n54335), .B(n56658), .Y(n54336) );
  NAND2X1 U57656 ( .A(n54337), .B(n54336), .Y(n56685) );
  NAND2X1 U57657 ( .A(n54338), .B(n56685), .Y(n54339) );
  NAND2X1 U57658 ( .A(n54340), .B(n54339), .Y(n56557) );
  NAND2X1 U57659 ( .A(n54341), .B(n56557), .Y(n54342) );
  NAND2X1 U57660 ( .A(n54343), .B(n54342), .Y(n56694) );
  NAND2X1 U57661 ( .A(n54344), .B(n56694), .Y(n54345) );
  NAND2X1 U57662 ( .A(n54346), .B(n54345), .Y(n56676) );
  NAND2X1 U57663 ( .A(n54347), .B(n56676), .Y(n54348) );
  NAND2X1 U57664 ( .A(n54349), .B(n54348), .Y(n56640) );
  NAND2X1 U57665 ( .A(n54350), .B(n56640), .Y(n54351) );
  NAND2X1 U57666 ( .A(n54352), .B(n54351), .Y(n56353) );
  INVX1 U57667 ( .A(n56353), .Y(n54354) );
  XNOR2X1 U57668 ( .A(n42852), .B(n54354), .Y(n54353) );
  NAND2X1 U57669 ( .A(n54353), .B(n43374), .Y(n54356) );
  MX2X1 U57670 ( .A(n37555), .B(n42219), .S0(n54354), .Y(n54355) );
  MX2X1 U57671 ( .A(n54356), .B(n54355), .S0(n44006), .Y(u_lsu_mem_addr_r[26])
         );
  NAND2X1 U57672 ( .A(n57895), .B(n44862), .Y(n56726) );
  NAND2X1 U57673 ( .A(n29655), .B(n56726), .Y(n17217) );
  NAND2X1 U57674 ( .A(challenge[99]), .B(n44855), .Y(n54357) );
  NAND2X1 U57675 ( .A(n54435), .B(n54357), .Y(n17307) );
  NOR2X1 U57676 ( .A(n43317), .B(n54376), .Y(net2411) );
  NAND2X1 U57677 ( .A(challenge[107]), .B(n44855), .Y(n54358) );
  NAND2X1 U57678 ( .A(n54437), .B(n54358), .Y(n17315) );
  NOR2X1 U57679 ( .A(n54383), .B(n42934), .Y(n54359) );
  NOR2X1 U57680 ( .A(n58363), .B(n58370), .Y(n54366) );
  NOR2X1 U57681 ( .A(n58338), .B(n58344), .Y(n54363) );
  NAND2X1 U57682 ( .A(opcode_pc_w[3]), .B(opcode_pc_w[2]), .Y(n54530) );
  INVX1 U57683 ( .A(n54530), .Y(n54478) );
  NAND2X1 U57684 ( .A(n54478), .B(opcode_pc_w[4]), .Y(n54609) );
  INVX1 U57685 ( .A(n54669), .Y(n54730) );
  NAND2X1 U57686 ( .A(n54730), .B(opcode_pc_w[7]), .Y(n54836) );
  INVX1 U57687 ( .A(n54836), .Y(n54832) );
  NAND2X1 U57688 ( .A(n42567), .B(opcode_pc_w[9]), .Y(n54912) );
  INVX1 U57689 ( .A(n54912), .Y(n54908) );
  NAND2X1 U57690 ( .A(n42568), .B(opcode_pc_w[11]), .Y(n55038) );
  INVX1 U57691 ( .A(n55038), .Y(n55043) );
  NAND2X1 U57692 ( .A(n55043), .B(opcode_pc_w[12]), .Y(n55059) );
  INVX1 U57693 ( .A(n55059), .Y(n55097) );
  NAND2X1 U57694 ( .A(n55097), .B(opcode_pc_w[13]), .Y(n55146) );
  INVX1 U57695 ( .A(n55146), .Y(n55150) );
  NAND2X1 U57696 ( .A(n55150), .B(opcode_pc_w[14]), .Y(n55202) );
  INVX1 U57697 ( .A(n55202), .Y(n55207) );
  NAND2X1 U57698 ( .A(n55207), .B(opcode_pc_w[15]), .Y(n55264) );
  INVX1 U57699 ( .A(n55264), .Y(n54360) );
  NAND2X1 U57700 ( .A(n54360), .B(opcode_pc_w[16]), .Y(n55324) );
  INVX1 U57701 ( .A(n55324), .Y(n54361) );
  NAND2X1 U57702 ( .A(n54361), .B(opcode_pc_w[17]), .Y(n55374) );
  INVX1 U57703 ( .A(n55374), .Y(n54362) );
  NAND2X1 U57704 ( .A(n54362), .B(opcode_pc_w[18]), .Y(n55375) );
  INVX1 U57705 ( .A(n55375), .Y(n55480) );
  NAND2X1 U57706 ( .A(n54363), .B(n55480), .Y(n55534) );
  INVX1 U57707 ( .A(n55534), .Y(n54364) );
  NAND2X1 U57708 ( .A(n54364), .B(opcode_pc_w[21]), .Y(n55585) );
  INVX1 U57709 ( .A(n55585), .Y(n54365) );
  NAND2X1 U57710 ( .A(n54365), .B(opcode_pc_w[22]), .Y(n55586) );
  INVX1 U57711 ( .A(n55586), .Y(n55683) );
  NAND2X1 U57712 ( .A(n54366), .B(n55683), .Y(n55731) );
  INVX1 U57713 ( .A(n55731), .Y(n54367) );
  NAND2X1 U57714 ( .A(n54367), .B(opcode_pc_w[25]), .Y(n55732) );
  NAND2X1 U57715 ( .A(n55732), .B(n58382), .Y(n54369) );
  INVX1 U57716 ( .A(n55732), .Y(n54368) );
  NAND2X1 U57717 ( .A(n54368), .B(opcode_pc_w[26]), .Y(n55954) );
  NAND2X1 U57718 ( .A(n54369), .B(n55954), .Y(n55779) );
  NOR2X1 U57719 ( .A(n43326), .B(n55779), .Y(n54371) );
  NOR2X1 U57720 ( .A(n54371), .B(n54370), .Y(n54380) );
  NOR2X1 U57721 ( .A(n42845), .B(n42933), .Y(n54372) );
  NOR2X1 U57722 ( .A(n2190), .B(n43320), .Y(n54378) );
  NOR2X1 U57723 ( .A(n43406), .B(n42845), .Y(n54375) );
  NOR2X1 U57724 ( .A(mem_i_valid_i), .B(u_fetch_fetch_page_fault_q), .Y(n54373) );
  NOR2X1 U57725 ( .A(n54373), .B(n42934), .Y(n54374) );
  NOR2X1 U57726 ( .A(n43323), .B(n54376), .Y(n54377) );
  NOR2X1 U57727 ( .A(n54378), .B(n54377), .Y(n54379) );
  NAND2X1 U57728 ( .A(n54380), .B(n54379), .Y(u_decode_N316) );
  NOR2X1 U57729 ( .A(n73390), .B(n54382), .Y(n54384) );
  NAND2X1 U57730 ( .A(challenge[35]), .B(n44855), .Y(n54385) );
  NAND2X1 U57731 ( .A(n54446), .B(n54385), .Y(n17243) );
  MX2X1 U57732 ( .A(n42689), .B(n40627), .S0(n73522), .Y(n25903) );
  NAND2X1 U57733 ( .A(opcode_pc_w[2]), .B(n36599), .Y(n54466) );
  NAND2X1 U57734 ( .A(n38919), .B(n54528), .Y(n54464) );
  NAND2X1 U57735 ( .A(n54466), .B(n54464), .Y(n54386) );
  XNOR2X1 U57736 ( .A(n54387), .B(n54386), .Y(n54388) );
  NOR2X1 U57737 ( .A(n43014), .B(n54388), .Y(n54392) );
  NAND2X1 U57738 ( .A(opcode_opcode_w[9]), .B(opcode_pc_w[2]), .Y(n54451) );
  NAND2X1 U57739 ( .A(n57436), .B(n54528), .Y(n54449) );
  NAND2X1 U57740 ( .A(n54451), .B(n54449), .Y(n54389) );
  XNOR2X1 U57741 ( .A(n54448), .B(n54389), .Y(n54390) );
  NOR2X1 U57742 ( .A(n54390), .B(n42872), .Y(n54391) );
  NOR2X1 U57743 ( .A(n54392), .B(n54391), .Y(n54398) );
  NAND2X1 U57744 ( .A(n54903), .B(n54396), .Y(n54397) );
  NAND2X1 U57745 ( .A(n54398), .B(n54397), .Y(n54432) );
  INVX1 U57746 ( .A(n54432), .Y(n54399) );
  NOR2X1 U57747 ( .A(n54399), .B(n57240), .Y(n54404) );
  NAND2X1 U57748 ( .A(n43286), .B(n54431), .Y(n54402) );
  NAND2X1 U57749 ( .A(n44281), .B(n25903), .Y(n54412) );
  NAND2X1 U57750 ( .A(n27560), .B(n54412), .Y(n54400) );
  NAND2X1 U57751 ( .A(u_csr_csr_mepc_q[2]), .B(n54400), .Y(n54401) );
  NAND2X1 U57752 ( .A(n54402), .B(n54401), .Y(n54403) );
  NOR2X1 U57753 ( .A(n54404), .B(n54403), .Y(n54411) );
  MX2X1 U57754 ( .A(n56578), .B(n43245), .S0(opcode_pc_w[2]), .Y(n54409) );
  INVX1 U57755 ( .A(n58222), .Y(n55540) );
  NAND2X1 U57756 ( .A(n3064), .B(n55540), .Y(n54407) );
  INVX1 U57757 ( .A(n25903), .Y(n73505) );
  NAND2X1 U57758 ( .A(n73505), .B(n42442), .Y(n58408) );
  INVX1 U57759 ( .A(n58408), .Y(n58452) );
  NAND2X1 U57760 ( .A(n58452), .B(n57247), .Y(n54406) );
  NAND2X1 U57761 ( .A(n54407), .B(n54406), .Y(n54408) );
  NOR2X1 U57762 ( .A(n54409), .B(n54408), .Y(n54410) );
  NAND2X1 U57763 ( .A(n54411), .B(n54410), .Y(u_csr_csr_mepc_r[2]) );
  NOR2X1 U57764 ( .A(n8845), .B(n57254), .Y(n54417) );
  NAND2X1 U57765 ( .A(n43289), .B(n54432), .Y(n54415) );
  NAND2X1 U57766 ( .A(n26456), .B(n54412), .Y(n54413) );
  NAND2X1 U57767 ( .A(u_csr_csr_sepc_q[2]), .B(n54413), .Y(n54414) );
  NAND2X1 U57768 ( .A(n54415), .B(n54414), .Y(n54416) );
  NOR2X1 U57769 ( .A(n54417), .B(n54416), .Y(n54424) );
  MX2X1 U57770 ( .A(n56590), .B(n43258), .S0(opcode_pc_w[2]), .Y(n54422) );
  INVX1 U57771 ( .A(n58251), .Y(n58279) );
  NAND2X1 U57772 ( .A(n3064), .B(n58279), .Y(n54420) );
  INVX1 U57773 ( .A(n58274), .Y(n55061) );
  NAND2X1 U57774 ( .A(n58452), .B(n55061), .Y(n54419) );
  NAND2X1 U57775 ( .A(n54420), .B(n54419), .Y(n54421) );
  NOR2X1 U57776 ( .A(n54422), .B(n54421), .Y(n54423) );
  NAND2X1 U57777 ( .A(n54424), .B(n54423), .Y(u_csr_csr_sepc_r[2]) );
  AND2X1 U57778 ( .A(n28494), .B(n28492), .Y(n54428) );
  NOR2X1 U57779 ( .A(n58488), .B(n43294), .Y(n54426) );
  NOR2X1 U57780 ( .A(n58487), .B(n43297), .Y(n54425) );
  NOR2X1 U57781 ( .A(n54426), .B(n54425), .Y(n54427) );
  NAND2X1 U57782 ( .A(n54428), .B(n54427), .Y(u_csr_N3667) );
  NAND2X1 U57783 ( .A(n43298), .B(n54432), .Y(n54430) );
  NAND2X1 U57784 ( .A(n43301), .B(n54431), .Y(n54429) );
  NAND2X1 U57785 ( .A(n54430), .B(n54429), .Y(net2283) );
  NOR2X1 U57786 ( .A(n2004), .B(n43304), .Y(n54433) );
  INVX1 U57787 ( .A(mem_i_pc_o[2]), .Y(n36343) );
  NAND2X1 U57788 ( .A(challenge[98]), .B(n44854), .Y(n54434) );
  NAND2X1 U57789 ( .A(n54435), .B(n54434), .Y(n17306) );
  NOR2X1 U57790 ( .A(n43317), .B(n54440), .Y(net2382) );
  NAND2X1 U57791 ( .A(challenge[106]), .B(n44854), .Y(n54436) );
  NAND2X1 U57792 ( .A(n54437), .B(n54436), .Y(n17314) );
  NOR2X1 U57793 ( .A(n2005), .B(n43320), .Y(n54439) );
  NOR2X1 U57794 ( .A(n54439), .B(n54438), .Y(n54444) );
  NOR2X1 U57795 ( .A(n43323), .B(n54440), .Y(n54442) );
  NOR2X1 U57796 ( .A(opcode_pc_w[2]), .B(n43328), .Y(n54441) );
  NOR2X1 U57797 ( .A(n54442), .B(n54441), .Y(n54443) );
  NAND2X1 U57798 ( .A(n54444), .B(n54443), .Y(u_decode_N292) );
  NAND2X1 U57799 ( .A(challenge[34]), .B(n44854), .Y(n54445) );
  NAND2X1 U57800 ( .A(n54446), .B(n54445), .Y(n17242) );
  MX2X1 U57801 ( .A(n42788), .B(n43470), .S0(n73522), .Y(n25860) );
  NAND2X1 U57802 ( .A(n43286), .B(n54571), .Y(n54477) );
  NAND2X1 U57803 ( .A(opcode_pc_w[3]), .B(opcode_opcode_w[10]), .Y(n54455) );
  NAND2X1 U57804 ( .A(n54447), .B(n54529), .Y(n54453) );
  INVX1 U57805 ( .A(n54448), .Y(n54450) );
  NAND2X1 U57806 ( .A(n54450), .B(n54449), .Y(n54452) );
  NAND2X1 U57807 ( .A(n54452), .B(n54451), .Y(n54511) );
  NAND2X1 U57808 ( .A(n54453), .B(n54511), .Y(n54454) );
  NAND2X1 U57809 ( .A(n54455), .B(n54454), .Y(n54587) );
  NOR2X1 U57810 ( .A(n54456), .B(n42873), .Y(n54463) );
  XNOR2X1 U57811 ( .A(n54458), .B(n54457), .Y(n54459) );
  XOR2X1 U57812 ( .A(n54460), .B(n54459), .Y(n54461) );
  NOR2X1 U57813 ( .A(n54461), .B(n42931), .Y(n54462) );
  NOR2X1 U57814 ( .A(n54463), .B(n54462), .Y(n54475) );
  NAND2X1 U57815 ( .A(opcode_pc_w[3]), .B(n40454), .Y(n54470) );
  NAND2X1 U57816 ( .A(n42760), .B(n54529), .Y(n54468) );
  NAND2X1 U57817 ( .A(n54465), .B(n54464), .Y(n54467) );
  NAND2X1 U57818 ( .A(n54467), .B(n54466), .Y(n54520) );
  NAND2X1 U57819 ( .A(n54468), .B(n54520), .Y(n54469) );
  NAND2X1 U57820 ( .A(n54470), .B(n54469), .Y(n54592) );
  INVX1 U57821 ( .A(n54592), .Y(n54472) );
  XNOR2X1 U57822 ( .A(n42747), .B(opcode_pc_w[4]), .Y(n54471) );
  XOR2X1 U57823 ( .A(n54472), .B(n54471), .Y(n54473) );
  NAND2X1 U57824 ( .A(n54473), .B(n54979), .Y(n54474) );
  NAND2X1 U57825 ( .A(n54475), .B(n54474), .Y(n54572) );
  NAND2X1 U57826 ( .A(n43246), .B(n54572), .Y(n54476) );
  NAND2X1 U57827 ( .A(n54477), .B(n54476), .Y(n54483) );
  XNOR2X1 U57828 ( .A(opcode_pc_w[4]), .B(n54478), .Y(n54578) );
  INVX1 U57829 ( .A(n54578), .Y(n54490) );
  NAND2X1 U57830 ( .A(n54490), .B(n43240), .Y(n54481) );
  NAND2X1 U57831 ( .A(n44281), .B(n25860), .Y(n54493) );
  NAND2X1 U57832 ( .A(n27560), .B(n54493), .Y(n54479) );
  NAND2X1 U57833 ( .A(u_csr_csr_mepc_q[4]), .B(n54479), .Y(n54480) );
  NAND2X1 U57834 ( .A(n54481), .B(n54480), .Y(n54482) );
  NOR2X1 U57835 ( .A(n54483), .B(n54482), .Y(n54489) );
  NOR2X1 U57836 ( .A(n42953), .B(n37763), .Y(n54487) );
  INVX1 U57837 ( .A(n25860), .Y(n73504) );
  NAND2X1 U57838 ( .A(n73504), .B(n42442), .Y(n58424) );
  INVX1 U57839 ( .A(n58424), .Y(n58454) );
  NAND2X1 U57840 ( .A(n58454), .B(n57247), .Y(n54485) );
  NAND2X1 U57841 ( .A(n43245), .B(opcode_pc_w[4]), .Y(n54484) );
  NAND2X1 U57842 ( .A(n54485), .B(n54484), .Y(n54486) );
  NOR2X1 U57843 ( .A(n54487), .B(n54486), .Y(n54488) );
  NAND2X1 U57844 ( .A(n54489), .B(n54488), .Y(u_csr_csr_mepc_r[4]) );
  INVX1 U57845 ( .A(n57254), .Y(n56600) );
  NAND2X1 U57846 ( .A(n43259), .B(n54571), .Y(n54492) );
  NAND2X1 U57847 ( .A(n54490), .B(n43250), .Y(n54491) );
  NAND2X1 U57848 ( .A(n54492), .B(n54491), .Y(n54498) );
  NAND2X1 U57849 ( .A(n43289), .B(n54572), .Y(n54496) );
  NAND2X1 U57850 ( .A(n26456), .B(n54493), .Y(n54494) );
  NAND2X1 U57851 ( .A(u_csr_csr_sepc_q[4]), .B(n54494), .Y(n54495) );
  NAND2X1 U57852 ( .A(n54496), .B(n54495), .Y(n54497) );
  NOR2X1 U57853 ( .A(n54498), .B(n54497), .Y(n54504) );
  NOR2X1 U57854 ( .A(n42957), .B(n37763), .Y(n54502) );
  NAND2X1 U57855 ( .A(n58454), .B(n55061), .Y(n54500) );
  NAND2X1 U57856 ( .A(n43258), .B(opcode_pc_w[4]), .Y(n54499) );
  NAND2X1 U57857 ( .A(n54500), .B(n54499), .Y(n54501) );
  NOR2X1 U57858 ( .A(n54502), .B(n54501), .Y(n54503) );
  NAND2X1 U57859 ( .A(n54504), .B(n54503), .Y(u_csr_csr_sepc_r[4]) );
  AND2X1 U57860 ( .A(n28478), .B(n28476), .Y(n54508) );
  NOR2X1 U57861 ( .A(n58494), .B(n43294), .Y(n54506) );
  NOR2X1 U57862 ( .A(n58493), .B(n43297), .Y(n54505) );
  NOR2X1 U57863 ( .A(n54506), .B(n54505), .Y(n54507) );
  NAND2X1 U57864 ( .A(n54508), .B(n54507), .Y(u_csr_N3669) );
  NAND2X1 U57865 ( .A(n43298), .B(n54572), .Y(n54510) );
  NAND2X1 U57866 ( .A(n43301), .B(n54571), .Y(n54509) );
  NAND2X1 U57867 ( .A(n54510), .B(n54509), .Y(net2285) );
  MX2X1 U57868 ( .A(n42663), .B(n43476), .S0(n73522), .Y(n25872) );
  NAND2X1 U57869 ( .A(n44281), .B(n25872), .Y(n26297) );
  NOR2X1 U57870 ( .A(n54512), .B(n42874), .Y(n54519) );
  XNOR2X1 U57871 ( .A(n54514), .B(n54513), .Y(n54515) );
  XOR2X1 U57872 ( .A(n54516), .B(n54515), .Y(n54517) );
  NOR2X1 U57873 ( .A(n54517), .B(n42930), .Y(n54518) );
  NOR2X1 U57874 ( .A(n54519), .B(n54518), .Y(n54525) );
  INVX1 U57875 ( .A(n54520), .Y(n54522) );
  XNOR2X1 U57876 ( .A(n42759), .B(opcode_pc_w[3]), .Y(n54521) );
  XOR2X1 U57877 ( .A(n54522), .B(n54521), .Y(n54523) );
  NAND2X1 U57878 ( .A(n54523), .B(n54979), .Y(n54524) );
  NAND2X1 U57879 ( .A(n54525), .B(n54524), .Y(n54565) );
  NAND2X1 U57880 ( .A(n43246), .B(n54565), .Y(n54527) );
  NAND2X1 U57881 ( .A(n43286), .B(n54564), .Y(n54526) );
  NAND2X1 U57882 ( .A(n54527), .B(n54526), .Y(n54536) );
  NAND2X1 U57883 ( .A(n54529), .B(n54528), .Y(n54531) );
  NAND2X1 U57884 ( .A(n54531), .B(n54530), .Y(n56790) );
  INVX1 U57885 ( .A(n56790), .Y(n54544) );
  NAND2X1 U57886 ( .A(n54544), .B(n43240), .Y(n54534) );
  NAND2X1 U57887 ( .A(n27560), .B(n26297), .Y(n54532) );
  NAND2X1 U57888 ( .A(u_csr_csr_mepc_q[3]), .B(n54532), .Y(n54533) );
  NAND2X1 U57889 ( .A(n54534), .B(n54533), .Y(n54535) );
  NOR2X1 U57890 ( .A(n54536), .B(n54535), .Y(n54543) );
  NOR2X1 U57891 ( .A(n42953), .B(n37764), .Y(n54541) );
  INVX1 U57892 ( .A(n25872), .Y(n54537) );
  NAND2X1 U57893 ( .A(n54537), .B(n42442), .Y(n58423) );
  INVX1 U57894 ( .A(n58423), .Y(n58453) );
  NAND2X1 U57895 ( .A(n58453), .B(n57247), .Y(n54539) );
  NAND2X1 U57896 ( .A(n43245), .B(opcode_pc_w[3]), .Y(n54538) );
  NAND2X1 U57897 ( .A(n54539), .B(n54538), .Y(n54540) );
  NOR2X1 U57898 ( .A(n54541), .B(n54540), .Y(n54542) );
  NAND2X1 U57899 ( .A(n54543), .B(n54542), .Y(u_csr_csr_mepc_r[3]) );
  NAND2X1 U57900 ( .A(n43259), .B(n54564), .Y(n54546) );
  NAND2X1 U57901 ( .A(n54544), .B(n43250), .Y(n54545) );
  NAND2X1 U57902 ( .A(n54546), .B(n54545), .Y(n54551) );
  NAND2X1 U57903 ( .A(n43289), .B(n54565), .Y(n54549) );
  NAND2X1 U57904 ( .A(n26456), .B(n26297), .Y(n54547) );
  NAND2X1 U57905 ( .A(u_csr_csr_sepc_q[3]), .B(n54547), .Y(n54548) );
  NAND2X1 U57906 ( .A(n54549), .B(n54548), .Y(n54550) );
  NOR2X1 U57907 ( .A(n54551), .B(n54550), .Y(n54557) );
  NOR2X1 U57908 ( .A(n42957), .B(n37764), .Y(n54555) );
  NAND2X1 U57909 ( .A(n58453), .B(n55061), .Y(n54553) );
  NAND2X1 U57910 ( .A(n43258), .B(opcode_pc_w[3]), .Y(n54552) );
  NAND2X1 U57911 ( .A(n54553), .B(n54552), .Y(n54554) );
  NOR2X1 U57912 ( .A(n54555), .B(n54554), .Y(n54556) );
  NAND2X1 U57913 ( .A(n54557), .B(n54556), .Y(u_csr_csr_sepc_r[3]) );
  AND2X1 U57914 ( .A(n28486), .B(n28484), .Y(n54561) );
  NOR2X1 U57915 ( .A(n58492), .B(n43294), .Y(n54559) );
  NOR2X1 U57916 ( .A(n58491), .B(n43297), .Y(n54558) );
  NOR2X1 U57917 ( .A(n54559), .B(n54558), .Y(n54560) );
  NAND2X1 U57918 ( .A(n54561), .B(n54560), .Y(u_csr_N3668) );
  NAND2X1 U57919 ( .A(n43298), .B(n54565), .Y(n54563) );
  NAND2X1 U57920 ( .A(n43301), .B(n54564), .Y(n54562) );
  NAND2X1 U57921 ( .A(n54563), .B(n54562), .Y(net2284) );
  NOR2X1 U57922 ( .A(n2035), .B(n43304), .Y(n54568) );
  NAND2X1 U57923 ( .A(n43307), .B(n54564), .Y(n54567) );
  NAND2X1 U57924 ( .A(n43312), .B(n54565), .Y(n54566) );
  NAND2X1 U57925 ( .A(n54567), .B(n54566), .Y(n56787) );
  NOR2X1 U57926 ( .A(n54568), .B(n56787), .Y(n54570) );
  OR2X1 U57927 ( .A(n1761), .B(n42847), .Y(n54569) );
  NAND2X1 U57928 ( .A(n54570), .B(n54569), .Y(mem_i_pc_o[3]) );
  NOR2X1 U57929 ( .A(n2066), .B(n43304), .Y(n54575) );
  NAND2X1 U57930 ( .A(n43307), .B(n54571), .Y(n54574) );
  NAND2X1 U57931 ( .A(n43312), .B(n54572), .Y(n54573) );
  NAND2X1 U57932 ( .A(n54574), .B(n54573), .Y(n54579) );
  NOR2X1 U57933 ( .A(n54575), .B(n54579), .Y(n54577) );
  OR2X1 U57934 ( .A(n1762), .B(n42846), .Y(n54576) );
  NAND2X1 U57935 ( .A(n54577), .B(n54576), .Y(mem_i_pc_o[4]) );
  NOR2X1 U57936 ( .A(n43317), .B(n54581), .Y(net2384) );
  NOR2X1 U57937 ( .A(n43328), .B(n54578), .Y(n54580) );
  NOR2X1 U57938 ( .A(n54580), .B(n54579), .Y(n54585) );
  NOR2X1 U57939 ( .A(n2067), .B(n43320), .Y(n54583) );
  NOR2X1 U57940 ( .A(n43323), .B(n54581), .Y(n54582) );
  NOR2X1 U57941 ( .A(n54583), .B(n54582), .Y(n54584) );
  NAND2X1 U57942 ( .A(n54585), .B(n54584), .Y(u_decode_N294) );
  NAND2X1 U57943 ( .A(opcode_pc_w[4]), .B(opcode_opcode_w[11]), .Y(n54590) );
  NAND2X1 U57944 ( .A(n54586), .B(n54591), .Y(n54588) );
  NAND2X1 U57945 ( .A(n54588), .B(n54587), .Y(n54589) );
  NAND2X1 U57946 ( .A(n54590), .B(n54589), .Y(n29776) );
  NAND2X1 U57947 ( .A(opcode_pc_w[4]), .B(n42748), .Y(n54595) );
  NAND2X1 U57948 ( .A(n42749), .B(n54591), .Y(n54593) );
  NAND2X1 U57949 ( .A(n54593), .B(n54592), .Y(n54594) );
  NAND2X1 U57950 ( .A(n54595), .B(n54594), .Y(n29786) );
  NAND2X1 U57951 ( .A(n42136), .B(n39940), .Y(n54608) );
  XOR2X1 U57952 ( .A(n29777), .B(n29776), .Y(n54596) );
  NOR2X1 U57953 ( .A(n42872), .B(n54596), .Y(n54603) );
  XNOR2X1 U57954 ( .A(n54598), .B(n54597), .Y(n54599) );
  XOR2X1 U57955 ( .A(n54600), .B(n54599), .Y(n54601) );
  NOR2X1 U57956 ( .A(n54601), .B(n42931), .Y(n54602) );
  NOR2X1 U57957 ( .A(n54603), .B(n54602), .Y(n54606) );
  XNOR2X1 U57958 ( .A(n29786), .B(n29777), .Y(n54604) );
  NAND2X1 U57959 ( .A(n54604), .B(n54979), .Y(n54605) );
  NAND2X1 U57960 ( .A(n54606), .B(n54605), .Y(n54643) );
  NAND2X1 U57961 ( .A(n43246), .B(n54643), .Y(n54607) );
  NAND2X1 U57962 ( .A(n54608), .B(n54607), .Y(n54615) );
  NAND2X1 U57963 ( .A(n54609), .B(n58426), .Y(n54610) );
  NAND2X1 U57964 ( .A(n54610), .B(n54668), .Y(n54649) );
  INVX1 U57965 ( .A(n54649), .Y(n54622) );
  NAND2X1 U57966 ( .A(n54622), .B(n43240), .Y(n54613) );
  NAND2X1 U57967 ( .A(n44281), .B(n39946), .Y(n58268) );
  NAND2X1 U57968 ( .A(n27477), .B(n58268), .Y(n54611) );
  NAND2X1 U57969 ( .A(u_csr_csr_mepc_q[5]), .B(n54611), .Y(n54612) );
  NAND2X1 U57970 ( .A(n54613), .B(n54612), .Y(n54614) );
  NOR2X1 U57971 ( .A(n54615), .B(n54614), .Y(n54621) );
  NOR2X1 U57972 ( .A(n42951), .B(n37765), .Y(n54619) );
  NAND2X1 U57973 ( .A(n43245), .B(opcode_pc_w[5]), .Y(n54617) );
  NAND2X1 U57974 ( .A(n43286), .B(n54642), .Y(n54616) );
  NAND2X1 U57975 ( .A(n54617), .B(n54616), .Y(n54618) );
  NOR2X1 U57976 ( .A(n54619), .B(n54618), .Y(n54620) );
  NAND2X1 U57977 ( .A(n54621), .B(n54620), .Y(u_csr_csr_mepc_r[5]) );
  NAND2X1 U57978 ( .A(n42137), .B(n39941), .Y(n54624) );
  NAND2X1 U57979 ( .A(n54622), .B(n43250), .Y(n54623) );
  NAND2X1 U57980 ( .A(n54624), .B(n54623), .Y(n54629) );
  NAND2X1 U57981 ( .A(n43289), .B(n54643), .Y(n54627) );
  NAND2X1 U57982 ( .A(n26373), .B(n58268), .Y(n54625) );
  NAND2X1 U57983 ( .A(u_csr_csr_sepc_q[5]), .B(n54625), .Y(n54626) );
  NAND2X1 U57984 ( .A(n54627), .B(n54626), .Y(n54628) );
  NOR2X1 U57985 ( .A(n54629), .B(n54628), .Y(n54635) );
  NOR2X1 U57986 ( .A(n42956), .B(n37765), .Y(n54633) );
  NAND2X1 U57987 ( .A(n43258), .B(opcode_pc_w[5]), .Y(n54631) );
  NAND2X1 U57988 ( .A(n43259), .B(n54642), .Y(n54630) );
  NAND2X1 U57989 ( .A(n54631), .B(n54630), .Y(n54632) );
  NOR2X1 U57990 ( .A(n54633), .B(n54632), .Y(n54634) );
  NAND2X1 U57991 ( .A(n54635), .B(n54634), .Y(u_csr_csr_sepc_r[5]) );
  AND2X1 U57992 ( .A(n28470), .B(n28468), .Y(n54639) );
  NOR2X1 U57993 ( .A(n58496), .B(n43294), .Y(n54637) );
  NOR2X1 U57994 ( .A(n58495), .B(n43297), .Y(n54636) );
  NOR2X1 U57995 ( .A(n54637), .B(n54636), .Y(n54638) );
  NAND2X1 U57996 ( .A(n54639), .B(n54638), .Y(u_csr_N3670) );
  NAND2X1 U57997 ( .A(n43298), .B(n54643), .Y(n54641) );
  NAND2X1 U57998 ( .A(n43301), .B(n54642), .Y(n54640) );
  NAND2X1 U57999 ( .A(n54641), .B(n54640), .Y(net2286) );
  NOR2X1 U58000 ( .A(n2098), .B(n43306), .Y(n54646) );
  NAND2X1 U58001 ( .A(n43307), .B(n54642), .Y(n54645) );
  NAND2X1 U58002 ( .A(n43311), .B(n54643), .Y(n54644) );
  NAND2X1 U58003 ( .A(n54645), .B(n54644), .Y(n54650) );
  NOR2X1 U58004 ( .A(n54646), .B(n54650), .Y(n54648) );
  OR2X1 U58005 ( .A(n1763), .B(n42847), .Y(n54647) );
  NAND2X1 U58006 ( .A(n54648), .B(n54647), .Y(mem_i_pc_o[5]) );
  INVX1 U58007 ( .A(mem_i_pc_o[5]), .Y(n54710) );
  NAND2X1 U58008 ( .A(n42401), .B(mem_i_pc_o[4]), .Y(n54769) );
  NOR2X1 U58009 ( .A(n43317), .B(n54652), .Y(net2385) );
  NOR2X1 U58010 ( .A(n43328), .B(n54649), .Y(n54651) );
  NOR2X1 U58011 ( .A(n54651), .B(n54650), .Y(n54656) );
  NOR2X1 U58012 ( .A(n2099), .B(n43320), .Y(n54654) );
  NOR2X1 U58013 ( .A(n43323), .B(n54652), .Y(n54653) );
  NOR2X1 U58014 ( .A(n54654), .B(n54653), .Y(n54655) );
  NAND2X1 U58015 ( .A(n54656), .B(n54655), .Y(u_decode_N295) );
  NAND2X1 U58016 ( .A(n43236), .B(n43843), .Y(n54667) );
  NOR2X1 U58017 ( .A(n29764), .B(n37342), .Y(n54665) );
  NAND2X1 U58018 ( .A(n29754), .B(n54897), .Y(n54663) );
  XNOR2X1 U58019 ( .A(n54660), .B(n54659), .Y(n54661) );
  NAND2X1 U58020 ( .A(n54903), .B(n54661), .Y(n54662) );
  NAND2X1 U58021 ( .A(n54663), .B(n54662), .Y(n54664) );
  OR2X1 U58022 ( .A(n54665), .B(n54664), .Y(n54704) );
  NAND2X1 U58023 ( .A(n43246), .B(n54704), .Y(n54666) );
  NAND2X1 U58024 ( .A(n54667), .B(n54666), .Y(n54675) );
  NAND2X1 U58025 ( .A(n54668), .B(n58431), .Y(n54670) );
  NAND2X1 U58026 ( .A(n54670), .B(n54669), .Y(n54712) );
  INVX1 U58027 ( .A(n54712), .Y(n54684) );
  NAND2X1 U58028 ( .A(n54684), .B(n43240), .Y(n54673) );
  NAND2X1 U58029 ( .A(n44281), .B(n43847), .Y(n54685) );
  NAND2X1 U58030 ( .A(n27477), .B(n54685), .Y(n54671) );
  NAND2X1 U58031 ( .A(u_csr_csr_mepc_q[6]), .B(n54671), .Y(n54672) );
  NAND2X1 U58032 ( .A(n54673), .B(n54672), .Y(n54674) );
  NOR2X1 U58033 ( .A(n54675), .B(n54674), .Y(n54681) );
  NOR2X1 U58034 ( .A(n42951), .B(n37766), .Y(n54679) );
  NAND2X1 U58035 ( .A(n43245), .B(opcode_pc_w[6]), .Y(n54677) );
  NAND2X1 U58036 ( .A(n43286), .B(n54703), .Y(n54676) );
  NAND2X1 U58037 ( .A(n54677), .B(n54676), .Y(n54678) );
  NOR2X1 U58038 ( .A(n54679), .B(n54678), .Y(n54680) );
  NAND2X1 U58039 ( .A(n54681), .B(n54680), .Y(u_csr_csr_mepc_r[6]) );
  NAND2X1 U58040 ( .A(n43253), .B(n43843), .Y(n54683) );
  NAND2X1 U58041 ( .A(n43289), .B(n54704), .Y(n54682) );
  NAND2X1 U58042 ( .A(n54683), .B(n54682), .Y(n54690) );
  NAND2X1 U58043 ( .A(n54684), .B(n43250), .Y(n54688) );
  NAND2X1 U58044 ( .A(n26373), .B(n54685), .Y(n54686) );
  NAND2X1 U58045 ( .A(u_csr_csr_sepc_q[6]), .B(n54686), .Y(n54687) );
  NAND2X1 U58046 ( .A(n54688), .B(n54687), .Y(n54689) );
  NOR2X1 U58047 ( .A(n54690), .B(n54689), .Y(n54696) );
  NOR2X1 U58048 ( .A(n42957), .B(n37766), .Y(n54694) );
  NAND2X1 U58049 ( .A(n43258), .B(opcode_pc_w[6]), .Y(n54692) );
  NAND2X1 U58050 ( .A(n43259), .B(n54703), .Y(n54691) );
  NAND2X1 U58051 ( .A(n54692), .B(n54691), .Y(n54693) );
  NOR2X1 U58052 ( .A(n54694), .B(n54693), .Y(n54695) );
  NAND2X1 U58053 ( .A(n54696), .B(n54695), .Y(u_csr_csr_sepc_r[6]) );
  AND2X1 U58054 ( .A(n28462), .B(n28460), .Y(n54700) );
  NOR2X1 U58055 ( .A(n58498), .B(n43293), .Y(n54698) );
  NOR2X1 U58056 ( .A(n58497), .B(n43296), .Y(n54697) );
  NOR2X1 U58057 ( .A(n54698), .B(n54697), .Y(n54699) );
  NAND2X1 U58058 ( .A(n54700), .B(n54699), .Y(u_csr_N3671) );
  NAND2X1 U58059 ( .A(n43298), .B(n54704), .Y(n54702) );
  NAND2X1 U58060 ( .A(n43301), .B(n54703), .Y(n54701) );
  NAND2X1 U58061 ( .A(n54702), .B(n54701), .Y(net2287) );
  NOR2X1 U58062 ( .A(n2130), .B(n43304), .Y(n54707) );
  NAND2X1 U58063 ( .A(n43307), .B(n54703), .Y(n54706) );
  NAND2X1 U58064 ( .A(n43312), .B(n54704), .Y(n54705) );
  NAND2X1 U58065 ( .A(n54706), .B(n54705), .Y(n54713) );
  OR2X1 U58066 ( .A(n1764), .B(n42847), .Y(n54708) );
  NAND2X1 U58067 ( .A(n54709), .B(n54708), .Y(mem_i_pc_o[6]) );
  INVX1 U58068 ( .A(mem_i_pc_o[6]), .Y(n54770) );
  NOR2X1 U58069 ( .A(n54710), .B(n54769), .Y(n54711) );
  XNOR2X1 U58070 ( .A(n54770), .B(n54711), .Y(u_fetch_N55) );
  NOR2X1 U58071 ( .A(n43317), .B(n54715), .Y(net2386) );
  NOR2X1 U58072 ( .A(n43328), .B(n54712), .Y(n54714) );
  NOR2X1 U58073 ( .A(n54714), .B(n54713), .Y(n54719) );
  NOR2X1 U58074 ( .A(n2131), .B(n43320), .Y(n54717) );
  NOR2X1 U58075 ( .A(n43323), .B(n54715), .Y(n54716) );
  NOR2X1 U58076 ( .A(n54717), .B(n54716), .Y(n54718) );
  NAND2X1 U58077 ( .A(n54719), .B(n54718), .Y(u_decode_N296) );
  NAND2X1 U58078 ( .A(n42136), .B(n38381), .Y(n54729) );
  NOR2X1 U58079 ( .A(n29743), .B(n43014), .Y(n54727) );
  NAND2X1 U58080 ( .A(n29733), .B(n54897), .Y(n54725) );
  XNOR2X1 U58081 ( .A(n37893), .B(n54722), .Y(n54723) );
  NAND2X1 U58082 ( .A(n54903), .B(n54723), .Y(n54724) );
  NAND2X1 U58083 ( .A(n54725), .B(n54724), .Y(n54726) );
  OR2X1 U58084 ( .A(n54727), .B(n54726), .Y(n54763) );
  NAND2X1 U58085 ( .A(n43246), .B(n54763), .Y(n54728) );
  NAND2X1 U58086 ( .A(n54729), .B(n54728), .Y(n54735) );
  XNOR2X1 U58087 ( .A(opcode_pc_w[7]), .B(n54730), .Y(n54772) );
  INVX1 U58088 ( .A(n54772), .Y(n54742) );
  NAND2X1 U58089 ( .A(n54742), .B(n43240), .Y(n54733) );
  NAND2X1 U58090 ( .A(n44281), .B(n38385), .Y(n58269) );
  NAND2X1 U58091 ( .A(n27477), .B(n58269), .Y(n54731) );
  NAND2X1 U58092 ( .A(u_csr_csr_mepc_q[7]), .B(n54731), .Y(n54732) );
  NAND2X1 U58093 ( .A(n54733), .B(n54732), .Y(n54734) );
  NOR2X1 U58094 ( .A(n54735), .B(n54734), .Y(n54741) );
  NOR2X1 U58095 ( .A(n42953), .B(n37767), .Y(n54739) );
  NAND2X1 U58096 ( .A(n43245), .B(opcode_pc_w[7]), .Y(n54737) );
  NAND2X1 U58097 ( .A(n43286), .B(n54762), .Y(n54736) );
  NAND2X1 U58098 ( .A(n54737), .B(n54736), .Y(n54738) );
  NOR2X1 U58099 ( .A(n54739), .B(n54738), .Y(n54740) );
  NAND2X1 U58100 ( .A(n54741), .B(n54740), .Y(u_csr_csr_mepc_r[7]) );
  NAND2X1 U58101 ( .A(n42137), .B(n38380), .Y(n54744) );
  NAND2X1 U58102 ( .A(n54742), .B(n43250), .Y(n54743) );
  NAND2X1 U58103 ( .A(n54744), .B(n54743), .Y(n54749) );
  NAND2X1 U58104 ( .A(n43289), .B(n54763), .Y(n54747) );
  NAND2X1 U58105 ( .A(n26373), .B(n58269), .Y(n54745) );
  NAND2X1 U58106 ( .A(u_csr_csr_sepc_q[7]), .B(n54745), .Y(n54746) );
  NAND2X1 U58107 ( .A(n54747), .B(n54746), .Y(n54748) );
  NOR2X1 U58108 ( .A(n54749), .B(n54748), .Y(n54755) );
  NOR2X1 U58109 ( .A(n42957), .B(n37767), .Y(n54753) );
  NAND2X1 U58110 ( .A(n43258), .B(opcode_pc_w[7]), .Y(n54751) );
  NAND2X1 U58111 ( .A(n43259), .B(n54762), .Y(n54750) );
  NAND2X1 U58112 ( .A(n54751), .B(n54750), .Y(n54752) );
  NOR2X1 U58113 ( .A(n54753), .B(n54752), .Y(n54754) );
  NAND2X1 U58114 ( .A(n54755), .B(n54754), .Y(u_csr_csr_sepc_r[7]) );
  AND2X1 U58115 ( .A(n28454), .B(n28452), .Y(n54759) );
  NOR2X1 U58116 ( .A(n58500), .B(n43293), .Y(n54757) );
  NOR2X1 U58117 ( .A(n58499), .B(n43296), .Y(n54756) );
  NOR2X1 U58118 ( .A(n54757), .B(n54756), .Y(n54758) );
  NAND2X1 U58119 ( .A(n54759), .B(n54758), .Y(u_csr_N3672) );
  NAND2X1 U58120 ( .A(n43298), .B(n54763), .Y(n54761) );
  NAND2X1 U58121 ( .A(n43301), .B(n54762), .Y(n54760) );
  NAND2X1 U58122 ( .A(n54761), .B(n54760), .Y(net2288) );
  NOR2X1 U58123 ( .A(n2133), .B(n43306), .Y(n54766) );
  NAND2X1 U58124 ( .A(n43307), .B(n54762), .Y(n54765) );
  NAND2X1 U58125 ( .A(n43311), .B(n54763), .Y(n54764) );
  NAND2X1 U58126 ( .A(n54765), .B(n54764), .Y(n54773) );
  NOR2X1 U58127 ( .A(n54766), .B(n54773), .Y(n54768) );
  OR2X1 U58128 ( .A(n1765), .B(n42847), .Y(n54767) );
  NAND2X1 U58129 ( .A(n54768), .B(n54767), .Y(mem_i_pc_o[7]) );
  NOR2X1 U58130 ( .A(n43317), .B(n54775), .Y(net2387) );
  NOR2X1 U58131 ( .A(n43328), .B(n54772), .Y(n54774) );
  NOR2X1 U58132 ( .A(n54774), .B(n54773), .Y(n54779) );
  NOR2X1 U58133 ( .A(n2134), .B(n43320), .Y(n54777) );
  NOR2X1 U58134 ( .A(n43323), .B(n54775), .Y(n54776) );
  NOR2X1 U58135 ( .A(n54777), .B(n54776), .Y(n54778) );
  NAND2X1 U58136 ( .A(n54779), .B(n54778), .Y(u_decode_N297) );
  NAND2X1 U58137 ( .A(n43237), .B(n43853), .Y(n54789) );
  NOR2X1 U58138 ( .A(n29701), .B(n37342), .Y(n54787) );
  NAND2X1 U58139 ( .A(n29690), .B(n54897), .Y(n54785) );
  XNOR2X1 U58140 ( .A(n37898), .B(n54782), .Y(n54783) );
  NAND2X1 U58141 ( .A(n54903), .B(n54783), .Y(n54784) );
  NAND2X1 U58142 ( .A(n54785), .B(n54784), .Y(n54786) );
  OR2X1 U58143 ( .A(n54787), .B(n54786), .Y(n54883) );
  NAND2X1 U58144 ( .A(n43246), .B(n54883), .Y(n54788) );
  NAND2X1 U58145 ( .A(n54789), .B(n54788), .Y(n54794) );
  XNOR2X1 U58146 ( .A(opcode_pc_w[9]), .B(n42567), .Y(n54889) );
  INVX1 U58147 ( .A(n54889), .Y(n54801) );
  NAND2X1 U58148 ( .A(n54801), .B(n43240), .Y(n54792) );
  NAND2X1 U58149 ( .A(n44281), .B(n43856), .Y(n54804) );
  NAND2X1 U58150 ( .A(n27477), .B(n54804), .Y(n54790) );
  NAND2X1 U58151 ( .A(u_csr_csr_mepc_q[9]), .B(n54790), .Y(n54791) );
  NAND2X1 U58152 ( .A(n54792), .B(n54791), .Y(n54793) );
  NOR2X1 U58153 ( .A(n54794), .B(n54793), .Y(n54800) );
  NOR2X1 U58154 ( .A(n42953), .B(n37768), .Y(n54798) );
  NAND2X1 U58155 ( .A(n43244), .B(opcode_pc_w[9]), .Y(n54796) );
  NAND2X1 U58156 ( .A(n43286), .B(n54882), .Y(n54795) );
  NAND2X1 U58157 ( .A(n54796), .B(n54795), .Y(n54797) );
  NOR2X1 U58158 ( .A(n54798), .B(n54797), .Y(n54799) );
  NAND2X1 U58159 ( .A(n54800), .B(n54799), .Y(u_csr_csr_mepc_r[9]) );
  NAND2X1 U58160 ( .A(n43254), .B(n43853), .Y(n54803) );
  NAND2X1 U58161 ( .A(n54801), .B(n43250), .Y(n54802) );
  NAND2X1 U58162 ( .A(n54803), .B(n54802), .Y(n54809) );
  NAND2X1 U58163 ( .A(n43289), .B(n54883), .Y(n54807) );
  NAND2X1 U58164 ( .A(n26373), .B(n54804), .Y(n54805) );
  NAND2X1 U58165 ( .A(u_csr_csr_sepc_q[9]), .B(n54805), .Y(n54806) );
  NAND2X1 U58166 ( .A(n54807), .B(n54806), .Y(n54808) );
  NOR2X1 U58167 ( .A(n54809), .B(n54808), .Y(n54815) );
  NOR2X1 U58168 ( .A(n42955), .B(n37768), .Y(n54813) );
  NAND2X1 U58169 ( .A(n43257), .B(opcode_pc_w[9]), .Y(n54811) );
  NAND2X1 U58170 ( .A(n43259), .B(n54882), .Y(n54810) );
  NAND2X1 U58171 ( .A(n54811), .B(n54810), .Y(n54812) );
  NOR2X1 U58172 ( .A(n54813), .B(n54812), .Y(n54814) );
  NAND2X1 U58173 ( .A(n54815), .B(n54814), .Y(u_csr_csr_sepc_r[9]) );
  AND2X1 U58174 ( .A(n28438), .B(n28436), .Y(n54819) );
  NOR2X1 U58175 ( .A(n58505), .B(n43293), .Y(n54817) );
  NOR2X1 U58176 ( .A(n58504), .B(n43296), .Y(n54816) );
  NOR2X1 U58177 ( .A(n54817), .B(n54816), .Y(n54818) );
  NAND2X1 U58178 ( .A(n54819), .B(n54818), .Y(u_csr_N3674) );
  NAND2X1 U58179 ( .A(n43298), .B(n54883), .Y(n54821) );
  NAND2X1 U58180 ( .A(n43301), .B(n54882), .Y(n54820) );
  NAND2X1 U58181 ( .A(n54821), .B(n54820), .Y(net2290) );
  NOR2X1 U58182 ( .A(n29722), .B(n43014), .Y(n54830) );
  NAND2X1 U58183 ( .A(n29712), .B(n54897), .Y(n54828) );
  XNOR2X1 U58184 ( .A(n54825), .B(n54824), .Y(n54826) );
  NAND2X1 U58185 ( .A(n54903), .B(n54826), .Y(n54827) );
  NAND2X1 U58186 ( .A(n54828), .B(n54827), .Y(n54829) );
  OR2X1 U58187 ( .A(n54830), .B(n54829), .Y(n54876) );
  NAND2X1 U58188 ( .A(n43246), .B(n54876), .Y(n54834) );
  INVX1 U58189 ( .A(n54831), .Y(n55208) );
  XNOR2X1 U58190 ( .A(opcode_pc_w[8]), .B(n54832), .Y(n56808) );
  INVX1 U58191 ( .A(n56808), .Y(n54851) );
  NAND2X1 U58192 ( .A(n55208), .B(n54851), .Y(n54833) );
  NAND2X1 U58193 ( .A(n54834), .B(n54833), .Y(n54841) );
  NAND2X1 U58194 ( .A(n44281), .B(n44040), .Y(n58272) );
  NAND2X1 U58195 ( .A(n27477), .B(n58272), .Y(n54835) );
  NAND2X1 U58196 ( .A(u_csr_csr_mepc_q[8]), .B(n54835), .Y(n54839) );
  NOR2X1 U58197 ( .A(n42567), .B(n55039), .Y(n54837) );
  NAND2X1 U58198 ( .A(n54836), .B(n58441), .Y(n54855) );
  NAND2X1 U58199 ( .A(n54837), .B(n54855), .Y(n54838) );
  NAND2X1 U58200 ( .A(n54839), .B(n54838), .Y(n54840) );
  NOR2X1 U58201 ( .A(n54841), .B(n54840), .Y(n54849) );
  NAND2X1 U58202 ( .A(n2138), .B(n55540), .Y(n54843) );
  NAND2X1 U58203 ( .A(n43244), .B(opcode_pc_w[8]), .Y(n54842) );
  NAND2X1 U58204 ( .A(n54843), .B(n54842), .Y(n54847) );
  NAND2X1 U58205 ( .A(n43286), .B(n54875), .Y(n54845) );
  NAND2X1 U58206 ( .A(n43237), .B(n44038), .Y(n54844) );
  NAND2X1 U58207 ( .A(n54845), .B(n54844), .Y(n54846) );
  NOR2X1 U58208 ( .A(n54847), .B(n54846), .Y(n54848) );
  NAND2X1 U58209 ( .A(n54849), .B(n54848), .Y(u_csr_csr_mepc_r[8]) );
  NAND2X1 U58210 ( .A(n43289), .B(n54876), .Y(n54853) );
  INVX1 U58211 ( .A(n54850), .Y(n55228) );
  NAND2X1 U58212 ( .A(n55228), .B(n54851), .Y(n54852) );
  NAND2X1 U58213 ( .A(n54853), .B(n54852), .Y(n54860) );
  NAND2X1 U58214 ( .A(n26373), .B(n58272), .Y(n54854) );
  NAND2X1 U58215 ( .A(u_csr_csr_sepc_q[8]), .B(n54854), .Y(n54858) );
  NOR2X1 U58216 ( .A(n42567), .B(n55058), .Y(n54856) );
  NAND2X1 U58217 ( .A(n54856), .B(n54855), .Y(n54857) );
  NAND2X1 U58218 ( .A(n54858), .B(n54857), .Y(n54859) );
  NOR2X1 U58219 ( .A(n54860), .B(n54859), .Y(n54868) );
  NAND2X1 U58220 ( .A(n2138), .B(n58279), .Y(n54862) );
  NAND2X1 U58221 ( .A(n43257), .B(opcode_pc_w[8]), .Y(n54861) );
  NAND2X1 U58222 ( .A(n54862), .B(n54861), .Y(n54866) );
  NAND2X1 U58223 ( .A(n43259), .B(n54875), .Y(n54864) );
  NAND2X1 U58224 ( .A(n43254), .B(n44038), .Y(n54863) );
  NAND2X1 U58225 ( .A(n54864), .B(n54863), .Y(n54865) );
  NOR2X1 U58226 ( .A(n54866), .B(n54865), .Y(n54867) );
  NAND2X1 U58227 ( .A(n54868), .B(n54867), .Y(u_csr_csr_sepc_r[8]) );
  AND2X1 U58228 ( .A(n28446), .B(n28444), .Y(n54872) );
  NOR2X1 U58229 ( .A(n58503), .B(n43293), .Y(n54870) );
  NOR2X1 U58230 ( .A(n58502), .B(n43296), .Y(n54869) );
  NOR2X1 U58231 ( .A(n54870), .B(n54869), .Y(n54871) );
  NAND2X1 U58232 ( .A(n54872), .B(n54871), .Y(u_csr_N3673) );
  NAND2X1 U58233 ( .A(n43298), .B(n54876), .Y(n54874) );
  NAND2X1 U58234 ( .A(n43301), .B(n54875), .Y(n54873) );
  NAND2X1 U58235 ( .A(n54874), .B(n54873), .Y(net2289) );
  NOR2X1 U58236 ( .A(n2136), .B(n43306), .Y(n54879) );
  NAND2X1 U58237 ( .A(n43307), .B(n54875), .Y(n54878) );
  NAND2X1 U58238 ( .A(n43313), .B(n54876), .Y(n54877) );
  NAND2X1 U58239 ( .A(n54878), .B(n54877), .Y(n56809) );
  NOR2X1 U58240 ( .A(n54879), .B(n56809), .Y(n54881) );
  OR2X1 U58241 ( .A(n1766), .B(n42846), .Y(n54880) );
  NAND2X1 U58242 ( .A(n54881), .B(n54880), .Y(mem_i_pc_o[8]) );
  NOR2X1 U58243 ( .A(n2139), .B(n43306), .Y(n54886) );
  NAND2X1 U58244 ( .A(n43307), .B(n54882), .Y(n54885) );
  NAND2X1 U58245 ( .A(n43311), .B(n54883), .Y(n54884) );
  NAND2X1 U58246 ( .A(n54885), .B(n54884), .Y(n54890) );
  NOR2X1 U58247 ( .A(n54886), .B(n54890), .Y(n54888) );
  OR2X1 U58248 ( .A(n1767), .B(n42846), .Y(n54887) );
  NAND2X1 U58249 ( .A(n54888), .B(n54887), .Y(mem_i_pc_o[9]) );
  INVX1 U58250 ( .A(mem_i_pc_o[9]), .Y(n54958) );
  NAND2X1 U58251 ( .A(n42416), .B(mem_i_pc_o[8]), .Y(n55023) );
  NOR2X1 U58252 ( .A(n43317), .B(n54892), .Y(net2389) );
  NOR2X1 U58253 ( .A(n43328), .B(n54889), .Y(n54891) );
  NOR2X1 U58254 ( .A(n54891), .B(n54890), .Y(n54896) );
  NOR2X1 U58255 ( .A(n2140), .B(n43320), .Y(n54894) );
  NOR2X1 U58256 ( .A(n43323), .B(n54892), .Y(n54893) );
  NOR2X1 U58257 ( .A(n54894), .B(n54893), .Y(n54895) );
  NAND2X1 U58258 ( .A(n54896), .B(n54895), .Y(u_decode_N299) );
  NOR2X1 U58259 ( .A(n29939), .B(n37342), .Y(n54907) );
  NAND2X1 U58260 ( .A(n29929), .B(n54897), .Y(n54905) );
  XNOR2X1 U58261 ( .A(n54901), .B(n54900), .Y(n54902) );
  NAND2X1 U58262 ( .A(n54903), .B(n54902), .Y(n54904) );
  NAND2X1 U58263 ( .A(n54905), .B(n54904), .Y(n54906) );
  OR2X1 U58264 ( .A(n54907), .B(n54906), .Y(n54952) );
  NAND2X1 U58265 ( .A(n43246), .B(n54952), .Y(n54910) );
  XNOR2X1 U58266 ( .A(opcode_pc_w[10]), .B(n54908), .Y(n54960) );
  INVX1 U58267 ( .A(n54960), .Y(n54926) );
  NAND2X1 U58268 ( .A(n54926), .B(n55208), .Y(n54909) );
  NAND2X1 U58269 ( .A(n54910), .B(n54909), .Y(n54917) );
  NAND2X1 U58270 ( .A(n44281), .B(n43866), .Y(n54929) );
  NAND2X1 U58271 ( .A(n27477), .B(n54929), .Y(n54911) );
  NAND2X1 U58272 ( .A(u_csr_csr_mepc_q[10]), .B(n54911), .Y(n54915) );
  NOR2X1 U58273 ( .A(n42568), .B(n55039), .Y(n54913) );
  NAND2X1 U58274 ( .A(n54912), .B(n58280), .Y(n54931) );
  NAND2X1 U58275 ( .A(n54913), .B(n54931), .Y(n54914) );
  NAND2X1 U58276 ( .A(n54915), .B(n54914), .Y(n54916) );
  NOR2X1 U58277 ( .A(n54917), .B(n54916), .Y(n54925) );
  NAND2X1 U58278 ( .A(n2144), .B(n55540), .Y(n54919) );
  NAND2X1 U58279 ( .A(n43244), .B(opcode_pc_w[10]), .Y(n54918) );
  NAND2X1 U58280 ( .A(n54919), .B(n54918), .Y(n54923) );
  NAND2X1 U58281 ( .A(n43286), .B(n54951), .Y(n54921) );
  NAND2X1 U58282 ( .A(n43237), .B(n43862), .Y(n54920) );
  NAND2X1 U58283 ( .A(n54921), .B(n54920), .Y(n54922) );
  NOR2X1 U58284 ( .A(n54923), .B(n54922), .Y(n54924) );
  NAND2X1 U58285 ( .A(n54925), .B(n54924), .Y(u_csr_csr_mepc_r[10]) );
  NAND2X1 U58286 ( .A(n43289), .B(n54952), .Y(n54928) );
  NAND2X1 U58287 ( .A(n54926), .B(n55228), .Y(n54927) );
  NAND2X1 U58288 ( .A(n54928), .B(n54927), .Y(n54936) );
  NAND2X1 U58289 ( .A(n26373), .B(n54929), .Y(n54930) );
  NAND2X1 U58290 ( .A(u_csr_csr_sepc_q[10]), .B(n54930), .Y(n54934) );
  NOR2X1 U58291 ( .A(n42568), .B(n55058), .Y(n54932) );
  NAND2X1 U58292 ( .A(n54932), .B(n54931), .Y(n54933) );
  NAND2X1 U58293 ( .A(n54934), .B(n54933), .Y(n54935) );
  NOR2X1 U58294 ( .A(n54936), .B(n54935), .Y(n54944) );
  NAND2X1 U58295 ( .A(n2144), .B(n58279), .Y(n54938) );
  NAND2X1 U58296 ( .A(n43257), .B(opcode_pc_w[10]), .Y(n54937) );
  NAND2X1 U58297 ( .A(n54938), .B(n54937), .Y(n54942) );
  NAND2X1 U58298 ( .A(n43259), .B(n54951), .Y(n54940) );
  NAND2X1 U58299 ( .A(n43254), .B(n43862), .Y(n54939) );
  NAND2X1 U58300 ( .A(n54940), .B(n54939), .Y(n54941) );
  NOR2X1 U58301 ( .A(n54942), .B(n54941), .Y(n54943) );
  NAND2X1 U58302 ( .A(n54944), .B(n54943), .Y(u_csr_csr_sepc_r[10]) );
  AND2X1 U58303 ( .A(n28430), .B(n28428), .Y(n54948) );
  NOR2X1 U58304 ( .A(n58464), .B(n43293), .Y(n54946) );
  NOR2X1 U58305 ( .A(n58463), .B(n43296), .Y(n54945) );
  NOR2X1 U58306 ( .A(n54946), .B(n54945), .Y(n54947) );
  NAND2X1 U58307 ( .A(n54948), .B(n54947), .Y(u_csr_N3675) );
  NAND2X1 U58308 ( .A(n43298), .B(n54952), .Y(n54950) );
  NAND2X1 U58309 ( .A(n43301), .B(n54951), .Y(n54949) );
  NAND2X1 U58310 ( .A(n54950), .B(n54949), .Y(net2291) );
  NOR2X1 U58311 ( .A(n2142), .B(n43305), .Y(n54955) );
  NAND2X1 U58312 ( .A(n43307), .B(n54951), .Y(n54954) );
  NAND2X1 U58313 ( .A(n43313), .B(n54952), .Y(n54953) );
  NAND2X1 U58314 ( .A(n54954), .B(n54953), .Y(n54961) );
  NOR2X1 U58315 ( .A(n54955), .B(n54961), .Y(n54957) );
  OR2X1 U58316 ( .A(n1768), .B(n42846), .Y(n54956) );
  NAND2X1 U58317 ( .A(n54957), .B(n54956), .Y(mem_i_pc_o[10]) );
  INVX1 U58318 ( .A(mem_i_pc_o[10]), .Y(n55024) );
  NOR2X1 U58319 ( .A(n54958), .B(n55023), .Y(n54959) );
  XNOR2X1 U58320 ( .A(n55024), .B(n54959), .Y(u_fetch_N59) );
  NOR2X1 U58321 ( .A(n43317), .B(n54963), .Y(net2390) );
  NOR2X1 U58322 ( .A(n43327), .B(n54960), .Y(n54962) );
  NOR2X1 U58323 ( .A(n54962), .B(n54961), .Y(n54967) );
  NOR2X1 U58324 ( .A(n2143), .B(n43320), .Y(n54965) );
  NOR2X1 U58325 ( .A(n43323), .B(n54963), .Y(n54964) );
  NOR2X1 U58326 ( .A(n54965), .B(n54964), .Y(n54966) );
  NAND2X1 U58327 ( .A(n54967), .B(n54966), .Y(u_decode_N300) );
  NAND2X1 U58328 ( .A(n43237), .B(n43965), .Y(n54984) );
  NOR2X1 U58329 ( .A(n54969), .B(n42872), .Y(n54975) );
  NOR2X1 U58330 ( .A(n54973), .B(n42930), .Y(n54974) );
  NOR2X1 U58331 ( .A(n54975), .B(n54974), .Y(n54982) );
  INVX1 U58332 ( .A(n54976), .Y(n54978) );
  XNOR2X1 U58333 ( .A(n39115), .B(opcode_pc_w[11]), .Y(n54977) );
  XOR2X1 U58334 ( .A(n54978), .B(n54977), .Y(n54980) );
  NAND2X1 U58335 ( .A(n54980), .B(n54979), .Y(n54981) );
  NAND2X1 U58336 ( .A(n54982), .B(n54981), .Y(n55017) );
  NAND2X1 U58337 ( .A(n43246), .B(n55017), .Y(n54983) );
  NAND2X1 U58338 ( .A(n54984), .B(n54983), .Y(n54989) );
  XNOR2X1 U58339 ( .A(opcode_pc_w[11]), .B(n42568), .Y(n55025) );
  INVX1 U58340 ( .A(n55025), .Y(n54996) );
  NAND2X1 U58341 ( .A(n54996), .B(n43240), .Y(n54987) );
  NAND2X1 U58342 ( .A(n44281), .B(n43967), .Y(n58257) );
  NAND2X1 U58343 ( .A(n27477), .B(n58257), .Y(n54985) );
  NAND2X1 U58344 ( .A(u_csr_csr_mepc_q[11]), .B(n54985), .Y(n54986) );
  NAND2X1 U58345 ( .A(n54987), .B(n54986), .Y(n54988) );
  NOR2X1 U58346 ( .A(n54989), .B(n54988), .Y(n54995) );
  NOR2X1 U58347 ( .A(n42953), .B(n37769), .Y(n54993) );
  NAND2X1 U58348 ( .A(n43244), .B(opcode_pc_w[11]), .Y(n54991) );
  NAND2X1 U58349 ( .A(n43286), .B(n55016), .Y(n54990) );
  NAND2X1 U58350 ( .A(n54991), .B(n54990), .Y(n54992) );
  NOR2X1 U58351 ( .A(n54993), .B(n54992), .Y(n54994) );
  NAND2X1 U58352 ( .A(n54995), .B(n54994), .Y(u_csr_csr_mepc_r[11]) );
  NAND2X1 U58353 ( .A(n54996), .B(n43250), .Y(n54998) );
  NAND2X1 U58354 ( .A(n43289), .B(n55017), .Y(n54997) );
  NAND2X1 U58355 ( .A(n54998), .B(n54997), .Y(n55003) );
  NAND2X1 U58356 ( .A(n43254), .B(n43965), .Y(n55001) );
  NAND2X1 U58357 ( .A(n26373), .B(n58257), .Y(n54999) );
  NAND2X1 U58358 ( .A(u_csr_csr_sepc_q[11]), .B(n54999), .Y(n55000) );
  NAND2X1 U58359 ( .A(n55001), .B(n55000), .Y(n55002) );
  NOR2X1 U58360 ( .A(n55003), .B(n55002), .Y(n55009) );
  NOR2X1 U58361 ( .A(n42957), .B(n37769), .Y(n55007) );
  NAND2X1 U58362 ( .A(n43257), .B(opcode_pc_w[11]), .Y(n55005) );
  NAND2X1 U58363 ( .A(n43259), .B(n55016), .Y(n55004) );
  NAND2X1 U58364 ( .A(n55005), .B(n55004), .Y(n55006) );
  NOR2X1 U58365 ( .A(n55007), .B(n55006), .Y(n55008) );
  NAND2X1 U58366 ( .A(n55009), .B(n55008), .Y(u_csr_csr_sepc_r[11]) );
  AND2X1 U58367 ( .A(n28422), .B(n28420), .Y(n55013) );
  NOR2X1 U58368 ( .A(n58466), .B(n43293), .Y(n55011) );
  NOR2X1 U58369 ( .A(n58465), .B(n43296), .Y(n55010) );
  NOR2X1 U58370 ( .A(n55011), .B(n55010), .Y(n55012) );
  NAND2X1 U58371 ( .A(n55013), .B(n55012), .Y(u_csr_N3676) );
  NAND2X1 U58372 ( .A(n43298), .B(n55017), .Y(n55015) );
  NAND2X1 U58373 ( .A(n43301), .B(n55016), .Y(n55014) );
  NAND2X1 U58374 ( .A(n55015), .B(n55014), .Y(net2292) );
  NOR2X1 U58375 ( .A(n1931), .B(n43306), .Y(n55020) );
  NAND2X1 U58376 ( .A(n43307), .B(n55016), .Y(n55019) );
  NAND2X1 U58377 ( .A(n43313), .B(n55017), .Y(n55018) );
  NAND2X1 U58378 ( .A(n55019), .B(n55018), .Y(n55026) );
  NOR2X1 U58379 ( .A(n55020), .B(n55026), .Y(n55022) );
  OR2X1 U58380 ( .A(n1769), .B(n42847), .Y(n55021) );
  NAND2X1 U58381 ( .A(n55022), .B(n55021), .Y(mem_i_pc_o[11]) );
  NOR2X1 U58382 ( .A(n43316), .B(n55028), .Y(net2391) );
  NOR2X1 U58383 ( .A(n43327), .B(n55025), .Y(n55027) );
  NOR2X1 U58384 ( .A(n55027), .B(n55026), .Y(n55032) );
  NOR2X1 U58385 ( .A(n1932), .B(n43320), .Y(n55030) );
  NOR2X1 U58386 ( .A(n43323), .B(n55028), .Y(n55029) );
  NOR2X1 U58387 ( .A(n55030), .B(n55029), .Y(n55031) );
  NAND2X1 U58388 ( .A(n55032), .B(n55031), .Y(u_decode_N301) );
  NOR2X1 U58389 ( .A(n57411), .B(n42933), .Y(u_decode_N334) );
  NAND2X1 U58390 ( .A(n29569), .B(n73576), .Y(n24877) );
  INVX1 U58391 ( .A(n24877), .Y(n73503) );
  NAND2X1 U58392 ( .A(n55034), .B(n55033), .Y(n29634) );
  NOR2X1 U58393 ( .A(n24422), .B(n55035), .Y(u_decode_N778) );
  NAND2X1 U58394 ( .A(n43286), .B(n55084), .Y(n55037) );
  NAND2X1 U58395 ( .A(n43237), .B(n43955), .Y(n55036) );
  NAND2X1 U58396 ( .A(n55037), .B(n55036), .Y(n55047) );
  INVX1 U58397 ( .A(n55039), .Y(n55203) );
  NAND2X1 U58398 ( .A(n55203), .B(n55059), .Y(n55040) );
  NOR2X1 U58399 ( .A(n42465), .B(n55040), .Y(n55042) );
  NAND2X1 U58400 ( .A(n43958), .B(n44082), .Y(n73267) );
  NAND2X1 U58401 ( .A(u_csr_csr_mepc_q[12]), .B(n42131), .Y(n58468) );
  NOR2X1 U58402 ( .A(n73267), .B(n58468), .Y(n55041) );
  NOR2X1 U58403 ( .A(n55042), .B(n55041), .Y(n55045) );
  XNOR2X1 U58404 ( .A(opcode_pc_w[12]), .B(n55043), .Y(n55087) );
  INVX1 U58405 ( .A(n55087), .Y(n55064) );
  NAND2X1 U58406 ( .A(n55064), .B(n55208), .Y(n55044) );
  NAND2X1 U58407 ( .A(n55045), .B(n55044), .Y(n55046) );
  NOR2X1 U58408 ( .A(n55047), .B(n55046), .Y(n55055) );
  NAND2X1 U58409 ( .A(u_csr_csr_mepc_q[12]), .B(n42443), .Y(n55049) );
  NAND2X1 U58410 ( .A(n2147), .B(n55540), .Y(n55048) );
  NAND2X1 U58411 ( .A(n55049), .B(n55048), .Y(n55053) );
  NAND2X1 U58412 ( .A(n43244), .B(opcode_pc_w[12]), .Y(n55051) );
  NAND2X1 U58413 ( .A(n43246), .B(n55083), .Y(n55050) );
  NAND2X1 U58414 ( .A(n55051), .B(n55050), .Y(n55052) );
  NOR2X1 U58415 ( .A(n55053), .B(n55052), .Y(n55054) );
  NAND2X1 U58416 ( .A(n55055), .B(n55054), .Y(u_csr_csr_mepc_r[12]) );
  NAND2X1 U58417 ( .A(n43289), .B(n55083), .Y(n55057) );
  NAND2X1 U58418 ( .A(n43254), .B(n43955), .Y(n55056) );
  NAND2X1 U58419 ( .A(n55057), .B(n55056), .Y(n55068) );
  INVX1 U58420 ( .A(n55058), .Y(n55223) );
  NAND2X1 U58421 ( .A(n55223), .B(n55059), .Y(n55060) );
  NOR2X1 U58422 ( .A(n42465), .B(n55060), .Y(n55063) );
  INVX1 U58423 ( .A(n42965), .Y(n73501) );
  NAND2X1 U58424 ( .A(u_csr_csr_sepc_q[12]), .B(n73501), .Y(n58467) );
  NOR2X1 U58425 ( .A(n58467), .B(n73267), .Y(n55062) );
  NOR2X1 U58426 ( .A(n55063), .B(n55062), .Y(n55066) );
  NAND2X1 U58427 ( .A(n55064), .B(n55228), .Y(n55065) );
  NAND2X1 U58428 ( .A(n55066), .B(n55065), .Y(n55067) );
  NOR2X1 U58429 ( .A(n55068), .B(n55067), .Y(n55076) );
  NAND2X1 U58430 ( .A(u_csr_csr_sepc_q[12]), .B(n42134), .Y(n55070) );
  NAND2X1 U58431 ( .A(n2147), .B(n58279), .Y(n55069) );
  NAND2X1 U58432 ( .A(n55070), .B(n55069), .Y(n55074) );
  NAND2X1 U58433 ( .A(n43257), .B(opcode_pc_w[12]), .Y(n55072) );
  NAND2X1 U58434 ( .A(n43259), .B(n55084), .Y(n55071) );
  NAND2X1 U58435 ( .A(n55072), .B(n55071), .Y(n55073) );
  NOR2X1 U58436 ( .A(n55074), .B(n55073), .Y(n55075) );
  NAND2X1 U58437 ( .A(n55076), .B(n55075), .Y(u_csr_csr_sepc_r[12]) );
  AND2X1 U58438 ( .A(n28414), .B(n28412), .Y(n55082) );
  NOR2X1 U58439 ( .A(n55077), .B(n43293), .Y(n55080) );
  NOR2X1 U58440 ( .A(n55078), .B(n43296), .Y(n55079) );
  NOR2X1 U58441 ( .A(n55080), .B(n55079), .Y(n55081) );
  NAND2X1 U58442 ( .A(n55082), .B(n55081), .Y(u_csr_N3677) );
  NAND2X1 U58443 ( .A(n43298), .B(n55083), .Y(n55086) );
  NAND2X1 U58444 ( .A(n43301), .B(n55084), .Y(n55085) );
  NAND2X1 U58445 ( .A(n55086), .B(n55085), .Y(net2293) );
  NOR2X1 U58446 ( .A(n43316), .B(n55090), .Y(net2392) );
  NOR2X1 U58447 ( .A(n43327), .B(n55087), .Y(n55089) );
  NOR2X1 U58448 ( .A(n55089), .B(n55088), .Y(n55094) );
  NOR2X1 U58449 ( .A(n2146), .B(n43320), .Y(n55092) );
  NOR2X1 U58450 ( .A(n43323), .B(n55090), .Y(n55091) );
  NOR2X1 U58451 ( .A(n55092), .B(n55091), .Y(n55093) );
  NAND2X1 U58452 ( .A(n55094), .B(n55093), .Y(u_decode_N302) );
  NAND2X1 U58453 ( .A(n43287), .B(n55133), .Y(n55096) );
  NAND2X1 U58454 ( .A(n43237), .B(n43872), .Y(n55095) );
  NAND2X1 U58455 ( .A(n55096), .B(n55095), .Y(n55101) );
  NAND2X1 U58456 ( .A(n43875), .B(n44084), .Y(n73193) );
  INVX1 U58457 ( .A(n73193), .Y(n55113) );
  NAND2X1 U58458 ( .A(n42564), .B(n55113), .Y(n55099) );
  XNOR2X1 U58459 ( .A(opcode_pc_w[13]), .B(n55097), .Y(n55136) );
  INVX1 U58460 ( .A(n55136), .Y(n55112) );
  NAND2X1 U58461 ( .A(n55112), .B(n43240), .Y(n55098) );
  NAND2X1 U58462 ( .A(n55099), .B(n55098), .Y(n55100) );
  NOR2X1 U58463 ( .A(n55101), .B(n55100), .Y(n55109) );
  NAND2X1 U58464 ( .A(u_csr_csr_mepc_q[13]), .B(n42443), .Y(n55103) );
  NAND2X1 U58465 ( .A(n2150), .B(n55540), .Y(n55102) );
  NAND2X1 U58466 ( .A(n55103), .B(n55102), .Y(n55107) );
  NAND2X1 U58467 ( .A(n43244), .B(opcode_pc_w[13]), .Y(n55105) );
  NAND2X1 U58468 ( .A(n43246), .B(n55132), .Y(n55104) );
  NAND2X1 U58469 ( .A(n55105), .B(n55104), .Y(n55106) );
  NOR2X1 U58470 ( .A(n55107), .B(n55106), .Y(n55108) );
  NAND2X1 U58471 ( .A(n55109), .B(n55108), .Y(u_csr_csr_mepc_r[13]) );
  NAND2X1 U58472 ( .A(n43290), .B(n55132), .Y(n55111) );
  NAND2X1 U58473 ( .A(n43254), .B(n43872), .Y(n55110) );
  NAND2X1 U58474 ( .A(n55111), .B(n55110), .Y(n55117) );
  NAND2X1 U58475 ( .A(n55112), .B(n43250), .Y(n55115) );
  NAND2X1 U58476 ( .A(n55113), .B(n42569), .Y(n55114) );
  NAND2X1 U58477 ( .A(n55115), .B(n55114), .Y(n55116) );
  NOR2X1 U58478 ( .A(n55117), .B(n55116), .Y(n55125) );
  NAND2X1 U58479 ( .A(u_csr_csr_sepc_q[13]), .B(n42134), .Y(n55119) );
  NAND2X1 U58480 ( .A(n2150), .B(n58279), .Y(n55118) );
  NAND2X1 U58481 ( .A(n55119), .B(n55118), .Y(n55123) );
  NAND2X1 U58482 ( .A(n43257), .B(opcode_pc_w[13]), .Y(n55121) );
  NAND2X1 U58483 ( .A(n43259), .B(n55133), .Y(n55120) );
  NAND2X1 U58484 ( .A(n55121), .B(n55120), .Y(n55122) );
  NOR2X1 U58485 ( .A(n55123), .B(n55122), .Y(n55124) );
  NAND2X1 U58486 ( .A(n55125), .B(n55124), .Y(u_csr_csr_sepc_r[13]) );
  AND2X1 U58487 ( .A(n28406), .B(n28404), .Y(n55131) );
  NOR2X1 U58488 ( .A(n55126), .B(n43293), .Y(n55129) );
  NOR2X1 U58489 ( .A(n55127), .B(n43296), .Y(n55128) );
  NOR2X1 U58490 ( .A(n55129), .B(n55128), .Y(n55130) );
  NAND2X1 U58491 ( .A(n55131), .B(n55130), .Y(u_csr_N3678) );
  NAND2X1 U58492 ( .A(n43299), .B(n55132), .Y(n55135) );
  NAND2X1 U58493 ( .A(n43302), .B(n55133), .Y(n55134) );
  NAND2X1 U58494 ( .A(n55135), .B(n55134), .Y(net2294) );
  NAND2X1 U58495 ( .A(n42415), .B(n21), .Y(n55251) );
  NOR2X1 U58496 ( .A(n43316), .B(n55139), .Y(net2393) );
  NOR2X1 U58497 ( .A(n43327), .B(n55136), .Y(n55138) );
  NOR2X1 U58498 ( .A(n55138), .B(n55137), .Y(n55143) );
  NOR2X1 U58499 ( .A(n2149), .B(n43320), .Y(n55141) );
  NOR2X1 U58500 ( .A(n43323), .B(n55139), .Y(n55140) );
  NOR2X1 U58501 ( .A(n55141), .B(n55140), .Y(n55142) );
  NAND2X1 U58502 ( .A(n55143), .B(n55142), .Y(u_decode_N303) );
  NAND2X1 U58503 ( .A(n43287), .B(n55188), .Y(n55145) );
  NAND2X1 U58504 ( .A(n43237), .B(n43882), .Y(n55144) );
  NAND2X1 U58505 ( .A(n55145), .B(n55144), .Y(n55154) );
  NAND2X1 U58506 ( .A(n55203), .B(n55202), .Y(n55147) );
  NOR2X1 U58507 ( .A(n42463), .B(n55147), .Y(n55149) );
  NAND2X1 U58508 ( .A(n43884), .B(n44084), .Y(n73200) );
  NAND2X1 U58509 ( .A(u_csr_csr_mepc_q[14]), .B(n42131), .Y(n58472) );
  NOR2X1 U58510 ( .A(n73200), .B(n58472), .Y(n55148) );
  NOR2X1 U58511 ( .A(n55149), .B(n55148), .Y(n55152) );
  XNOR2X1 U58512 ( .A(opcode_pc_w[14]), .B(n55150), .Y(n55192) );
  INVX1 U58513 ( .A(n55192), .Y(n55168) );
  NAND2X1 U58514 ( .A(n55168), .B(n55208), .Y(n55151) );
  NAND2X1 U58515 ( .A(n55152), .B(n55151), .Y(n55153) );
  NOR2X1 U58516 ( .A(n55154), .B(n55153), .Y(n55162) );
  NAND2X1 U58517 ( .A(u_csr_csr_mepc_q[14]), .B(n42443), .Y(n55156) );
  NAND2X1 U58518 ( .A(n2153), .B(n55540), .Y(n55155) );
  NAND2X1 U58519 ( .A(n55156), .B(n55155), .Y(n55160) );
  NAND2X1 U58520 ( .A(n43244), .B(opcode_pc_w[14]), .Y(n55158) );
  NAND2X1 U58521 ( .A(n43246), .B(n55187), .Y(n55157) );
  NAND2X1 U58522 ( .A(n55158), .B(n55157), .Y(n55159) );
  NOR2X1 U58523 ( .A(n55160), .B(n55159), .Y(n55161) );
  NAND2X1 U58524 ( .A(n55162), .B(n55161), .Y(u_csr_csr_mepc_r[14]) );
  NAND2X1 U58525 ( .A(n43290), .B(n55187), .Y(n55164) );
  NAND2X1 U58526 ( .A(n43254), .B(n43882), .Y(n55163) );
  NAND2X1 U58527 ( .A(n55164), .B(n55163), .Y(n55172) );
  NAND2X1 U58528 ( .A(n55223), .B(n55202), .Y(n55165) );
  NOR2X1 U58529 ( .A(n42463), .B(n55165), .Y(n55167) );
  NAND2X1 U58530 ( .A(u_csr_csr_sepc_q[14]), .B(n73501), .Y(n58471) );
  NOR2X1 U58531 ( .A(n58471), .B(n73200), .Y(n55166) );
  NOR2X1 U58532 ( .A(n55167), .B(n55166), .Y(n55170) );
  NAND2X1 U58533 ( .A(n55168), .B(n55228), .Y(n55169) );
  NAND2X1 U58534 ( .A(n55170), .B(n55169), .Y(n55171) );
  NOR2X1 U58535 ( .A(n55172), .B(n55171), .Y(n55180) );
  NAND2X1 U58536 ( .A(u_csr_csr_sepc_q[14]), .B(n42134), .Y(n55174) );
  NAND2X1 U58537 ( .A(n2153), .B(n58279), .Y(n55173) );
  NAND2X1 U58538 ( .A(n55174), .B(n55173), .Y(n55178) );
  NAND2X1 U58539 ( .A(n43257), .B(opcode_pc_w[14]), .Y(n55176) );
  NAND2X1 U58540 ( .A(n43259), .B(n55188), .Y(n55175) );
  NAND2X1 U58541 ( .A(n55176), .B(n55175), .Y(n55177) );
  NOR2X1 U58542 ( .A(n55178), .B(n55177), .Y(n55179) );
  NAND2X1 U58543 ( .A(n55180), .B(n55179), .Y(u_csr_csr_sepc_r[14]) );
  AND2X1 U58544 ( .A(n28398), .B(n28396), .Y(n55186) );
  NOR2X1 U58545 ( .A(n55181), .B(n43293), .Y(n55184) );
  NOR2X1 U58546 ( .A(n55182), .B(n43296), .Y(n55183) );
  NOR2X1 U58547 ( .A(n55184), .B(n55183), .Y(n55185) );
  NAND2X1 U58548 ( .A(n55186), .B(n55185), .Y(u_csr_N3679) );
  NAND2X1 U58549 ( .A(n43299), .B(n55187), .Y(n55190) );
  NAND2X1 U58550 ( .A(n43302), .B(n55188), .Y(n55189) );
  NAND2X1 U58551 ( .A(n55190), .B(n55189), .Y(net2295) );
  INVX1 U58552 ( .A(n24), .Y(n55252) );
  NOR2X1 U58553 ( .A(n42406), .B(n55251), .Y(n55191) );
  XNOR2X1 U58554 ( .A(n55252), .B(n55191), .Y(u_fetch_N63) );
  NOR2X1 U58555 ( .A(n43316), .B(n55195), .Y(net2394) );
  NOR2X1 U58556 ( .A(n43327), .B(n55192), .Y(n55194) );
  NOR2X1 U58557 ( .A(n55194), .B(n55193), .Y(n55199) );
  NOR2X1 U58558 ( .A(n2152), .B(n43320), .Y(n55197) );
  NOR2X1 U58559 ( .A(n43323), .B(n55195), .Y(n55196) );
  NOR2X1 U58560 ( .A(n55197), .B(n55196), .Y(n55198) );
  NAND2X1 U58561 ( .A(n55199), .B(n55198), .Y(u_decode_N304) );
  NAND2X1 U58562 ( .A(n43287), .B(n55248), .Y(n55201) );
  NAND2X1 U58563 ( .A(n43237), .B(n43892), .Y(n55200) );
  NAND2X1 U58564 ( .A(n55201), .B(n55200), .Y(n55212) );
  NAND2X1 U58565 ( .A(n55203), .B(n55264), .Y(n55204) );
  NOR2X1 U58566 ( .A(n42462), .B(n55204), .Y(n55206) );
  NAND2X1 U58567 ( .A(n43894), .B(n44084), .Y(n73207) );
  NAND2X1 U58568 ( .A(u_csr_csr_mepc_q[15]), .B(n42131), .Y(n58474) );
  NOR2X1 U58569 ( .A(n73207), .B(n58474), .Y(n55205) );
  NOR2X1 U58570 ( .A(n55206), .B(n55205), .Y(n55210) );
  XNOR2X1 U58571 ( .A(opcode_pc_w[15]), .B(n55207), .Y(n55253) );
  INVX1 U58572 ( .A(n55253), .Y(n55227) );
  NAND2X1 U58573 ( .A(n55208), .B(n55227), .Y(n55209) );
  NAND2X1 U58574 ( .A(n55210), .B(n55209), .Y(n55211) );
  NOR2X1 U58575 ( .A(n55212), .B(n55211), .Y(n55220) );
  NAND2X1 U58576 ( .A(u_csr_csr_mepc_q[15]), .B(n42443), .Y(n55214) );
  NAND2X1 U58577 ( .A(n1896), .B(n55540), .Y(n55213) );
  NAND2X1 U58578 ( .A(n55214), .B(n55213), .Y(n55218) );
  NAND2X1 U58579 ( .A(n43244), .B(opcode_pc_w[15]), .Y(n55216) );
  NAND2X1 U58580 ( .A(n43247), .B(n55247), .Y(n55215) );
  NAND2X1 U58581 ( .A(n55216), .B(n55215), .Y(n55217) );
  NOR2X1 U58582 ( .A(n55218), .B(n55217), .Y(n55219) );
  NAND2X1 U58583 ( .A(n55220), .B(n55219), .Y(u_csr_csr_mepc_r[15]) );
  NAND2X1 U58584 ( .A(n43290), .B(n55247), .Y(n55222) );
  NAND2X1 U58585 ( .A(n43254), .B(n43892), .Y(n55221) );
  NAND2X1 U58586 ( .A(n55222), .B(n55221), .Y(n55232) );
  NAND2X1 U58587 ( .A(n55223), .B(n55264), .Y(n55224) );
  NOR2X1 U58588 ( .A(n42462), .B(n55224), .Y(n55226) );
  NAND2X1 U58589 ( .A(u_csr_csr_sepc_q[15]), .B(n73501), .Y(n58473) );
  NOR2X1 U58590 ( .A(n58473), .B(n73207), .Y(n55225) );
  NOR2X1 U58591 ( .A(n55226), .B(n55225), .Y(n55230) );
  NAND2X1 U58592 ( .A(n55228), .B(n55227), .Y(n55229) );
  NAND2X1 U58593 ( .A(n55230), .B(n55229), .Y(n55231) );
  NOR2X1 U58594 ( .A(n55232), .B(n55231), .Y(n55240) );
  NAND2X1 U58595 ( .A(u_csr_csr_sepc_q[15]), .B(n42134), .Y(n55234) );
  NAND2X1 U58596 ( .A(n1896), .B(n58279), .Y(n55233) );
  NAND2X1 U58597 ( .A(n55234), .B(n55233), .Y(n55238) );
  NAND2X1 U58598 ( .A(n43257), .B(opcode_pc_w[15]), .Y(n55236) );
  NAND2X1 U58599 ( .A(n43260), .B(n55248), .Y(n55235) );
  NAND2X1 U58600 ( .A(n55236), .B(n55235), .Y(n55237) );
  NOR2X1 U58601 ( .A(n55238), .B(n55237), .Y(n55239) );
  NAND2X1 U58602 ( .A(n55240), .B(n55239), .Y(u_csr_csr_sepc_r[15]) );
  AND2X1 U58603 ( .A(n28390), .B(n28388), .Y(n55246) );
  NOR2X1 U58604 ( .A(n55241), .B(n43293), .Y(n55244) );
  NOR2X1 U58605 ( .A(n55242), .B(n43296), .Y(n55243) );
  NOR2X1 U58606 ( .A(n55244), .B(n55243), .Y(n55245) );
  NAND2X1 U58607 ( .A(n55246), .B(n55245), .Y(u_csr_N3680) );
  NAND2X1 U58608 ( .A(n43299), .B(n55247), .Y(n55250) );
  NAND2X1 U58609 ( .A(n43302), .B(n55248), .Y(n55249) );
  NAND2X1 U58610 ( .A(n55250), .B(n55249), .Y(net2296) );
  NOR2X1 U58611 ( .A(n43316), .B(n55256), .Y(net2395) );
  NOR2X1 U58612 ( .A(n43327), .B(n55253), .Y(n55255) );
  NOR2X1 U58613 ( .A(n55255), .B(n55254), .Y(n55260) );
  NOR2X1 U58614 ( .A(n2156), .B(n43321), .Y(n55258) );
  NOR2X1 U58615 ( .A(n43324), .B(n55256), .Y(n55257) );
  NOR2X1 U58616 ( .A(n55258), .B(n55257), .Y(n55259) );
  NAND2X1 U58617 ( .A(n55260), .B(n55259), .Y(u_decode_N305) );
  NAND2X1 U58618 ( .A(u_csr_csr_mepc_q[16]), .B(n42131), .Y(n25458) );
  NAND2X1 U58619 ( .A(n43287), .B(n55301), .Y(n55262) );
  NAND2X1 U58620 ( .A(n43237), .B(n43899), .Y(n55261) );
  NAND2X1 U58621 ( .A(n55262), .B(n55261), .Y(n55269) );
  NAND2X1 U58622 ( .A(n43901), .B(n44084), .Y(n73214) );
  INVX1 U58623 ( .A(n73214), .Y(n55281) );
  INVX1 U58624 ( .A(n25458), .Y(n55263) );
  NAND2X1 U58625 ( .A(n55281), .B(n55263), .Y(n55267) );
  NAND2X1 U58626 ( .A(n55264), .B(n58319), .Y(n55265) );
  NAND2X1 U58627 ( .A(n55265), .B(n55324), .Y(n55313) );
  INVX1 U58628 ( .A(n55313), .Y(n55280) );
  NAND2X1 U58629 ( .A(n55280), .B(n43240), .Y(n55266) );
  NAND2X1 U58630 ( .A(n55267), .B(n55266), .Y(n55268) );
  NOR2X1 U58631 ( .A(n55269), .B(n55268), .Y(n55277) );
  NAND2X1 U58632 ( .A(u_csr_csr_mepc_q[16]), .B(n42443), .Y(n55271) );
  NAND2X1 U58633 ( .A(n2161), .B(n55540), .Y(n55270) );
  NAND2X1 U58634 ( .A(n55271), .B(n55270), .Y(n55275) );
  NAND2X1 U58635 ( .A(n43244), .B(opcode_pc_w[16]), .Y(n55273) );
  NAND2X1 U58636 ( .A(n43247), .B(n55300), .Y(n55272) );
  NAND2X1 U58637 ( .A(n55273), .B(n55272), .Y(n55274) );
  NOR2X1 U58638 ( .A(n55275), .B(n55274), .Y(n55276) );
  NAND2X1 U58639 ( .A(n55277), .B(n55276), .Y(u_csr_csr_mepc_r[16]) );
  NAND2X1 U58640 ( .A(n43290), .B(n55300), .Y(n55279) );
  NAND2X1 U58641 ( .A(n43254), .B(n43899), .Y(n55278) );
  NAND2X1 U58642 ( .A(n55279), .B(n55278), .Y(n55285) );
  NAND2X1 U58643 ( .A(n55280), .B(n43250), .Y(n55283) );
  NAND2X1 U58644 ( .A(n55281), .B(n42573), .Y(n55282) );
  NAND2X1 U58645 ( .A(n55283), .B(n55282), .Y(n55284) );
  NOR2X1 U58646 ( .A(n55285), .B(n55284), .Y(n55293) );
  NAND2X1 U58647 ( .A(u_csr_csr_sepc_q[16]), .B(n42134), .Y(n55287) );
  NAND2X1 U58648 ( .A(n2161), .B(n58279), .Y(n55286) );
  NAND2X1 U58649 ( .A(n55287), .B(n55286), .Y(n55291) );
  NAND2X1 U58650 ( .A(n43257), .B(opcode_pc_w[16]), .Y(n55289) );
  NAND2X1 U58651 ( .A(n43260), .B(n55301), .Y(n55288) );
  NAND2X1 U58652 ( .A(n55289), .B(n55288), .Y(n55290) );
  NOR2X1 U58653 ( .A(n55291), .B(n55290), .Y(n55292) );
  NAND2X1 U58654 ( .A(n55293), .B(n55292), .Y(u_csr_csr_sepc_r[16]) );
  AND2X1 U58655 ( .A(n28382), .B(n28380), .Y(n55299) );
  NOR2X1 U58656 ( .A(n43292), .B(n55294), .Y(n55297) );
  NOR2X1 U58657 ( .A(n55295), .B(n43296), .Y(n55296) );
  NOR2X1 U58658 ( .A(n55297), .B(n55296), .Y(n55298) );
  NAND2X1 U58659 ( .A(n55299), .B(n55298), .Y(u_csr_N3681) );
  NAND2X1 U58660 ( .A(n43299), .B(n55300), .Y(n55303) );
  NAND2X1 U58661 ( .A(n43302), .B(n55301), .Y(n55302) );
  NAND2X1 U58662 ( .A(n55303), .B(n55302), .Y(net2302) );
  NAND2X1 U58663 ( .A(challenge[101]), .B(n44854), .Y(n55304) );
  NAND2X1 U58664 ( .A(n42254), .B(n55304), .Y(n17309) );
  XNOR2X1 U58665 ( .A(n55305), .B(n42402), .Y(u_fetch_N65) );
  NOR2X1 U58666 ( .A(n44848), .B(n55306), .Y(n55311) );
  NOR2X1 U58667 ( .A(n55307), .B(n58179), .Y(n55309) );
  NOR2X1 U58668 ( .A(n55309), .B(n55308), .Y(n55310) );
  NAND2X1 U58669 ( .A(n55311), .B(n55310), .Y(n56771) );
  NAND2X1 U58670 ( .A(challenge[103]), .B(n44854), .Y(n55312) );
  NAND2X1 U58671 ( .A(n56771), .B(n55312), .Y(n17311) );
  NOR2X1 U58672 ( .A(n43316), .B(n55316), .Y(net2401) );
  NOR2X1 U58673 ( .A(n43327), .B(n55313), .Y(n55315) );
  NOR2X1 U58674 ( .A(n55315), .B(n55314), .Y(n55320) );
  NOR2X1 U58675 ( .A(n2160), .B(n43321), .Y(n55318) );
  NOR2X1 U58676 ( .A(n43324), .B(n55316), .Y(n55317) );
  NOR2X1 U58677 ( .A(n55318), .B(n55317), .Y(n55319) );
  NAND2X1 U58678 ( .A(n55320), .B(n55319), .Y(u_decode_N306) );
  NAND2X1 U58679 ( .A(u_csr_csr_mepc_q[17]), .B(n42131), .Y(n25438) );
  NAND2X1 U58680 ( .A(n43287), .B(n55361), .Y(n55322) );
  NAND2X1 U58681 ( .A(n43237), .B(n43906), .Y(n55321) );
  NAND2X1 U58682 ( .A(n55322), .B(n55321), .Y(n55329) );
  NAND2X1 U58683 ( .A(n43908), .B(n44084), .Y(n73222) );
  INVX1 U58684 ( .A(n73222), .Y(n55341) );
  INVX1 U58685 ( .A(n25438), .Y(n55323) );
  NAND2X1 U58686 ( .A(n55341), .B(n55323), .Y(n55327) );
  NAND2X1 U58687 ( .A(n55324), .B(n58324), .Y(n55325) );
  NAND2X1 U58688 ( .A(n55325), .B(n55374), .Y(n55364) );
  INVX1 U58689 ( .A(n55364), .Y(n55340) );
  NAND2X1 U58690 ( .A(n55340), .B(n43240), .Y(n55326) );
  NAND2X1 U58691 ( .A(n55327), .B(n55326), .Y(n55328) );
  NOR2X1 U58692 ( .A(n55329), .B(n55328), .Y(n55337) );
  NAND2X1 U58693 ( .A(u_csr_csr_mepc_q[17]), .B(n42443), .Y(n55331) );
  NAND2X1 U58694 ( .A(n2164), .B(n55540), .Y(n55330) );
  NAND2X1 U58695 ( .A(n55331), .B(n55330), .Y(n55335) );
  NAND2X1 U58696 ( .A(n43244), .B(opcode_pc_w[17]), .Y(n55333) );
  NAND2X1 U58697 ( .A(n43247), .B(n55360), .Y(n55332) );
  NAND2X1 U58698 ( .A(n55333), .B(n55332), .Y(n55334) );
  NOR2X1 U58699 ( .A(n55335), .B(n55334), .Y(n55336) );
  NAND2X1 U58700 ( .A(n55337), .B(n55336), .Y(u_csr_csr_mepc_r[17]) );
  NAND2X1 U58701 ( .A(n43290), .B(n55360), .Y(n55339) );
  NAND2X1 U58702 ( .A(n43254), .B(n43906), .Y(n55338) );
  NAND2X1 U58703 ( .A(n55339), .B(n55338), .Y(n55345) );
  NAND2X1 U58704 ( .A(n55340), .B(n43250), .Y(n55343) );
  NAND2X1 U58705 ( .A(n55341), .B(n42572), .Y(n55342) );
  NAND2X1 U58706 ( .A(n55343), .B(n55342), .Y(n55344) );
  NOR2X1 U58707 ( .A(n55345), .B(n55344), .Y(n55353) );
  NAND2X1 U58708 ( .A(u_csr_csr_sepc_q[17]), .B(n42134), .Y(n55347) );
  NAND2X1 U58709 ( .A(n2164), .B(n58279), .Y(n55346) );
  NAND2X1 U58710 ( .A(n55347), .B(n55346), .Y(n55351) );
  NAND2X1 U58711 ( .A(n43257), .B(opcode_pc_w[17]), .Y(n55349) );
  NAND2X1 U58712 ( .A(n43260), .B(n55361), .Y(n55348) );
  NAND2X1 U58713 ( .A(n55349), .B(n55348), .Y(n55350) );
  NOR2X1 U58714 ( .A(n55351), .B(n55350), .Y(n55352) );
  NAND2X1 U58715 ( .A(n55353), .B(n55352), .Y(u_csr_csr_sepc_r[17]) );
  AND2X1 U58716 ( .A(n28374), .B(n28372), .Y(n55359) );
  NOR2X1 U58717 ( .A(n43292), .B(n55354), .Y(n55357) );
  NOR2X1 U58718 ( .A(n55355), .B(n43296), .Y(n55356) );
  NOR2X1 U58719 ( .A(n55357), .B(n55356), .Y(n55358) );
  NAND2X1 U58720 ( .A(n55359), .B(n55358), .Y(u_csr_N3682) );
  NAND2X1 U58721 ( .A(n43299), .B(n55360), .Y(n55363) );
  NAND2X1 U58722 ( .A(n43302), .B(n55361), .Y(n55362) );
  NAND2X1 U58723 ( .A(n55363), .B(n55362), .Y(net2303) );
  NAND2X1 U58724 ( .A(n42402), .B(n8), .Y(n55467) );
  NOR2X1 U58725 ( .A(n43316), .B(n55367), .Y(net2402) );
  NOR2X1 U58726 ( .A(n43327), .B(n55364), .Y(n55366) );
  NOR2X1 U58727 ( .A(n55366), .B(n55365), .Y(n55371) );
  NOR2X1 U58728 ( .A(n2163), .B(n43321), .Y(n55369) );
  NOR2X1 U58729 ( .A(n43324), .B(n55367), .Y(n55368) );
  NOR2X1 U58730 ( .A(n55369), .B(n55368), .Y(n55370) );
  NAND2X1 U58731 ( .A(n55371), .B(n55370), .Y(u_decode_N307) );
  NAND2X1 U58732 ( .A(n43247), .B(n55412), .Y(n55373) );
  NAND2X1 U58733 ( .A(n43287), .B(n55413), .Y(n55372) );
  NAND2X1 U58734 ( .A(n55373), .B(n55372), .Y(n55380) );
  NAND2X1 U58735 ( .A(n43237), .B(n43912), .Y(n55378) );
  NAND2X1 U58736 ( .A(n55374), .B(n58331), .Y(n55376) );
  NAND2X1 U58737 ( .A(n55376), .B(n55375), .Y(n55418) );
  INVX1 U58738 ( .A(n55418), .Y(n55391) );
  NAND2X1 U58739 ( .A(n55391), .B(n43240), .Y(n55377) );
  NAND2X1 U58740 ( .A(n55378), .B(n55377), .Y(n55379) );
  NOR2X1 U58741 ( .A(n55380), .B(n55379), .Y(n55388) );
  NAND2X1 U58742 ( .A(u_csr_csr_mepc_q[18]), .B(n42443), .Y(n55382) );
  NAND2X1 U58743 ( .A(n43914), .B(n44084), .Y(n73230) );
  INVX1 U58744 ( .A(n73230), .Y(n55397) );
  NAND2X1 U58745 ( .A(n42566), .B(n55397), .Y(n55381) );
  NAND2X1 U58746 ( .A(n55382), .B(n55381), .Y(n55386) );
  NAND2X1 U58747 ( .A(n2167), .B(n55540), .Y(n55384) );
  NAND2X1 U58748 ( .A(n43244), .B(opcode_pc_w[18]), .Y(n55383) );
  NAND2X1 U58749 ( .A(n55384), .B(n55383), .Y(n55385) );
  NOR2X1 U58750 ( .A(n55386), .B(n55385), .Y(n55387) );
  NAND2X1 U58751 ( .A(n55388), .B(n55387), .Y(u_csr_csr_mepc_r[18]) );
  NAND2X1 U58752 ( .A(u_csr_csr_sepc_q[18]), .B(n73501), .Y(n25420) );
  NAND2X1 U58753 ( .A(n43260), .B(n55413), .Y(n55390) );
  NAND2X1 U58754 ( .A(n43290), .B(n55412), .Y(n55389) );
  NAND2X1 U58755 ( .A(n55390), .B(n55389), .Y(n55395) );
  NAND2X1 U58756 ( .A(n43254), .B(n43912), .Y(n55393) );
  NAND2X1 U58757 ( .A(n55391), .B(n43250), .Y(n55392) );
  NAND2X1 U58758 ( .A(n55393), .B(n55392), .Y(n55394) );
  NOR2X1 U58759 ( .A(n55395), .B(n55394), .Y(n55405) );
  NAND2X1 U58760 ( .A(u_csr_csr_sepc_q[18]), .B(n42134), .Y(n55399) );
  INVX1 U58761 ( .A(n25420), .Y(n55396) );
  NAND2X1 U58762 ( .A(n55397), .B(n55396), .Y(n55398) );
  NAND2X1 U58763 ( .A(n55399), .B(n55398), .Y(n55403) );
  NAND2X1 U58764 ( .A(n2167), .B(n58279), .Y(n55401) );
  NAND2X1 U58765 ( .A(n43257), .B(opcode_pc_w[18]), .Y(n55400) );
  NAND2X1 U58766 ( .A(n55401), .B(n55400), .Y(n55402) );
  NOR2X1 U58767 ( .A(n55403), .B(n55402), .Y(n55404) );
  NAND2X1 U58768 ( .A(n55405), .B(n55404), .Y(u_csr_csr_sepc_r[18]) );
  AND2X1 U58769 ( .A(n28366), .B(n28364), .Y(n55411) );
  NOR2X1 U58770 ( .A(n55406), .B(n43293), .Y(n55409) );
  NOR2X1 U58771 ( .A(n43295), .B(n55407), .Y(n55408) );
  NOR2X1 U58772 ( .A(n55409), .B(n55408), .Y(n55410) );
  NAND2X1 U58773 ( .A(n55411), .B(n55410), .Y(u_csr_N3683) );
  NAND2X1 U58774 ( .A(n43299), .B(n55412), .Y(n55415) );
  NAND2X1 U58775 ( .A(n43302), .B(n55413), .Y(n55414) );
  NAND2X1 U58776 ( .A(n55415), .B(n55414), .Y(net2304) );
  INVX1 U58777 ( .A(n10), .Y(n55468) );
  NOR2X1 U58778 ( .A(n55416), .B(n55467), .Y(n55417) );
  XNOR2X1 U58779 ( .A(n55468), .B(n55417), .Y(u_fetch_N67) );
  NOR2X1 U58780 ( .A(n43316), .B(n55421), .Y(net2403) );
  NOR2X1 U58781 ( .A(n43327), .B(n55418), .Y(n55420) );
  NOR2X1 U58782 ( .A(n55420), .B(n55419), .Y(n55425) );
  NOR2X1 U58783 ( .A(n2166), .B(n43321), .Y(n55423) );
  NOR2X1 U58784 ( .A(n43324), .B(n55421), .Y(n55422) );
  NOR2X1 U58785 ( .A(n55423), .B(n55422), .Y(n55424) );
  NAND2X1 U58786 ( .A(n55425), .B(n55424), .Y(u_decode_N308) );
  NAND2X1 U58787 ( .A(u_csr_csr_mepc_q[19]), .B(n42131), .Y(n25396) );
  NAND2X1 U58788 ( .A(n43287), .B(n55464), .Y(n55427) );
  NAND2X1 U58789 ( .A(n43237), .B(n43921), .Y(n55426) );
  NAND2X1 U58790 ( .A(n55427), .B(n55426), .Y(n55432) );
  NAND2X1 U58791 ( .A(n43922), .B(n44084), .Y(n73238) );
  INVX1 U58792 ( .A(n73238), .Y(n55444) );
  INVX1 U58793 ( .A(n25396), .Y(n55428) );
  NAND2X1 U58794 ( .A(n55444), .B(n55428), .Y(n55430) );
  XNOR2X1 U58795 ( .A(opcode_pc_w[19]), .B(n55480), .Y(n55470) );
  INVX1 U58796 ( .A(n55470), .Y(n55443) );
  NAND2X1 U58797 ( .A(n55443), .B(n43240), .Y(n55429) );
  NAND2X1 U58798 ( .A(n55430), .B(n55429), .Y(n55431) );
  NOR2X1 U58799 ( .A(n55432), .B(n55431), .Y(n55440) );
  NAND2X1 U58800 ( .A(u_csr_csr_mepc_q[19]), .B(n42443), .Y(n55434) );
  NAND2X1 U58801 ( .A(n2170), .B(n55540), .Y(n55433) );
  NAND2X1 U58802 ( .A(n55434), .B(n55433), .Y(n55438) );
  NAND2X1 U58803 ( .A(n43244), .B(opcode_pc_w[19]), .Y(n55436) );
  NAND2X1 U58804 ( .A(n43247), .B(n55463), .Y(n55435) );
  NAND2X1 U58805 ( .A(n55436), .B(n55435), .Y(n55437) );
  NOR2X1 U58806 ( .A(n55438), .B(n55437), .Y(n55439) );
  NAND2X1 U58807 ( .A(n55440), .B(n55439), .Y(u_csr_csr_mepc_r[19]) );
  NAND2X1 U58808 ( .A(n43290), .B(n55463), .Y(n55442) );
  NAND2X1 U58809 ( .A(n43254), .B(n43921), .Y(n55441) );
  NAND2X1 U58810 ( .A(n55442), .B(n55441), .Y(n55448) );
  NAND2X1 U58811 ( .A(n55443), .B(n43250), .Y(n55446) );
  NAND2X1 U58812 ( .A(n55444), .B(n42571), .Y(n55445) );
  NAND2X1 U58813 ( .A(n55446), .B(n55445), .Y(n55447) );
  NOR2X1 U58814 ( .A(n55448), .B(n55447), .Y(n55456) );
  NAND2X1 U58815 ( .A(u_csr_csr_sepc_q[19]), .B(n42134), .Y(n55450) );
  NAND2X1 U58816 ( .A(n2170), .B(n58279), .Y(n55449) );
  NAND2X1 U58817 ( .A(n55450), .B(n55449), .Y(n55454) );
  NAND2X1 U58818 ( .A(n43257), .B(opcode_pc_w[19]), .Y(n55452) );
  NAND2X1 U58819 ( .A(n43260), .B(n55464), .Y(n55451) );
  NAND2X1 U58820 ( .A(n55452), .B(n55451), .Y(n55453) );
  NOR2X1 U58821 ( .A(n55454), .B(n55453), .Y(n55455) );
  NAND2X1 U58822 ( .A(n55456), .B(n55455), .Y(u_csr_csr_sepc_r[19]) );
  AND2X1 U58823 ( .A(n28358), .B(n28356), .Y(n55462) );
  NOR2X1 U58824 ( .A(n43292), .B(n55457), .Y(n55460) );
  NOR2X1 U58825 ( .A(n55458), .B(n43296), .Y(n55459) );
  NOR2X1 U58826 ( .A(n55460), .B(n55459), .Y(n55461) );
  NAND2X1 U58827 ( .A(n55462), .B(n55461), .Y(u_csr_N3684) );
  NAND2X1 U58828 ( .A(n43299), .B(n55463), .Y(n55466) );
  NAND2X1 U58829 ( .A(n43302), .B(n55464), .Y(n55465) );
  NAND2X1 U58830 ( .A(n55466), .B(n55465), .Y(net2305) );
  XNOR2X1 U58831 ( .A(n55469), .B(n42397), .Y(u_fetch_N68) );
  NOR2X1 U58832 ( .A(n43316), .B(n55473), .Y(net2404) );
  NOR2X1 U58833 ( .A(n43327), .B(n55470), .Y(n55472) );
  NOR2X1 U58834 ( .A(n55472), .B(n55471), .Y(n55477) );
  NOR2X1 U58835 ( .A(n2169), .B(n43321), .Y(n55475) );
  NOR2X1 U58836 ( .A(n43324), .B(n55473), .Y(n55474) );
  NOR2X1 U58837 ( .A(n55475), .B(n55474), .Y(n55476) );
  NAND2X1 U58838 ( .A(n55477), .B(n55476), .Y(u_decode_N309) );
  NAND2X1 U58839 ( .A(n43287), .B(n55519), .Y(n55479) );
  NAND2X1 U58840 ( .A(n43236), .B(n43929), .Y(n55478) );
  NAND2X1 U58841 ( .A(n55479), .B(n55478), .Y(n55486) );
  NAND2X1 U58842 ( .A(n43931), .B(n44084), .Y(n73245) );
  INVX1 U58843 ( .A(n73245), .Y(n55499) );
  NAND2X1 U58844 ( .A(n42565), .B(n55499), .Y(n55484) );
  NAND2X1 U58845 ( .A(n55480), .B(opcode_pc_w[19]), .Y(n55481) );
  NAND2X1 U58846 ( .A(n55481), .B(n58344), .Y(n55482) );
  NAND2X1 U58847 ( .A(n55482), .B(n55534), .Y(n55523) );
  INVX1 U58848 ( .A(n55523), .Y(n55497) );
  NAND2X1 U58849 ( .A(n55497), .B(n43239), .Y(n55483) );
  NAND2X1 U58850 ( .A(n55484), .B(n55483), .Y(n55485) );
  NOR2X1 U58851 ( .A(n55486), .B(n55485), .Y(n55494) );
  NAND2X1 U58852 ( .A(u_csr_csr_mepc_q[20]), .B(n42443), .Y(n55488) );
  NAND2X1 U58853 ( .A(n2173), .B(n55540), .Y(n55487) );
  NAND2X1 U58854 ( .A(n55488), .B(n55487), .Y(n55492) );
  NAND2X1 U58855 ( .A(n43243), .B(opcode_pc_w[20]), .Y(n55490) );
  NAND2X1 U58856 ( .A(n43247), .B(n55518), .Y(n55489) );
  NAND2X1 U58857 ( .A(n55490), .B(n55489), .Y(n55491) );
  NOR2X1 U58858 ( .A(n55492), .B(n55491), .Y(n55493) );
  NAND2X1 U58859 ( .A(n55494), .B(n55493), .Y(u_csr_csr_mepc_r[20]) );
  NAND2X1 U58860 ( .A(u_csr_csr_sepc_q[20]), .B(n73501), .Y(n25343) );
  NAND2X1 U58861 ( .A(n43290), .B(n55518), .Y(n55496) );
  NAND2X1 U58862 ( .A(n43253), .B(n43929), .Y(n55495) );
  NAND2X1 U58863 ( .A(n55496), .B(n55495), .Y(n55503) );
  NAND2X1 U58864 ( .A(n55497), .B(n43249), .Y(n55501) );
  INVX1 U58865 ( .A(n25343), .Y(n55498) );
  NAND2X1 U58866 ( .A(n55499), .B(n55498), .Y(n55500) );
  NAND2X1 U58867 ( .A(n55501), .B(n55500), .Y(n55502) );
  NOR2X1 U58868 ( .A(n55503), .B(n55502), .Y(n55511) );
  NAND2X1 U58869 ( .A(u_csr_csr_sepc_q[20]), .B(n42134), .Y(n55505) );
  NAND2X1 U58870 ( .A(n2173), .B(n58279), .Y(n55504) );
  NAND2X1 U58871 ( .A(n55505), .B(n55504), .Y(n55509) );
  NAND2X1 U58872 ( .A(n43256), .B(opcode_pc_w[20]), .Y(n55507) );
  NAND2X1 U58873 ( .A(n43260), .B(n55519), .Y(n55506) );
  NAND2X1 U58874 ( .A(n55507), .B(n55506), .Y(n55508) );
  NOR2X1 U58875 ( .A(n55509), .B(n55508), .Y(n55510) );
  NAND2X1 U58876 ( .A(n55511), .B(n55510), .Y(u_csr_csr_sepc_r[20]) );
  AND2X1 U58877 ( .A(n28350), .B(n28348), .Y(n55517) );
  NOR2X1 U58878 ( .A(n55512), .B(n43292), .Y(n55515) );
  NOR2X1 U58879 ( .A(n43295), .B(n55513), .Y(n55514) );
  NOR2X1 U58880 ( .A(n55515), .B(n55514), .Y(n55516) );
  NAND2X1 U58881 ( .A(n55517), .B(n55516), .Y(u_csr_N3685) );
  NAND2X1 U58882 ( .A(n43299), .B(n55518), .Y(n55521) );
  NAND2X1 U58883 ( .A(n43302), .B(n55519), .Y(n55520) );
  NAND2X1 U58884 ( .A(n55521), .B(n55520), .Y(net2306) );
  XNOR2X1 U58885 ( .A(n55522), .B(n42412), .Y(u_fetch_N69) );
  NOR2X1 U58886 ( .A(n43316), .B(n55526), .Y(net2405) );
  NOR2X1 U58887 ( .A(n43327), .B(n55523), .Y(n55525) );
  NOR2X1 U58888 ( .A(n55525), .B(n55524), .Y(n55530) );
  NOR2X1 U58889 ( .A(n2172), .B(n43321), .Y(n55528) );
  NOR2X1 U58890 ( .A(n43324), .B(n55526), .Y(n55527) );
  NOR2X1 U58891 ( .A(n55528), .B(n55527), .Y(n55529) );
  NAND2X1 U58892 ( .A(n55530), .B(n55529), .Y(u_decode_N310) );
  NAND2X1 U58893 ( .A(u_csr_csr_mepc_q[21]), .B(n42131), .Y(n25320) );
  NAND2X1 U58894 ( .A(n43287), .B(n55572), .Y(n55532) );
  NAND2X1 U58895 ( .A(n43236), .B(n43936), .Y(n55531) );
  NAND2X1 U58896 ( .A(n55532), .B(n55531), .Y(n55539) );
  NAND2X1 U58897 ( .A(n43939), .B(n44084), .Y(n73252) );
  INVX1 U58898 ( .A(n73252), .Y(n55552) );
  INVX1 U58899 ( .A(n25320), .Y(n55533) );
  NAND2X1 U58900 ( .A(n55552), .B(n55533), .Y(n55537) );
  NAND2X1 U58901 ( .A(n55534), .B(n58349), .Y(n55535) );
  NAND2X1 U58902 ( .A(n55535), .B(n55585), .Y(n55575) );
  INVX1 U58903 ( .A(n55575), .Y(n55551) );
  NAND2X1 U58904 ( .A(n55551), .B(n43239), .Y(n55536) );
  NAND2X1 U58905 ( .A(n55537), .B(n55536), .Y(n55538) );
  NOR2X1 U58906 ( .A(n55539), .B(n55538), .Y(n55548) );
  NAND2X1 U58907 ( .A(u_csr_csr_mepc_q[21]), .B(n42443), .Y(n55542) );
  NAND2X1 U58908 ( .A(n2176), .B(n55540), .Y(n55541) );
  NAND2X1 U58909 ( .A(n55542), .B(n55541), .Y(n55546) );
  NAND2X1 U58910 ( .A(n43243), .B(opcode_pc_w[21]), .Y(n55544) );
  NAND2X1 U58911 ( .A(n43247), .B(n55571), .Y(n55543) );
  NAND2X1 U58912 ( .A(n55544), .B(n55543), .Y(n55545) );
  NOR2X1 U58913 ( .A(n55546), .B(n55545), .Y(n55547) );
  NAND2X1 U58914 ( .A(n55548), .B(n55547), .Y(u_csr_csr_mepc_r[21]) );
  NAND2X1 U58915 ( .A(n43290), .B(n55571), .Y(n55550) );
  NAND2X1 U58916 ( .A(n43253), .B(n43936), .Y(n55549) );
  NAND2X1 U58917 ( .A(n55550), .B(n55549), .Y(n55556) );
  NAND2X1 U58918 ( .A(n55551), .B(n43249), .Y(n55554) );
  NAND2X1 U58919 ( .A(n55552), .B(n42570), .Y(n55553) );
  NAND2X1 U58920 ( .A(n55554), .B(n55553), .Y(n55555) );
  NOR2X1 U58921 ( .A(n55556), .B(n55555), .Y(n55564) );
  NAND2X1 U58922 ( .A(u_csr_csr_sepc_q[21]), .B(n42134), .Y(n55558) );
  NAND2X1 U58923 ( .A(n2176), .B(n58279), .Y(n55557) );
  NAND2X1 U58924 ( .A(n55558), .B(n55557), .Y(n55562) );
  NAND2X1 U58925 ( .A(n43256), .B(opcode_pc_w[21]), .Y(n55560) );
  NAND2X1 U58926 ( .A(n43260), .B(n55572), .Y(n55559) );
  NAND2X1 U58927 ( .A(n55560), .B(n55559), .Y(n55561) );
  NOR2X1 U58928 ( .A(n55562), .B(n55561), .Y(n55563) );
  NAND2X1 U58929 ( .A(n55564), .B(n55563), .Y(u_csr_csr_sepc_r[21]) );
  AND2X1 U58930 ( .A(n28342), .B(n28340), .Y(n55570) );
  NOR2X1 U58931 ( .A(n43292), .B(n55565), .Y(n55568) );
  NOR2X1 U58932 ( .A(n55566), .B(n43295), .Y(n55567) );
  NOR2X1 U58933 ( .A(n55568), .B(n55567), .Y(n55569) );
  NAND2X1 U58934 ( .A(n55570), .B(n55569), .Y(u_csr_N3686) );
  NAND2X1 U58935 ( .A(n43299), .B(n55571), .Y(n55574) );
  NAND2X1 U58936 ( .A(n43302), .B(n55572), .Y(n55573) );
  NAND2X1 U58937 ( .A(n55574), .B(n55573), .Y(net2307) );
  INVX1 U58938 ( .A(n12), .Y(n55623) );
  NAND2X1 U58939 ( .A(n42412), .B(n7), .Y(n55670) );
  NOR2X1 U58940 ( .A(n43316), .B(n55578), .Y(net2406) );
  NOR2X1 U58941 ( .A(n43326), .B(n55575), .Y(n55577) );
  NOR2X1 U58942 ( .A(n55577), .B(n55576), .Y(n55582) );
  NOR2X1 U58943 ( .A(n2175), .B(n43321), .Y(n55580) );
  NOR2X1 U58944 ( .A(n43324), .B(n55578), .Y(n55579) );
  NOR2X1 U58945 ( .A(n55580), .B(n55579), .Y(n55581) );
  NAND2X1 U58946 ( .A(n55582), .B(n55581), .Y(u_decode_N311) );
  NAND2X1 U58947 ( .A(n43287), .B(n55620), .Y(n55584) );
  NAND2X1 U58948 ( .A(n43236), .B(n43945), .Y(n55583) );
  NAND2X1 U58949 ( .A(n55584), .B(n55583), .Y(n55592) );
  NAND2X1 U58950 ( .A(n55585), .B(n58356), .Y(n55587) );
  NAND2X1 U58951 ( .A(n55587), .B(n55586), .Y(n55625) );
  INVX1 U58952 ( .A(n55625), .Y(n55601) );
  NAND2X1 U58953 ( .A(n55601), .B(n43239), .Y(n55590) );
  NAND2X1 U58954 ( .A(n44282), .B(n43949), .Y(n55602) );
  NAND2X1 U58955 ( .A(n27477), .B(n55602), .Y(n55588) );
  NAND2X1 U58956 ( .A(u_csr_csr_mepc_q[22]), .B(n55588), .Y(n55589) );
  NAND2X1 U58957 ( .A(n55590), .B(n55589), .Y(n55591) );
  NOR2X1 U58958 ( .A(n55592), .B(n55591), .Y(n55598) );
  NOR2X1 U58959 ( .A(n42952), .B(n37770), .Y(n55596) );
  NAND2X1 U58960 ( .A(n43243), .B(opcode_pc_w[22]), .Y(n55594) );
  NAND2X1 U58961 ( .A(n43247), .B(n55619), .Y(n55593) );
  NAND2X1 U58962 ( .A(n55594), .B(n55593), .Y(n55595) );
  NOR2X1 U58963 ( .A(n55596), .B(n55595), .Y(n55597) );
  NAND2X1 U58964 ( .A(n55598), .B(n55597), .Y(u_csr_csr_mepc_r[22]) );
  NAND2X1 U58965 ( .A(n43290), .B(n55619), .Y(n55600) );
  NAND2X1 U58966 ( .A(n43253), .B(n43945), .Y(n55599) );
  NAND2X1 U58967 ( .A(n55600), .B(n55599), .Y(n55607) );
  NAND2X1 U58968 ( .A(n55601), .B(n43249), .Y(n55605) );
  NAND2X1 U58969 ( .A(n26373), .B(n55602), .Y(n55603) );
  NAND2X1 U58970 ( .A(u_csr_csr_sepc_q[22]), .B(n55603), .Y(n55604) );
  NAND2X1 U58971 ( .A(n55605), .B(n55604), .Y(n55606) );
  NOR2X1 U58972 ( .A(n55607), .B(n55606), .Y(n55613) );
  NOR2X1 U58973 ( .A(n42955), .B(n37770), .Y(n55611) );
  NAND2X1 U58974 ( .A(n43256), .B(opcode_pc_w[22]), .Y(n55609) );
  NAND2X1 U58975 ( .A(n43260), .B(n55620), .Y(n55608) );
  NAND2X1 U58976 ( .A(n55609), .B(n55608), .Y(n55610) );
  NOR2X1 U58977 ( .A(n55611), .B(n55610), .Y(n55612) );
  NAND2X1 U58978 ( .A(n55613), .B(n55612), .Y(u_csr_csr_sepc_r[22]) );
  AND2X1 U58979 ( .A(n28334), .B(n28332), .Y(n55618) );
  NOR2X1 U58980 ( .A(n55614), .B(n43293), .Y(n55616) );
  NOR2X1 U58981 ( .A(n58479), .B(n43295), .Y(n55615) );
  NOR2X1 U58982 ( .A(n55616), .B(n55615), .Y(n55617) );
  NAND2X1 U58983 ( .A(n55618), .B(n55617), .Y(u_csr_N3687) );
  NAND2X1 U58984 ( .A(n43299), .B(n55619), .Y(n55622) );
  NAND2X1 U58985 ( .A(n43302), .B(n55620), .Y(n55621) );
  NAND2X1 U58986 ( .A(n55622), .B(n55621), .Y(net2308) );
  INVX1 U58987 ( .A(n17), .Y(n55671) );
  NOR2X1 U58988 ( .A(n55623), .B(n55670), .Y(n55624) );
  XNOR2X1 U58989 ( .A(n55671), .B(n55624), .Y(u_fetch_N71) );
  NOR2X1 U58990 ( .A(n43316), .B(n55628), .Y(net2407) );
  NOR2X1 U58991 ( .A(n43326), .B(n55625), .Y(n55627) );
  NOR2X1 U58992 ( .A(n55627), .B(n55626), .Y(n55632) );
  NOR2X1 U58993 ( .A(n2178), .B(n43321), .Y(n55630) );
  NOR2X1 U58994 ( .A(n43324), .B(n55628), .Y(n55629) );
  NOR2X1 U58995 ( .A(n55630), .B(n55629), .Y(n55631) );
  NAND2X1 U58996 ( .A(n55632), .B(n55631), .Y(u_decode_N312) );
  NAND2X1 U58997 ( .A(n43287), .B(n55667), .Y(n55634) );
  NAND2X1 U58998 ( .A(n43236), .B(n43975), .Y(n55633) );
  NAND2X1 U58999 ( .A(n55634), .B(n55633), .Y(n55639) );
  XNOR2X1 U59000 ( .A(opcode_pc_w[23]), .B(n55683), .Y(n55673) );
  INVX1 U59001 ( .A(n55673), .Y(n55648) );
  NAND2X1 U59002 ( .A(n55648), .B(n43239), .Y(n55637) );
  NAND2X1 U59003 ( .A(n44282), .B(n43979), .Y(n55649) );
  NAND2X1 U59004 ( .A(n27477), .B(n55649), .Y(n55635) );
  NAND2X1 U59005 ( .A(u_csr_csr_mepc_q[23]), .B(n55635), .Y(n55636) );
  NAND2X1 U59006 ( .A(n55637), .B(n55636), .Y(n55638) );
  NOR2X1 U59007 ( .A(n55639), .B(n55638), .Y(n55645) );
  NOR2X1 U59008 ( .A(n42953), .B(n37771), .Y(n55643) );
  NAND2X1 U59009 ( .A(n43243), .B(opcode_pc_w[23]), .Y(n55641) );
  NAND2X1 U59010 ( .A(n43247), .B(n55666), .Y(n55640) );
  NAND2X1 U59011 ( .A(n55641), .B(n55640), .Y(n55642) );
  NOR2X1 U59012 ( .A(n55643), .B(n55642), .Y(n55644) );
  NAND2X1 U59013 ( .A(n55645), .B(n55644), .Y(u_csr_csr_mepc_r[23]) );
  NAND2X1 U59014 ( .A(n43290), .B(n55666), .Y(n55647) );
  NAND2X1 U59015 ( .A(n43253), .B(n43975), .Y(n55646) );
  NAND2X1 U59016 ( .A(n55647), .B(n55646), .Y(n55654) );
  NAND2X1 U59017 ( .A(n55648), .B(n43249), .Y(n55652) );
  NAND2X1 U59018 ( .A(n26373), .B(n55649), .Y(n55650) );
  NAND2X1 U59019 ( .A(u_csr_csr_sepc_q[23]), .B(n55650), .Y(n55651) );
  NAND2X1 U59020 ( .A(n55652), .B(n55651), .Y(n55653) );
  NOR2X1 U59021 ( .A(n55654), .B(n55653), .Y(n55660) );
  NOR2X1 U59022 ( .A(n42957), .B(n37771), .Y(n55658) );
  NAND2X1 U59023 ( .A(n43256), .B(opcode_pc_w[23]), .Y(n55656) );
  NAND2X1 U59024 ( .A(n43260), .B(n55667), .Y(n55655) );
  NAND2X1 U59025 ( .A(n55656), .B(n55655), .Y(n55657) );
  NOR2X1 U59026 ( .A(n55658), .B(n55657), .Y(n55659) );
  NAND2X1 U59027 ( .A(n55660), .B(n55659), .Y(u_csr_csr_sepc_r[23]) );
  AND2X1 U59028 ( .A(n28326), .B(n28324), .Y(n55665) );
  NOR2X1 U59029 ( .A(n55661), .B(n43293), .Y(n55663) );
  NOR2X1 U59030 ( .A(n58480), .B(n43295), .Y(n55662) );
  NOR2X1 U59031 ( .A(n55663), .B(n55662), .Y(n55664) );
  NAND2X1 U59032 ( .A(n55665), .B(n55664), .Y(u_csr_N3688) );
  NAND2X1 U59033 ( .A(n43299), .B(n55666), .Y(n55669) );
  NAND2X1 U59034 ( .A(n43302), .B(n55667), .Y(n55668) );
  NAND2X1 U59035 ( .A(n55669), .B(n55668), .Y(net2309) );
  XNOR2X1 U59036 ( .A(n55672), .B(n42403), .Y(u_fetch_N72) );
  NOR2X1 U59037 ( .A(n43315), .B(n55676), .Y(net2408) );
  NOR2X1 U59038 ( .A(n43326), .B(n55673), .Y(n55675) );
  NOR2X1 U59039 ( .A(n55675), .B(n55674), .Y(n55680) );
  NOR2X1 U59040 ( .A(n2181), .B(n43321), .Y(n55678) );
  NOR2X1 U59041 ( .A(n43324), .B(n55676), .Y(n55677) );
  NOR2X1 U59042 ( .A(n55678), .B(n55677), .Y(n55679) );
  NAND2X1 U59043 ( .A(n55680), .B(n55679), .Y(u_decode_N313) );
  NAND2X1 U59044 ( .A(n43287), .B(n55718), .Y(n55682) );
  NAND2X1 U59045 ( .A(n43236), .B(n43985), .Y(n55681) );
  NAND2X1 U59046 ( .A(n55682), .B(n55681), .Y(n55690) );
  NAND2X1 U59047 ( .A(n55683), .B(opcode_pc_w[23]), .Y(n55684) );
  NAND2X1 U59048 ( .A(n55684), .B(n58370), .Y(n55685) );
  NAND2X1 U59049 ( .A(n55685), .B(n55731), .Y(n55721) );
  INVX1 U59050 ( .A(n55721), .Y(n55699) );
  NAND2X1 U59051 ( .A(n55699), .B(n43239), .Y(n55688) );
  NAND2X1 U59052 ( .A(n44282), .B(n43987), .Y(n55700) );
  NAND2X1 U59053 ( .A(n27477), .B(n55700), .Y(n55686) );
  NAND2X1 U59054 ( .A(u_csr_csr_mepc_q[24]), .B(n55686), .Y(n55687) );
  NAND2X1 U59055 ( .A(n55688), .B(n55687), .Y(n55689) );
  NOR2X1 U59056 ( .A(n55690), .B(n55689), .Y(n55696) );
  NOR2X1 U59057 ( .A(n42951), .B(n37772), .Y(n55694) );
  NAND2X1 U59058 ( .A(n43243), .B(opcode_pc_w[24]), .Y(n55692) );
  NAND2X1 U59059 ( .A(n43247), .B(n55717), .Y(n55691) );
  NAND2X1 U59060 ( .A(n55692), .B(n55691), .Y(n55693) );
  NOR2X1 U59061 ( .A(n55694), .B(n55693), .Y(n55695) );
  NAND2X1 U59062 ( .A(n55696), .B(n55695), .Y(u_csr_csr_mepc_r[24]) );
  NAND2X1 U59063 ( .A(n43290), .B(n55717), .Y(n55698) );
  NAND2X1 U59064 ( .A(n43253), .B(n43985), .Y(n55697) );
  NAND2X1 U59065 ( .A(n55698), .B(n55697), .Y(n55705) );
  NAND2X1 U59066 ( .A(n55699), .B(n43249), .Y(n55703) );
  NAND2X1 U59067 ( .A(n26373), .B(n55700), .Y(n55701) );
  NAND2X1 U59068 ( .A(u_csr_csr_sepc_q[24]), .B(n55701), .Y(n55702) );
  NAND2X1 U59069 ( .A(n55703), .B(n55702), .Y(n55704) );
  NOR2X1 U59070 ( .A(n55705), .B(n55704), .Y(n55711) );
  NOR2X1 U59071 ( .A(n42955), .B(n37772), .Y(n55709) );
  NAND2X1 U59072 ( .A(n43256), .B(opcode_pc_w[24]), .Y(n55707) );
  NAND2X1 U59073 ( .A(n43260), .B(n55718), .Y(n55706) );
  NAND2X1 U59074 ( .A(n55707), .B(n55706), .Y(n55708) );
  NOR2X1 U59075 ( .A(n55709), .B(n55708), .Y(n55710) );
  NAND2X1 U59076 ( .A(n55711), .B(n55710), .Y(u_csr_csr_sepc_r[24]) );
  AND2X1 U59077 ( .A(n28318), .B(n28316), .Y(n55716) );
  NOR2X1 U59078 ( .A(n55712), .B(n43292), .Y(n55714) );
  NOR2X1 U59079 ( .A(n58481), .B(n43295), .Y(n55713) );
  NOR2X1 U59080 ( .A(n55714), .B(n55713), .Y(n55715) );
  NAND2X1 U59081 ( .A(n55716), .B(n55715), .Y(u_csr_N3689) );
  NAND2X1 U59082 ( .A(n43299), .B(n55717), .Y(n55720) );
  NAND2X1 U59083 ( .A(n43302), .B(n55718), .Y(n55719) );
  NAND2X1 U59084 ( .A(n55720), .B(n55719), .Y(net2310) );
  NOR2X1 U59085 ( .A(n43315), .B(n55724), .Y(net2409) );
  NOR2X1 U59086 ( .A(n43326), .B(n55721), .Y(n55723) );
  NOR2X1 U59087 ( .A(n55723), .B(n55722), .Y(n55728) );
  NOR2X1 U59088 ( .A(n2184), .B(n43321), .Y(n55726) );
  NOR2X1 U59089 ( .A(n43324), .B(n55724), .Y(n55725) );
  NOR2X1 U59090 ( .A(n55726), .B(n55725), .Y(n55727) );
  NAND2X1 U59091 ( .A(n55728), .B(n55727), .Y(u_decode_N314) );
  NAND2X1 U59092 ( .A(n43288), .B(n55766), .Y(n55730) );
  NAND2X1 U59093 ( .A(n43236), .B(n43994), .Y(n55729) );
  NAND2X1 U59094 ( .A(n55730), .B(n55729), .Y(n55738) );
  NAND2X1 U59095 ( .A(n55731), .B(n58377), .Y(n55733) );
  NAND2X1 U59096 ( .A(n55733), .B(n55732), .Y(n55769) );
  INVX1 U59097 ( .A(n55769), .Y(n55747) );
  NAND2X1 U59098 ( .A(n55747), .B(n43239), .Y(n55736) );
  NAND2X1 U59099 ( .A(n44282), .B(n43995), .Y(n55748) );
  NAND2X1 U59100 ( .A(n27477), .B(n55748), .Y(n55734) );
  NAND2X1 U59101 ( .A(u_csr_csr_mepc_q[25]), .B(n55734), .Y(n55735) );
  NAND2X1 U59102 ( .A(n55736), .B(n55735), .Y(n55737) );
  NOR2X1 U59103 ( .A(n55738), .B(n55737), .Y(n55744) );
  NOR2X1 U59104 ( .A(n42952), .B(n37773), .Y(n55742) );
  NAND2X1 U59105 ( .A(n43243), .B(opcode_pc_w[25]), .Y(n55740) );
  NAND2X1 U59106 ( .A(n43247), .B(n55765), .Y(n55739) );
  NAND2X1 U59107 ( .A(n55740), .B(n55739), .Y(n55741) );
  NOR2X1 U59108 ( .A(n55742), .B(n55741), .Y(n55743) );
  NAND2X1 U59109 ( .A(n55744), .B(n55743), .Y(u_csr_csr_mepc_r[25]) );
  NAND2X1 U59110 ( .A(n43291), .B(n55765), .Y(n55746) );
  NAND2X1 U59111 ( .A(n43253), .B(n43994), .Y(n55745) );
  NAND2X1 U59112 ( .A(n55746), .B(n55745), .Y(n55753) );
  NAND2X1 U59113 ( .A(n55747), .B(n43249), .Y(n55751) );
  NAND2X1 U59114 ( .A(n26373), .B(n55748), .Y(n55749) );
  NAND2X1 U59115 ( .A(u_csr_csr_sepc_q[25]), .B(n55749), .Y(n55750) );
  NAND2X1 U59116 ( .A(n55751), .B(n55750), .Y(n55752) );
  NOR2X1 U59117 ( .A(n55753), .B(n55752), .Y(n55759) );
  NOR2X1 U59118 ( .A(n42956), .B(n37773), .Y(n55757) );
  NAND2X1 U59119 ( .A(n43256), .B(opcode_pc_w[25]), .Y(n55755) );
  NAND2X1 U59120 ( .A(n43260), .B(n55766), .Y(n55754) );
  NAND2X1 U59121 ( .A(n55755), .B(n55754), .Y(n55756) );
  NOR2X1 U59122 ( .A(n55757), .B(n55756), .Y(n55758) );
  NAND2X1 U59123 ( .A(n55759), .B(n55758), .Y(u_csr_csr_sepc_r[25]) );
  AND2X1 U59124 ( .A(n28310), .B(n28308), .Y(n55764) );
  NOR2X1 U59125 ( .A(n55760), .B(n43292), .Y(n55762) );
  NOR2X1 U59126 ( .A(n58482), .B(n43295), .Y(n55761) );
  NOR2X1 U59127 ( .A(n55762), .B(n55761), .Y(n55763) );
  NAND2X1 U59128 ( .A(n55764), .B(n55763), .Y(u_csr_N3690) );
  NAND2X1 U59129 ( .A(n43300), .B(n55765), .Y(n55768) );
  NAND2X1 U59130 ( .A(n43303), .B(n55766), .Y(n55767) );
  NAND2X1 U59131 ( .A(n55768), .B(n55767), .Y(net2311) );
  NAND2X1 U59132 ( .A(n42413), .B(n11), .Y(n55992) );
  NOR2X1 U59133 ( .A(n43315), .B(n55772), .Y(net2410) );
  NOR2X1 U59134 ( .A(n43326), .B(n55769), .Y(n55771) );
  NOR2X1 U59135 ( .A(n55771), .B(n55770), .Y(n55776) );
  NOR2X1 U59136 ( .A(n2187), .B(n43321), .Y(n55774) );
  NOR2X1 U59137 ( .A(n43324), .B(n55772), .Y(n55773) );
  NOR2X1 U59138 ( .A(n55774), .B(n55773), .Y(n55775) );
  NAND2X1 U59139 ( .A(n55776), .B(n55775), .Y(u_decode_N315) );
  NAND2X1 U59140 ( .A(n43288), .B(n55812), .Y(n55778) );
  NAND2X1 U59141 ( .A(n43236), .B(n44002), .Y(n55777) );
  NAND2X1 U59142 ( .A(n55778), .B(n55777), .Y(n55784) );
  INVX1 U59143 ( .A(n55779), .Y(n55793) );
  NAND2X1 U59144 ( .A(n55793), .B(n43239), .Y(n55782) );
  NAND2X1 U59145 ( .A(n44282), .B(n44005), .Y(n55794) );
  NAND2X1 U59146 ( .A(n27477), .B(n55794), .Y(n55780) );
  NAND2X1 U59147 ( .A(u_csr_csr_mepc_q[26]), .B(n55780), .Y(n55781) );
  NAND2X1 U59148 ( .A(n55782), .B(n55781), .Y(n55783) );
  NOR2X1 U59149 ( .A(n55784), .B(n55783), .Y(n55790) );
  NOR2X1 U59150 ( .A(n42951), .B(n37774), .Y(n55788) );
  NAND2X1 U59151 ( .A(n43243), .B(opcode_pc_w[26]), .Y(n55786) );
  NAND2X1 U59152 ( .A(n43247), .B(n55811), .Y(n55785) );
  NAND2X1 U59153 ( .A(n55786), .B(n55785), .Y(n55787) );
  NOR2X1 U59154 ( .A(n55788), .B(n55787), .Y(n55789) );
  NAND2X1 U59155 ( .A(n55790), .B(n55789), .Y(u_csr_csr_mepc_r[26]) );
  NAND2X1 U59156 ( .A(n43291), .B(n55811), .Y(n55792) );
  NAND2X1 U59157 ( .A(n43253), .B(n44002), .Y(n55791) );
  NAND2X1 U59158 ( .A(n55792), .B(n55791), .Y(n55799) );
  NAND2X1 U59159 ( .A(n55793), .B(n43249), .Y(n55797) );
  NAND2X1 U59160 ( .A(n26373), .B(n55794), .Y(n55795) );
  NAND2X1 U59161 ( .A(u_csr_csr_sepc_q[26]), .B(n55795), .Y(n55796) );
  NAND2X1 U59162 ( .A(n55797), .B(n55796), .Y(n55798) );
  NOR2X1 U59163 ( .A(n55799), .B(n55798), .Y(n55805) );
  NOR2X1 U59164 ( .A(n42955), .B(n37774), .Y(n55803) );
  NAND2X1 U59165 ( .A(n43256), .B(opcode_pc_w[26]), .Y(n55801) );
  NAND2X1 U59166 ( .A(n43260), .B(n55812), .Y(n55800) );
  NAND2X1 U59167 ( .A(n55801), .B(n55800), .Y(n55802) );
  NOR2X1 U59168 ( .A(n55803), .B(n55802), .Y(n55804) );
  NAND2X1 U59169 ( .A(n55805), .B(n55804), .Y(u_csr_csr_sepc_r[26]) );
  AND2X1 U59170 ( .A(n28302), .B(n28300), .Y(n55810) );
  NOR2X1 U59171 ( .A(n55806), .B(n43292), .Y(n55808) );
  NOR2X1 U59172 ( .A(n58483), .B(n43295), .Y(n55807) );
  NOR2X1 U59173 ( .A(n55808), .B(n55807), .Y(n55809) );
  NAND2X1 U59174 ( .A(n55810), .B(n55809), .Y(u_csr_N3691) );
  NAND2X1 U59175 ( .A(n43300), .B(n55811), .Y(n55814) );
  NAND2X1 U59176 ( .A(n43303), .B(n55812), .Y(n55813) );
  NAND2X1 U59177 ( .A(n55814), .B(n55813), .Y(net2312) );
  INVX1 U59178 ( .A(n13), .Y(n55993) );
  NOR2X1 U59179 ( .A(n42409), .B(n55992), .Y(n55815) );
  XNOR2X1 U59180 ( .A(n55993), .B(n55815), .Y(u_fetch_N75) );
  INVX1 U59181 ( .A(n55816), .Y(n55817) );
  MX2X1 U59182 ( .A(n55819), .B(n55818), .S0(n55817), .Y(n56767) );
  INVX1 U59183 ( .A(n56767), .Y(n55820) );
  NOR2X1 U59184 ( .A(n2617), .B(n40672), .Y(n55822) );
  NOR2X1 U59185 ( .A(n8326), .B(n40687), .Y(n55821) );
  NOR2X1 U59186 ( .A(n55822), .B(n55821), .Y(n55824) );
  NAND2X1 U59187 ( .A(n56767), .B(n13), .Y(n55823) );
  NAND2X1 U59188 ( .A(n55824), .B(n55823), .Y(u_mmu_request_addr_w[26]) );
  MX2X1 U59189 ( .A(u_mmu_itlb_va_addr_q[26]), .B(n57389), .S0(n37548), .Y(
        n8433) );
  NOR2X1 U59190 ( .A(n16104), .B(n16105), .Y(n55826) );
  NOR2X1 U59191 ( .A(n16149), .B(n16150), .Y(n55825) );
  NAND2X1 U59192 ( .A(n55826), .B(n55825), .Y(u_exec_alu_p_w[27]) );
  NOR2X1 U59193 ( .A(n44539), .B(n55947), .Y(n55828) );
  NOR2X1 U59194 ( .A(n44537), .B(n43215), .Y(n55827) );
  NOR2X1 U59195 ( .A(n55828), .B(n55827), .Y(n55830) );
  NOR2X1 U59196 ( .A(n19705), .B(n19704), .Y(n55829) );
  NAND2X1 U59197 ( .A(n55830), .B(n55829), .Y(u_decode_u_regfile_N682) );
  NOR2X1 U59198 ( .A(n44603), .B(n55947), .Y(n55832) );
  NOR2X1 U59199 ( .A(n44600), .B(n43215), .Y(n55831) );
  NOR2X1 U59200 ( .A(n55832), .B(n55831), .Y(n55834) );
  NOR2X1 U59201 ( .A(n18118), .B(n18116), .Y(n55833) );
  NAND2X1 U59202 ( .A(n55834), .B(n55833), .Y(u_decode_u_regfile_N978) );
  NOR2X1 U59203 ( .A(n43210), .B(n57131), .Y(n55836) );
  NOR2X1 U59204 ( .A(n43213), .B(n43386), .Y(n55835) );
  NOR2X1 U59205 ( .A(n55836), .B(n55835), .Y(n55838) );
  NOR2X1 U59206 ( .A(n21275), .B(n21274), .Y(n55837) );
  NAND2X1 U59207 ( .A(n55838), .B(n55837), .Y(u_decode_u_regfile_N386) );
  NOR2X1 U59208 ( .A(n44474), .B(n55947), .Y(n55840) );
  NOR2X1 U59209 ( .A(n44471), .B(n43215), .Y(n55839) );
  NOR2X1 U59210 ( .A(n55840), .B(n55839), .Y(n55842) );
  NOR2X1 U59211 ( .A(n20882), .B(n20881), .Y(n55841) );
  NAND2X1 U59212 ( .A(n55842), .B(n55841), .Y(u_decode_u_regfile_N460) );
  NOR2X1 U59213 ( .A(n44561), .B(n55947), .Y(n55844) );
  NOR2X1 U59214 ( .A(n44558), .B(n43215), .Y(n55843) );
  NOR2X1 U59215 ( .A(n55844), .B(n55843), .Y(n55846) );
  NOR2X1 U59216 ( .A(n19310), .B(n19309), .Y(n55845) );
  NAND2X1 U59217 ( .A(n55846), .B(n55845), .Y(u_decode_u_regfile_N756) );
  NOR2X1 U59218 ( .A(n22425), .B(n43211), .Y(n55848) );
  NOR2X1 U59219 ( .A(n44381), .B(n43214), .Y(n55847) );
  NOR2X1 U59220 ( .A(n55848), .B(n55847), .Y(n55850) );
  NOR2X1 U59221 ( .A(n22452), .B(n22451), .Y(n55849) );
  NAND2X1 U59222 ( .A(n55850), .B(n55849), .Y(u_decode_u_regfile_N164) );
  NOR2X1 U59223 ( .A(n23761), .B(n43211), .Y(n55852) );
  NOR2X1 U59224 ( .A(n44303), .B(n43214), .Y(n55851) );
  NOR2X1 U59225 ( .A(n55852), .B(n55851), .Y(n55854) );
  NOR2X1 U59226 ( .A(n23788), .B(n23787), .Y(n55853) );
  NAND2X1 U59227 ( .A(n55854), .B(n55853), .Y(u_decode_u_regfile_N1052) );
  NOR2X1 U59228 ( .A(n44573), .B(n43211), .Y(n55856) );
  NOR2X1 U59229 ( .A(n44570), .B(n43214), .Y(n55855) );
  NOR2X1 U59230 ( .A(n55856), .B(n55855), .Y(n55858) );
  NOR2X1 U59231 ( .A(n18918), .B(n18917), .Y(n55857) );
  NAND2X1 U59232 ( .A(n55858), .B(n55857), .Y(u_decode_u_regfile_N830) );
  NOR2X1 U59233 ( .A(n43210), .B(n57209), .Y(n55860) );
  NOR2X1 U59234 ( .A(n43213), .B(n43383), .Y(n55859) );
  NOR2X1 U59235 ( .A(n55860), .B(n55859), .Y(n55862) );
  NOR2X1 U59236 ( .A(n20490), .B(n20489), .Y(n55861) );
  NAND2X1 U59237 ( .A(n55862), .B(n55861), .Y(u_decode_u_regfile_N534) );
  NOR2X1 U59238 ( .A(n22033), .B(n43211), .Y(n55864) );
  NOR2X1 U59239 ( .A(n44405), .B(n43214), .Y(n55863) );
  NOR2X1 U59240 ( .A(n55864), .B(n55863), .Y(n55866) );
  NOR2X1 U59241 ( .A(n22060), .B(n22059), .Y(n55865) );
  NAND2X1 U59242 ( .A(n55866), .B(n55865), .Y(u_decode_u_regfile_N238) );
  NOR2X1 U59243 ( .A(n23321), .B(n43211), .Y(n55868) );
  NOR2X1 U59244 ( .A(n44327), .B(n43214), .Y(n55867) );
  NOR2X1 U59245 ( .A(n55868), .B(n55867), .Y(n55870) );
  NOR2X1 U59246 ( .A(n23354), .B(n23353), .Y(n55869) );
  NAND2X1 U59247 ( .A(n55870), .B(n55869), .Y(u_decode_u_regfile_N1126) );
  NOR2X1 U59248 ( .A(n44585), .B(n43211), .Y(n55872) );
  NOR2X1 U59249 ( .A(n44582), .B(n43214), .Y(n55871) );
  NOR2X1 U59250 ( .A(n55872), .B(n55871), .Y(n55874) );
  NOR2X1 U59251 ( .A(n18526), .B(n18525), .Y(n55873) );
  NAND2X1 U59252 ( .A(n55874), .B(n55873), .Y(u_decode_u_regfile_N904) );
  NOR2X1 U59253 ( .A(n21641), .B(n43211), .Y(n55876) );
  NOR2X1 U59254 ( .A(n44429), .B(n43214), .Y(n55875) );
  NOR2X1 U59255 ( .A(n55876), .B(n55875), .Y(n55878) );
  NOR2X1 U59256 ( .A(n21668), .B(n21667), .Y(n55877) );
  NAND2X1 U59257 ( .A(n55878), .B(n55877), .Y(u_decode_u_regfile_N312) );
  NOR2X1 U59258 ( .A(n20071), .B(n43211), .Y(n55880) );
  NOR2X1 U59259 ( .A(n44513), .B(n43214), .Y(n55879) );
  NOR2X1 U59260 ( .A(n55880), .B(n55879), .Y(n55882) );
  NOR2X1 U59261 ( .A(n20098), .B(n20097), .Y(n55881) );
  NAND2X1 U59262 ( .A(n55882), .B(n55881), .Y(u_decode_u_regfile_N608) );
  NOR2X1 U59263 ( .A(n22887), .B(n43211), .Y(n55884) );
  NOR2X1 U59264 ( .A(n44351), .B(n43214), .Y(n55883) );
  NOR2X1 U59265 ( .A(n55884), .B(n55883), .Y(n55886) );
  NOR2X1 U59266 ( .A(n22914), .B(n22913), .Y(n55885) );
  NAND2X1 U59267 ( .A(n55886), .B(n55885), .Y(u_decode_u_regfile_N1200) );
  NOR2X1 U59268 ( .A(n18002), .B(n43211), .Y(n55888) );
  NOR2X1 U59269 ( .A(n44606), .B(n43214), .Y(n55887) );
  NOR2X1 U59270 ( .A(n55888), .B(n55887), .Y(n55890) );
  NOR2X1 U59271 ( .A(n24004), .B(n24003), .Y(n55889) );
  NAND2X1 U59272 ( .A(n55890), .B(n55889), .Y(u_decode_u_regfile_N1015) );
  NOR2X1 U59273 ( .A(n43210), .B(n57144), .Y(n55892) );
  NOR2X1 U59274 ( .A(n43213), .B(n43389), .Y(n55891) );
  NOR2X1 U59275 ( .A(n55892), .B(n55891), .Y(n55894) );
  NOR2X1 U59276 ( .A(n22648), .B(n22647), .Y(n55893) );
  NAND2X1 U59277 ( .A(n55894), .B(n55893), .Y(u_decode_u_regfile_N127) );
  NOR2X1 U59278 ( .A(n21051), .B(n43211), .Y(n55896) );
  NOR2X1 U59279 ( .A(n44459), .B(n43214), .Y(n55895) );
  NOR2X1 U59280 ( .A(n55896), .B(n55895), .Y(n55898) );
  NOR2X1 U59281 ( .A(n21078), .B(n21077), .Y(n55897) );
  NAND2X1 U59282 ( .A(n55898), .B(n55897), .Y(u_decode_u_regfile_N423) );
  NOR2X1 U59283 ( .A(n19481), .B(n43211), .Y(n55900) );
  NOR2X1 U59284 ( .A(n44549), .B(n43214), .Y(n55899) );
  NOR2X1 U59285 ( .A(n55900), .B(n55899), .Y(n55902) );
  NOR2X1 U59286 ( .A(n19508), .B(n19507), .Y(n55901) );
  NAND2X1 U59287 ( .A(n55902), .B(n55901), .Y(u_decode_u_regfile_N719) );
  NOR2X1 U59288 ( .A(n19088), .B(n43210), .Y(n55904) );
  NOR2X1 U59289 ( .A(n44564), .B(n43213), .Y(n55903) );
  NOR2X1 U59290 ( .A(n55904), .B(n55903), .Y(n55906) );
  NOR2X1 U59291 ( .A(n19114), .B(n19113), .Y(n55905) );
  NAND2X1 U59292 ( .A(n55906), .B(n55905), .Y(u_decode_u_regfile_N793) );
  NOR2X1 U59293 ( .A(n23541), .B(n43210), .Y(n55908) );
  NOR2X1 U59294 ( .A(n44315), .B(n43213), .Y(n55907) );
  NOR2X1 U59295 ( .A(n55908), .B(n55907), .Y(n55910) );
  NOR2X1 U59296 ( .A(n23574), .B(n23573), .Y(n55909) );
  NAND2X1 U59297 ( .A(n55910), .B(n55909), .Y(u_decode_u_regfile_N1089) );
  NOR2X1 U59298 ( .A(n22229), .B(n43210), .Y(n55912) );
  NOR2X1 U59299 ( .A(n44393), .B(n43213), .Y(n55911) );
  NOR2X1 U59300 ( .A(n55912), .B(n55911), .Y(n55914) );
  NOR2X1 U59301 ( .A(n22256), .B(n22255), .Y(n55913) );
  NAND2X1 U59302 ( .A(n55914), .B(n55913), .Y(u_decode_u_regfile_N201) );
  NOR2X1 U59303 ( .A(n20659), .B(n43210), .Y(n55916) );
  NOR2X1 U59304 ( .A(n44483), .B(n43214), .Y(n55915) );
  NOR2X1 U59305 ( .A(n55916), .B(n55915), .Y(n55918) );
  NOR2X1 U59306 ( .A(n20686), .B(n20685), .Y(n55917) );
  NAND2X1 U59307 ( .A(n55918), .B(n55917), .Y(u_decode_u_regfile_N497) );
  NOR2X1 U59308 ( .A(n21837), .B(n43210), .Y(n55920) );
  NOR2X1 U59309 ( .A(n44417), .B(n43213), .Y(n55919) );
  NOR2X1 U59310 ( .A(n55920), .B(n55919), .Y(n55922) );
  NOR2X1 U59311 ( .A(n21864), .B(n21863), .Y(n55921) );
  NAND2X1 U59312 ( .A(n55922), .B(n55921), .Y(u_decode_u_regfile_N275) );
  NOR2X1 U59313 ( .A(n23107), .B(n43210), .Y(n55924) );
  NOR2X1 U59314 ( .A(n44339), .B(n43213), .Y(n55923) );
  NOR2X1 U59315 ( .A(n55924), .B(n55923), .Y(n55926) );
  NOR2X1 U59316 ( .A(n23134), .B(n23133), .Y(n55925) );
  NAND2X1 U59317 ( .A(n55926), .B(n55925), .Y(u_decode_u_regfile_N1163) );
  NOR2X1 U59318 ( .A(n20267), .B(n43210), .Y(n55928) );
  NOR2X1 U59319 ( .A(n44501), .B(n43213), .Y(n55927) );
  NOR2X1 U59320 ( .A(n55928), .B(n55927), .Y(n55930) );
  NOR2X1 U59321 ( .A(n20294), .B(n20293), .Y(n55929) );
  NAND2X1 U59322 ( .A(n55930), .B(n55929), .Y(u_decode_u_regfile_N571) );
  NOR2X1 U59323 ( .A(n18696), .B(n43210), .Y(n55932) );
  NOR2X1 U59324 ( .A(n44576), .B(n43213), .Y(n55931) );
  NOR2X1 U59325 ( .A(n55932), .B(n55931), .Y(n55934) );
  NOR2X1 U59326 ( .A(n18722), .B(n18721), .Y(n55933) );
  NAND2X1 U59327 ( .A(n55934), .B(n55933), .Y(u_decode_u_regfile_N867) );
  NOR2X1 U59328 ( .A(n19875), .B(n43210), .Y(n55936) );
  NOR2X1 U59329 ( .A(n44525), .B(n43213), .Y(n55935) );
  NOR2X1 U59330 ( .A(n55936), .B(n55935), .Y(n55938) );
  NOR2X1 U59331 ( .A(n19902), .B(n19901), .Y(n55937) );
  NAND2X1 U59332 ( .A(n55938), .B(n55937), .Y(u_decode_u_regfile_N645) );
  NOR2X1 U59333 ( .A(n18305), .B(n43211), .Y(n55940) );
  NOR2X1 U59334 ( .A(n44591), .B(n43213), .Y(n55939) );
  NOR2X1 U59335 ( .A(n55940), .B(n55939), .Y(n55942) );
  NOR2X1 U59336 ( .A(n18332), .B(n18331), .Y(n55941) );
  NAND2X1 U59337 ( .A(n55942), .B(n55941), .Y(u_decode_u_regfile_N941) );
  NOR2X1 U59338 ( .A(n22667), .B(n43210), .Y(n55944) );
  NOR2X1 U59339 ( .A(n44363), .B(n43213), .Y(n55943) );
  NOR2X1 U59340 ( .A(n55944), .B(n55943), .Y(n55946) );
  NOR2X1 U59341 ( .A(n22700), .B(n22699), .Y(n55945) );
  NAND2X1 U59342 ( .A(n55946), .B(n55945), .Y(u_decode_u_regfile_N1237) );
  NOR2X1 U59343 ( .A(n21445), .B(n43211), .Y(n55949) );
  NOR2X1 U59344 ( .A(n44441), .B(n43214), .Y(n55948) );
  NOR2X1 U59345 ( .A(n55949), .B(n55948), .Y(n55951) );
  NOR2X1 U59346 ( .A(n21472), .B(n21471), .Y(n55950) );
  NAND2X1 U59347 ( .A(n55951), .B(n55950), .Y(u_decode_u_regfile_N349) );
  MX2X1 U59348 ( .A(u_csr_pc_m_q[27]), .B(opcode_pc_w[27]), .S0(n58128), .Y(
        n8502) );
  NAND2X1 U59349 ( .A(n43288), .B(n55989), .Y(n55953) );
  NAND2X1 U59350 ( .A(n43236), .B(n44010), .Y(n55952) );
  NAND2X1 U59351 ( .A(n55953), .B(n55952), .Y(n55961) );
  NAND2X1 U59352 ( .A(n55954), .B(n58389), .Y(n55956) );
  INVX1 U59353 ( .A(n55954), .Y(n55955) );
  NAND2X1 U59354 ( .A(n55955), .B(opcode_pc_w[27]), .Y(n56131) );
  NAND2X1 U59355 ( .A(n55956), .B(n56131), .Y(n55994) );
  INVX1 U59356 ( .A(n55994), .Y(n55970) );
  NAND2X1 U59357 ( .A(n55970), .B(n43239), .Y(n55959) );
  NAND2X1 U59358 ( .A(n44282), .B(n44012), .Y(n55971) );
  NAND2X1 U59359 ( .A(n27477), .B(n55971), .Y(n55957) );
  NAND2X1 U59360 ( .A(u_csr_csr_mepc_q[27]), .B(n55957), .Y(n55958) );
  NAND2X1 U59361 ( .A(n55959), .B(n55958), .Y(n55960) );
  NOR2X1 U59362 ( .A(n55961), .B(n55960), .Y(n55967) );
  NOR2X1 U59363 ( .A(n42952), .B(n37757), .Y(n55965) );
  NAND2X1 U59364 ( .A(n43243), .B(opcode_pc_w[27]), .Y(n55963) );
  NAND2X1 U59365 ( .A(n43248), .B(n55988), .Y(n55962) );
  NAND2X1 U59366 ( .A(n55963), .B(n55962), .Y(n55964) );
  NOR2X1 U59367 ( .A(n55965), .B(n55964), .Y(n55966) );
  NAND2X1 U59368 ( .A(n55967), .B(n55966), .Y(u_csr_csr_mepc_r[27]) );
  NAND2X1 U59369 ( .A(n43291), .B(n55988), .Y(n55969) );
  NAND2X1 U59370 ( .A(n43253), .B(n44010), .Y(n55968) );
  NAND2X1 U59371 ( .A(n55969), .B(n55968), .Y(n55976) );
  NAND2X1 U59372 ( .A(n55970), .B(n43249), .Y(n55974) );
  NAND2X1 U59373 ( .A(n26373), .B(n55971), .Y(n55972) );
  NAND2X1 U59374 ( .A(u_csr_csr_sepc_q[27]), .B(n55972), .Y(n55973) );
  NAND2X1 U59375 ( .A(n55974), .B(n55973), .Y(n55975) );
  NOR2X1 U59376 ( .A(n55976), .B(n55975), .Y(n55982) );
  NOR2X1 U59377 ( .A(n42956), .B(n37757), .Y(n55980) );
  NAND2X1 U59378 ( .A(n43256), .B(opcode_pc_w[27]), .Y(n55978) );
  NAND2X1 U59379 ( .A(n56600), .B(n55989), .Y(n55977) );
  NAND2X1 U59380 ( .A(n55978), .B(n55977), .Y(n55979) );
  NOR2X1 U59381 ( .A(n55980), .B(n55979), .Y(n55981) );
  NAND2X1 U59382 ( .A(n55982), .B(n55981), .Y(u_csr_csr_sepc_r[27]) );
  AND2X1 U59383 ( .A(n28294), .B(n28292), .Y(n55987) );
  NOR2X1 U59384 ( .A(n55983), .B(n43292), .Y(n55985) );
  NOR2X1 U59385 ( .A(n58484), .B(n43295), .Y(n55984) );
  NOR2X1 U59386 ( .A(n55985), .B(n55984), .Y(n55986) );
  NAND2X1 U59387 ( .A(n55987), .B(n55986), .Y(u_csr_N3692) );
  NAND2X1 U59388 ( .A(n43300), .B(n55988), .Y(n55991) );
  NAND2X1 U59389 ( .A(n43303), .B(n55989), .Y(n55990) );
  NAND2X1 U59390 ( .A(n55991), .B(n55990), .Y(net2313) );
  NOR2X1 U59391 ( .A(n43315), .B(n55997), .Y(net2412) );
  NOR2X1 U59392 ( .A(n43327), .B(n55994), .Y(n55996) );
  NOR2X1 U59393 ( .A(n55996), .B(n55995), .Y(n56001) );
  NOR2X1 U59394 ( .A(n1939), .B(n43321), .Y(n55999) );
  NOR2X1 U59395 ( .A(n43324), .B(n55997), .Y(n55998) );
  NOR2X1 U59396 ( .A(n55999), .B(n55998), .Y(n56000) );
  NAND2X1 U59397 ( .A(n56001), .B(n56000), .Y(u_decode_N317) );
  NOR2X1 U59398 ( .A(n16028), .B(n16029), .Y(n56003) );
  NOR2X1 U59399 ( .A(n16085), .B(n16086), .Y(n56002) );
  NAND2X1 U59400 ( .A(n56003), .B(n56002), .Y(u_exec_alu_p_w[28]) );
  NOR2X1 U59401 ( .A(n44539), .B(n56124), .Y(n56005) );
  NOR2X1 U59402 ( .A(n44537), .B(n37685), .Y(n56004) );
  NOR2X1 U59403 ( .A(n56005), .B(n56004), .Y(n56007) );
  NOR2X1 U59404 ( .A(n19699), .B(n19698), .Y(n56006) );
  NAND2X1 U59405 ( .A(n56007), .B(n56006), .Y(u_decode_u_regfile_N683) );
  NOR2X1 U59406 ( .A(n44603), .B(n56124), .Y(n56009) );
  NOR2X1 U59407 ( .A(n44600), .B(n37685), .Y(n56008) );
  NOR2X1 U59408 ( .A(n56009), .B(n56008), .Y(n56011) );
  NOR2X1 U59409 ( .A(n18111), .B(n18109), .Y(n56010) );
  NAND2X1 U59410 ( .A(n56011), .B(n56010), .Y(u_decode_u_regfile_N979) );
  NOR2X1 U59411 ( .A(n43217), .B(n57131), .Y(n56013) );
  NOR2X1 U59412 ( .A(n43220), .B(n43386), .Y(n56012) );
  NOR2X1 U59413 ( .A(n56013), .B(n56012), .Y(n56015) );
  NOR2X1 U59414 ( .A(n21269), .B(n21268), .Y(n56014) );
  NAND2X1 U59415 ( .A(n56015), .B(n56014), .Y(u_decode_u_regfile_N387) );
  NOR2X1 U59416 ( .A(n44474), .B(n56124), .Y(n56017) );
  NOR2X1 U59417 ( .A(n44471), .B(n37685), .Y(n56016) );
  NOR2X1 U59418 ( .A(n56017), .B(n56016), .Y(n56019) );
  NOR2X1 U59419 ( .A(n20876), .B(n20875), .Y(n56018) );
  NAND2X1 U59420 ( .A(n56019), .B(n56018), .Y(u_decode_u_regfile_N461) );
  NOR2X1 U59421 ( .A(n44561), .B(n56124), .Y(n56021) );
  NOR2X1 U59422 ( .A(n44558), .B(n37685), .Y(n56020) );
  NOR2X1 U59423 ( .A(n56021), .B(n56020), .Y(n56023) );
  NOR2X1 U59424 ( .A(n19304), .B(n19303), .Y(n56022) );
  NAND2X1 U59425 ( .A(n56023), .B(n56022), .Y(u_decode_u_regfile_N757) );
  NOR2X1 U59426 ( .A(n22425), .B(n43218), .Y(n56025) );
  NOR2X1 U59427 ( .A(n44381), .B(n43221), .Y(n56024) );
  NOR2X1 U59428 ( .A(n56025), .B(n56024), .Y(n56027) );
  NOR2X1 U59429 ( .A(n22446), .B(n22445), .Y(n56026) );
  NAND2X1 U59430 ( .A(n56027), .B(n56026), .Y(u_decode_u_regfile_N165) );
  NOR2X1 U59431 ( .A(n23761), .B(n43218), .Y(n56029) );
  NOR2X1 U59432 ( .A(n44303), .B(n43221), .Y(n56028) );
  NOR2X1 U59433 ( .A(n56029), .B(n56028), .Y(n56031) );
  NOR2X1 U59434 ( .A(n23782), .B(n23781), .Y(n56030) );
  NAND2X1 U59435 ( .A(n56031), .B(n56030), .Y(u_decode_u_regfile_N1053) );
  NOR2X1 U59436 ( .A(n44573), .B(n43218), .Y(n56033) );
  NOR2X1 U59437 ( .A(n44570), .B(n43221), .Y(n56032) );
  NOR2X1 U59438 ( .A(n56033), .B(n56032), .Y(n56035) );
  NOR2X1 U59439 ( .A(n18912), .B(n18911), .Y(n56034) );
  NAND2X1 U59440 ( .A(n56035), .B(n56034), .Y(u_decode_u_regfile_N831) );
  NOR2X1 U59441 ( .A(n43217), .B(n57209), .Y(n56037) );
  NOR2X1 U59442 ( .A(n43220), .B(n43383), .Y(n56036) );
  NOR2X1 U59443 ( .A(n56037), .B(n56036), .Y(n56039) );
  NOR2X1 U59444 ( .A(n20484), .B(n20483), .Y(n56038) );
  NAND2X1 U59445 ( .A(n56039), .B(n56038), .Y(u_decode_u_regfile_N535) );
  NOR2X1 U59446 ( .A(n22033), .B(n43218), .Y(n56041) );
  NOR2X1 U59447 ( .A(n44405), .B(n43221), .Y(n56040) );
  NOR2X1 U59448 ( .A(n56041), .B(n56040), .Y(n56043) );
  NOR2X1 U59449 ( .A(n22054), .B(n22053), .Y(n56042) );
  NAND2X1 U59450 ( .A(n56043), .B(n56042), .Y(u_decode_u_regfile_N239) );
  NOR2X1 U59451 ( .A(n23321), .B(n43218), .Y(n56045) );
  NOR2X1 U59452 ( .A(n44327), .B(n43221), .Y(n56044) );
  NOR2X1 U59453 ( .A(n56045), .B(n56044), .Y(n56047) );
  NOR2X1 U59454 ( .A(n23348), .B(n23347), .Y(n56046) );
  NAND2X1 U59455 ( .A(n56047), .B(n56046), .Y(u_decode_u_regfile_N1127) );
  NOR2X1 U59456 ( .A(n44585), .B(n43218), .Y(n56049) );
  NOR2X1 U59457 ( .A(n44582), .B(n43221), .Y(n56048) );
  NOR2X1 U59458 ( .A(n56049), .B(n56048), .Y(n56051) );
  NOR2X1 U59459 ( .A(n18520), .B(n18519), .Y(n56050) );
  NAND2X1 U59460 ( .A(n56051), .B(n56050), .Y(u_decode_u_regfile_N905) );
  NOR2X1 U59461 ( .A(n21641), .B(n43218), .Y(n56053) );
  NOR2X1 U59462 ( .A(n44429), .B(n43221), .Y(n56052) );
  NOR2X1 U59463 ( .A(n56053), .B(n56052), .Y(n56055) );
  NOR2X1 U59464 ( .A(n21662), .B(n21661), .Y(n56054) );
  NAND2X1 U59465 ( .A(n56055), .B(n56054), .Y(u_decode_u_regfile_N313) );
  NOR2X1 U59466 ( .A(n20071), .B(n43218), .Y(n56057) );
  NOR2X1 U59467 ( .A(n44513), .B(n43221), .Y(n56056) );
  NOR2X1 U59468 ( .A(n56057), .B(n56056), .Y(n56059) );
  NOR2X1 U59469 ( .A(n20092), .B(n20091), .Y(n56058) );
  NAND2X1 U59470 ( .A(n56059), .B(n56058), .Y(u_decode_u_regfile_N609) );
  NOR2X1 U59471 ( .A(n22887), .B(n43218), .Y(n56061) );
  NOR2X1 U59472 ( .A(n44351), .B(n43221), .Y(n56060) );
  NOR2X1 U59473 ( .A(n56061), .B(n56060), .Y(n56063) );
  NOR2X1 U59474 ( .A(n22908), .B(n22907), .Y(n56062) );
  NAND2X1 U59475 ( .A(n56063), .B(n56062), .Y(u_decode_u_regfile_N1201) );
  NOR2X1 U59476 ( .A(n18002), .B(n43218), .Y(n56065) );
  NOR2X1 U59477 ( .A(n44606), .B(n43221), .Y(n56064) );
  NOR2X1 U59478 ( .A(n56065), .B(n56064), .Y(n56067) );
  NOR2X1 U59479 ( .A(n23998), .B(n23997), .Y(n56066) );
  NAND2X1 U59480 ( .A(n56067), .B(n56066), .Y(u_decode_u_regfile_N1016) );
  NOR2X1 U59481 ( .A(n43217), .B(n57144), .Y(n56069) );
  NOR2X1 U59482 ( .A(n43220), .B(n43389), .Y(n56068) );
  NOR2X1 U59483 ( .A(n56069), .B(n56068), .Y(n56071) );
  NOR2X1 U59484 ( .A(n22642), .B(n22641), .Y(n56070) );
  NAND2X1 U59485 ( .A(n56071), .B(n56070), .Y(u_decode_u_regfile_N128) );
  NOR2X1 U59486 ( .A(n21051), .B(n43218), .Y(n56073) );
  NOR2X1 U59487 ( .A(n44459), .B(n43221), .Y(n56072) );
  NOR2X1 U59488 ( .A(n56073), .B(n56072), .Y(n56075) );
  NOR2X1 U59489 ( .A(n21072), .B(n21071), .Y(n56074) );
  NAND2X1 U59490 ( .A(n56075), .B(n56074), .Y(u_decode_u_regfile_N424) );
  NOR2X1 U59491 ( .A(n19481), .B(n43218), .Y(n56077) );
  NOR2X1 U59492 ( .A(n44549), .B(n43221), .Y(n56076) );
  NOR2X1 U59493 ( .A(n56077), .B(n56076), .Y(n56079) );
  NOR2X1 U59494 ( .A(n19502), .B(n19501), .Y(n56078) );
  NAND2X1 U59495 ( .A(n56079), .B(n56078), .Y(u_decode_u_regfile_N720) );
  NOR2X1 U59496 ( .A(n44565), .B(n43217), .Y(n56081) );
  NOR2X1 U59497 ( .A(n44564), .B(n43220), .Y(n56080) );
  NOR2X1 U59498 ( .A(n56081), .B(n56080), .Y(n56083) );
  NOR2X1 U59499 ( .A(n19108), .B(n19107), .Y(n56082) );
  NAND2X1 U59500 ( .A(n56083), .B(n56082), .Y(u_decode_u_regfile_N794) );
  NOR2X1 U59501 ( .A(n23541), .B(n43217), .Y(n56085) );
  NOR2X1 U59502 ( .A(n44315), .B(n43220), .Y(n56084) );
  NOR2X1 U59503 ( .A(n56085), .B(n56084), .Y(n56087) );
  NOR2X1 U59504 ( .A(n23562), .B(n23561), .Y(n56086) );
  NAND2X1 U59505 ( .A(n56087), .B(n56086), .Y(u_decode_u_regfile_N1090) );
  NOR2X1 U59506 ( .A(n22229), .B(n43217), .Y(n56089) );
  NOR2X1 U59507 ( .A(n44393), .B(n43220), .Y(n56088) );
  NOR2X1 U59508 ( .A(n56089), .B(n56088), .Y(n56091) );
  NOR2X1 U59509 ( .A(n22250), .B(n22249), .Y(n56090) );
  NAND2X1 U59510 ( .A(n56091), .B(n56090), .Y(u_decode_u_regfile_N202) );
  NOR2X1 U59511 ( .A(n20659), .B(n43217), .Y(n56093) );
  NOR2X1 U59512 ( .A(n44483), .B(n43220), .Y(n56092) );
  NOR2X1 U59513 ( .A(n56093), .B(n56092), .Y(n56095) );
  NOR2X1 U59514 ( .A(n20680), .B(n20679), .Y(n56094) );
  NAND2X1 U59515 ( .A(n56095), .B(n56094), .Y(u_decode_u_regfile_N498) );
  NOR2X1 U59516 ( .A(n44419), .B(n43217), .Y(n56097) );
  NOR2X1 U59517 ( .A(n44417), .B(n43220), .Y(n56096) );
  NOR2X1 U59518 ( .A(n56097), .B(n56096), .Y(n56099) );
  NOR2X1 U59519 ( .A(n21858), .B(n21857), .Y(n56098) );
  NAND2X1 U59520 ( .A(n56099), .B(n56098), .Y(u_decode_u_regfile_N276) );
  NOR2X1 U59521 ( .A(n23107), .B(n43217), .Y(n56101) );
  NOR2X1 U59522 ( .A(n44339), .B(n43220), .Y(n56100) );
  NOR2X1 U59523 ( .A(n56101), .B(n56100), .Y(n56103) );
  NOR2X1 U59524 ( .A(n23128), .B(n23127), .Y(n56102) );
  NAND2X1 U59525 ( .A(n56103), .B(n56102), .Y(u_decode_u_regfile_N1164) );
  NOR2X1 U59526 ( .A(n20267), .B(n43217), .Y(n56105) );
  NOR2X1 U59527 ( .A(n44501), .B(n43220), .Y(n56104) );
  NOR2X1 U59528 ( .A(n56105), .B(n56104), .Y(n56107) );
  NOR2X1 U59529 ( .A(n20288), .B(n20287), .Y(n56106) );
  NAND2X1 U59530 ( .A(n56107), .B(n56106), .Y(u_decode_u_regfile_N572) );
  NOR2X1 U59531 ( .A(n44578), .B(n43217), .Y(n56109) );
  NOR2X1 U59532 ( .A(n44576), .B(n43220), .Y(n56108) );
  NOR2X1 U59533 ( .A(n56109), .B(n56108), .Y(n56111) );
  NOR2X1 U59534 ( .A(n18716), .B(n18715), .Y(n56110) );
  NAND2X1 U59535 ( .A(n56111), .B(n56110), .Y(u_decode_u_regfile_N868) );
  NOR2X1 U59536 ( .A(n19875), .B(n43217), .Y(n56113) );
  NOR2X1 U59537 ( .A(n44525), .B(n43220), .Y(n56112) );
  NOR2X1 U59538 ( .A(n56113), .B(n56112), .Y(n56115) );
  NOR2X1 U59539 ( .A(n19896), .B(n19895), .Y(n56114) );
  NAND2X1 U59540 ( .A(n56115), .B(n56114), .Y(u_decode_u_regfile_N646) );
  NOR2X1 U59541 ( .A(n18305), .B(n43218), .Y(n56117) );
  NOR2X1 U59542 ( .A(n44591), .B(n43221), .Y(n56116) );
  NOR2X1 U59543 ( .A(n56117), .B(n56116), .Y(n56119) );
  NOR2X1 U59544 ( .A(n18326), .B(n18325), .Y(n56118) );
  NAND2X1 U59545 ( .A(n56119), .B(n56118), .Y(u_decode_u_regfile_N942) );
  NOR2X1 U59546 ( .A(n22667), .B(n43217), .Y(n56121) );
  NOR2X1 U59547 ( .A(n44363), .B(n43220), .Y(n56120) );
  NOR2X1 U59548 ( .A(n56121), .B(n56120), .Y(n56123) );
  NOR2X1 U59549 ( .A(n22694), .B(n22693), .Y(n56122) );
  NAND2X1 U59550 ( .A(n56123), .B(n56122), .Y(u_decode_u_regfile_N1238) );
  NOR2X1 U59551 ( .A(n21445), .B(n43218), .Y(n56126) );
  NOR2X1 U59552 ( .A(n44441), .B(n43221), .Y(n56125) );
  NOR2X1 U59553 ( .A(n56126), .B(n56125), .Y(n56128) );
  NOR2X1 U59554 ( .A(n21466), .B(n21465), .Y(n56127) );
  NAND2X1 U59555 ( .A(n56128), .B(n56127), .Y(u_decode_u_regfile_N350) );
  MX2X1 U59556 ( .A(u_csr_pc_m_q[28]), .B(opcode_pc_w[28]), .S0(n58128), .Y(
        n8501) );
  NAND2X1 U59557 ( .A(n43288), .B(n56166), .Y(n56130) );
  NAND2X1 U59558 ( .A(n43236), .B(n44019), .Y(n56129) );
  NAND2X1 U59559 ( .A(n56130), .B(n56129), .Y(n56138) );
  NAND2X1 U59560 ( .A(n56131), .B(n58396), .Y(n56133) );
  INVX1 U59561 ( .A(n56131), .Y(n56132) );
  NAND2X1 U59562 ( .A(n56132), .B(opcode_pc_w[28]), .Y(n56178) );
  NAND2X1 U59563 ( .A(n56133), .B(n56178), .Y(n56170) );
  INVX1 U59564 ( .A(n56170), .Y(n56147) );
  NAND2X1 U59565 ( .A(n56147), .B(n43239), .Y(n56136) );
  NAND2X1 U59566 ( .A(n44282), .B(n44021), .Y(n56148) );
  NAND2X1 U59567 ( .A(n27477), .B(n56148), .Y(n56134) );
  NAND2X1 U59568 ( .A(u_csr_csr_mepc_q[28]), .B(n56134), .Y(n56135) );
  NAND2X1 U59569 ( .A(n56136), .B(n56135), .Y(n56137) );
  NOR2X1 U59570 ( .A(n56138), .B(n56137), .Y(n56144) );
  NOR2X1 U59571 ( .A(n42951), .B(n37758), .Y(n56142) );
  NAND2X1 U59572 ( .A(n43243), .B(opcode_pc_w[28]), .Y(n56140) );
  NAND2X1 U59573 ( .A(n43248), .B(n56165), .Y(n56139) );
  NAND2X1 U59574 ( .A(n56140), .B(n56139), .Y(n56141) );
  NOR2X1 U59575 ( .A(n56142), .B(n56141), .Y(n56143) );
  NAND2X1 U59576 ( .A(n56144), .B(n56143), .Y(u_csr_csr_mepc_r[28]) );
  NAND2X1 U59577 ( .A(n43291), .B(n56165), .Y(n56146) );
  NAND2X1 U59578 ( .A(n43253), .B(n44019), .Y(n56145) );
  NAND2X1 U59579 ( .A(n56146), .B(n56145), .Y(n56153) );
  NAND2X1 U59580 ( .A(n56147), .B(n43249), .Y(n56151) );
  NAND2X1 U59581 ( .A(n26373), .B(n56148), .Y(n56149) );
  NAND2X1 U59582 ( .A(u_csr_csr_sepc_q[28]), .B(n56149), .Y(n56150) );
  NAND2X1 U59583 ( .A(n56151), .B(n56150), .Y(n56152) );
  NOR2X1 U59584 ( .A(n56153), .B(n56152), .Y(n56159) );
  NOR2X1 U59585 ( .A(n42955), .B(n37758), .Y(n56157) );
  NAND2X1 U59586 ( .A(n43256), .B(opcode_pc_w[28]), .Y(n56155) );
  NAND2X1 U59587 ( .A(n56600), .B(n56166), .Y(n56154) );
  NAND2X1 U59588 ( .A(n56155), .B(n56154), .Y(n56156) );
  NOR2X1 U59589 ( .A(n56157), .B(n56156), .Y(n56158) );
  NAND2X1 U59590 ( .A(n56159), .B(n56158), .Y(u_csr_csr_sepc_r[28]) );
  AND2X1 U59591 ( .A(n28286), .B(n28284), .Y(n56164) );
  NOR2X1 U59592 ( .A(n56160), .B(n43292), .Y(n56162) );
  NOR2X1 U59593 ( .A(n58485), .B(n43295), .Y(n56161) );
  NOR2X1 U59594 ( .A(n56162), .B(n56161), .Y(n56163) );
  NAND2X1 U59595 ( .A(n56164), .B(n56163), .Y(u_csr_N3693) );
  NAND2X1 U59596 ( .A(n43300), .B(n56165), .Y(n56168) );
  NAND2X1 U59597 ( .A(n43303), .B(n56166), .Y(n56167) );
  NAND2X1 U59598 ( .A(n56168), .B(n56167), .Y(net2314) );
  XNOR2X1 U59599 ( .A(n56169), .B(n42411), .Y(u_fetch_N77) );
  NOR2X1 U59600 ( .A(n43315), .B(n56173), .Y(net2413) );
  NOR2X1 U59601 ( .A(n43326), .B(n56170), .Y(n56172) );
  NOR2X1 U59602 ( .A(n56172), .B(n56171), .Y(n56177) );
  NOR2X1 U59603 ( .A(n1937), .B(n43322), .Y(n56175) );
  NOR2X1 U59604 ( .A(n43325), .B(n56173), .Y(n56174) );
  NOR2X1 U59605 ( .A(n56175), .B(n56174), .Y(n56176) );
  NAND2X1 U59606 ( .A(n56177), .B(n56176), .Y(u_decode_N318) );
  NOR2X1 U59607 ( .A(n43315), .B(n56183), .Y(net2414) );
  NAND2X1 U59608 ( .A(n56178), .B(n58403), .Y(n56180) );
  INVX1 U59609 ( .A(n56178), .Y(n56179) );
  NAND2X1 U59610 ( .A(n56179), .B(opcode_pc_w[29]), .Y(n56566) );
  NAND2X1 U59611 ( .A(n56180), .B(n56566), .Y(n56316) );
  NOR2X1 U59612 ( .A(n43326), .B(n56316), .Y(n56182) );
  NOR2X1 U59613 ( .A(n56182), .B(n56181), .Y(n56187) );
  NOR2X1 U59614 ( .A(n1935), .B(n43322), .Y(n56185) );
  NOR2X1 U59615 ( .A(n43325), .B(n56183), .Y(n56184) );
  NOR2X1 U59616 ( .A(n56185), .B(n56184), .Y(n56186) );
  NAND2X1 U59617 ( .A(n56187), .B(n56186), .Y(u_decode_N319) );
  NOR2X1 U59618 ( .A(n15953), .B(n15954), .Y(n56189) );
  NOR2X1 U59619 ( .A(n16013), .B(n16014), .Y(n56188) );
  NAND2X1 U59620 ( .A(n56189), .B(n56188), .Y(u_exec_alu_p_w[29]) );
  NOR2X1 U59621 ( .A(n44539), .B(n43225), .Y(n56191) );
  NOR2X1 U59622 ( .A(n44537), .B(n37686), .Y(n56190) );
  NOR2X1 U59623 ( .A(n56191), .B(n56190), .Y(n56193) );
  NOR2X1 U59624 ( .A(n19693), .B(n19692), .Y(n56192) );
  NAND2X1 U59625 ( .A(n56193), .B(n56192), .Y(u_decode_u_regfile_N684) );
  NOR2X1 U59626 ( .A(n44603), .B(n43225), .Y(n56195) );
  NOR2X1 U59627 ( .A(n44600), .B(n37686), .Y(n56194) );
  NOR2X1 U59628 ( .A(n56195), .B(n56194), .Y(n56197) );
  NOR2X1 U59629 ( .A(n18104), .B(n18102), .Y(n56196) );
  NAND2X1 U59630 ( .A(n56197), .B(n56196), .Y(u_decode_u_regfile_N980) );
  NOR2X1 U59631 ( .A(n43223), .B(n57131), .Y(n56199) );
  NOR2X1 U59632 ( .A(n43226), .B(n43386), .Y(n56198) );
  NOR2X1 U59633 ( .A(n56199), .B(n56198), .Y(n56201) );
  NOR2X1 U59634 ( .A(n21263), .B(n21262), .Y(n56200) );
  NAND2X1 U59635 ( .A(n56201), .B(n56200), .Y(u_decode_u_regfile_N388) );
  NOR2X1 U59636 ( .A(n44474), .B(n43225), .Y(n56203) );
  NOR2X1 U59637 ( .A(n44471), .B(n37686), .Y(n56202) );
  NOR2X1 U59638 ( .A(n56203), .B(n56202), .Y(n56205) );
  NOR2X1 U59639 ( .A(n20870), .B(n20869), .Y(n56204) );
  NAND2X1 U59640 ( .A(n56205), .B(n56204), .Y(u_decode_u_regfile_N462) );
  NOR2X1 U59641 ( .A(n44561), .B(n43225), .Y(n56207) );
  NOR2X1 U59642 ( .A(n44558), .B(n37686), .Y(n56206) );
  NOR2X1 U59643 ( .A(n56207), .B(n56206), .Y(n56209) );
  NOR2X1 U59644 ( .A(n19298), .B(n19297), .Y(n56208) );
  NAND2X1 U59645 ( .A(n56209), .B(n56208), .Y(u_decode_u_regfile_N758) );
  NOR2X1 U59646 ( .A(n22425), .B(n43224), .Y(n56211) );
  NOR2X1 U59647 ( .A(n44381), .B(n43227), .Y(n56210) );
  NOR2X1 U59648 ( .A(n56211), .B(n56210), .Y(n56213) );
  NOR2X1 U59649 ( .A(n22440), .B(n22439), .Y(n56212) );
  NAND2X1 U59650 ( .A(n56213), .B(n56212), .Y(u_decode_u_regfile_N166) );
  NOR2X1 U59651 ( .A(n23761), .B(n43224), .Y(n56215) );
  NOR2X1 U59652 ( .A(n44303), .B(n43227), .Y(n56214) );
  NOR2X1 U59653 ( .A(n56215), .B(n56214), .Y(n56217) );
  NOR2X1 U59654 ( .A(n23776), .B(n23775), .Y(n56216) );
  NAND2X1 U59655 ( .A(n56217), .B(n56216), .Y(u_decode_u_regfile_N1054) );
  NOR2X1 U59656 ( .A(n44573), .B(n43224), .Y(n56219) );
  NOR2X1 U59657 ( .A(n44570), .B(n43227), .Y(n56218) );
  NOR2X1 U59658 ( .A(n56219), .B(n56218), .Y(n56221) );
  NOR2X1 U59659 ( .A(n18906), .B(n18905), .Y(n56220) );
  NAND2X1 U59660 ( .A(n56221), .B(n56220), .Y(u_decode_u_regfile_N832) );
  NOR2X1 U59661 ( .A(n43223), .B(n57209), .Y(n56223) );
  NOR2X1 U59662 ( .A(n43226), .B(n43383), .Y(n56222) );
  NOR2X1 U59663 ( .A(n56223), .B(n56222), .Y(n56225) );
  NOR2X1 U59664 ( .A(n20478), .B(n20477), .Y(n56224) );
  NAND2X1 U59665 ( .A(n56225), .B(n56224), .Y(u_decode_u_regfile_N536) );
  NOR2X1 U59666 ( .A(n22033), .B(n43224), .Y(n56227) );
  NOR2X1 U59667 ( .A(n44405), .B(n43227), .Y(n56226) );
  NOR2X1 U59668 ( .A(n56227), .B(n56226), .Y(n56229) );
  NOR2X1 U59669 ( .A(n22048), .B(n22047), .Y(n56228) );
  NAND2X1 U59670 ( .A(n56229), .B(n56228), .Y(u_decode_u_regfile_N240) );
  NOR2X1 U59671 ( .A(n23321), .B(n43224), .Y(n56231) );
  NOR2X1 U59672 ( .A(n44327), .B(n43227), .Y(n56230) );
  NOR2X1 U59673 ( .A(n56231), .B(n56230), .Y(n56233) );
  NOR2X1 U59674 ( .A(n23342), .B(n23341), .Y(n56232) );
  NAND2X1 U59675 ( .A(n56233), .B(n56232), .Y(u_decode_u_regfile_N1128) );
  NOR2X1 U59676 ( .A(n44585), .B(n43224), .Y(n56235) );
  NOR2X1 U59677 ( .A(n44582), .B(n43227), .Y(n56234) );
  NOR2X1 U59678 ( .A(n56235), .B(n56234), .Y(n56237) );
  NOR2X1 U59679 ( .A(n18514), .B(n18513), .Y(n56236) );
  NAND2X1 U59680 ( .A(n56237), .B(n56236), .Y(u_decode_u_regfile_N906) );
  NOR2X1 U59681 ( .A(n21641), .B(n43224), .Y(n56239) );
  NOR2X1 U59682 ( .A(n44429), .B(n43227), .Y(n56238) );
  NOR2X1 U59683 ( .A(n56239), .B(n56238), .Y(n56241) );
  NOR2X1 U59684 ( .A(n21656), .B(n21655), .Y(n56240) );
  NAND2X1 U59685 ( .A(n56241), .B(n56240), .Y(u_decode_u_regfile_N314) );
  NOR2X1 U59686 ( .A(n20071), .B(n43224), .Y(n56243) );
  NOR2X1 U59687 ( .A(n44513), .B(n43227), .Y(n56242) );
  NOR2X1 U59688 ( .A(n56243), .B(n56242), .Y(n56245) );
  NOR2X1 U59689 ( .A(n20086), .B(n20085), .Y(n56244) );
  NAND2X1 U59690 ( .A(n56245), .B(n56244), .Y(u_decode_u_regfile_N610) );
  NOR2X1 U59691 ( .A(n22887), .B(n43224), .Y(n56247) );
  NOR2X1 U59692 ( .A(n44351), .B(n43227), .Y(n56246) );
  NOR2X1 U59693 ( .A(n56247), .B(n56246), .Y(n56249) );
  NOR2X1 U59694 ( .A(n22902), .B(n22901), .Y(n56248) );
  NAND2X1 U59695 ( .A(n56249), .B(n56248), .Y(u_decode_u_regfile_N1202) );
  NOR2X1 U59696 ( .A(n18002), .B(n43224), .Y(n56251) );
  NOR2X1 U59697 ( .A(n44606), .B(n43227), .Y(n56250) );
  NOR2X1 U59698 ( .A(n56251), .B(n56250), .Y(n56253) );
  NOR2X1 U59699 ( .A(n23992), .B(n23991), .Y(n56252) );
  NAND2X1 U59700 ( .A(n56253), .B(n56252), .Y(u_decode_u_regfile_N1017) );
  NOR2X1 U59701 ( .A(n43223), .B(n57144), .Y(n56255) );
  NOR2X1 U59702 ( .A(n43226), .B(n43389), .Y(n56254) );
  NOR2X1 U59703 ( .A(n56255), .B(n56254), .Y(n56257) );
  NOR2X1 U59704 ( .A(n22636), .B(n22635), .Y(n56256) );
  NAND2X1 U59705 ( .A(n56257), .B(n56256), .Y(u_decode_u_regfile_N129) );
  NOR2X1 U59706 ( .A(n21051), .B(n43224), .Y(n56259) );
  NOR2X1 U59707 ( .A(n44459), .B(n43227), .Y(n56258) );
  NOR2X1 U59708 ( .A(n56259), .B(n56258), .Y(n56261) );
  NOR2X1 U59709 ( .A(n21066), .B(n21065), .Y(n56260) );
  NAND2X1 U59710 ( .A(n56261), .B(n56260), .Y(u_decode_u_regfile_N425) );
  NOR2X1 U59711 ( .A(n19481), .B(n43224), .Y(n56263) );
  NOR2X1 U59712 ( .A(n44549), .B(n43227), .Y(n56262) );
  NOR2X1 U59713 ( .A(n56263), .B(n56262), .Y(n56265) );
  NOR2X1 U59714 ( .A(n19496), .B(n19495), .Y(n56264) );
  NAND2X1 U59715 ( .A(n56265), .B(n56264), .Y(u_decode_u_regfile_N721) );
  NOR2X1 U59716 ( .A(n19088), .B(n43223), .Y(n56267) );
  NOR2X1 U59717 ( .A(n44564), .B(n43226), .Y(n56266) );
  NOR2X1 U59718 ( .A(n56267), .B(n56266), .Y(n56269) );
  NOR2X1 U59719 ( .A(n19102), .B(n19101), .Y(n56268) );
  NAND2X1 U59720 ( .A(n56269), .B(n56268), .Y(u_decode_u_regfile_N795) );
  NOR2X1 U59721 ( .A(n23541), .B(n43223), .Y(n56271) );
  NOR2X1 U59722 ( .A(n44315), .B(n43226), .Y(n56270) );
  NOR2X1 U59723 ( .A(n56271), .B(n56270), .Y(n56273) );
  NOR2X1 U59724 ( .A(n23556), .B(n23555), .Y(n56272) );
  NAND2X1 U59725 ( .A(n56273), .B(n56272), .Y(u_decode_u_regfile_N1091) );
  NOR2X1 U59726 ( .A(n22229), .B(n43223), .Y(n56275) );
  NOR2X1 U59727 ( .A(n44393), .B(n43226), .Y(n56274) );
  NOR2X1 U59728 ( .A(n56275), .B(n56274), .Y(n56277) );
  NOR2X1 U59729 ( .A(n22244), .B(n22243), .Y(n56276) );
  NAND2X1 U59730 ( .A(n56277), .B(n56276), .Y(u_decode_u_regfile_N203) );
  NOR2X1 U59731 ( .A(n20659), .B(n43224), .Y(n56279) );
  NOR2X1 U59732 ( .A(n44483), .B(n43226), .Y(n56278) );
  NOR2X1 U59733 ( .A(n56279), .B(n56278), .Y(n56281) );
  NOR2X1 U59734 ( .A(n20674), .B(n20673), .Y(n56280) );
  NAND2X1 U59735 ( .A(n56281), .B(n56280), .Y(u_decode_u_regfile_N499) );
  NOR2X1 U59736 ( .A(n21837), .B(n43223), .Y(n56283) );
  NOR2X1 U59737 ( .A(n44417), .B(n43226), .Y(n56282) );
  NOR2X1 U59738 ( .A(n56283), .B(n56282), .Y(n56285) );
  NOR2X1 U59739 ( .A(n21852), .B(n21851), .Y(n56284) );
  NAND2X1 U59740 ( .A(n56285), .B(n56284), .Y(u_decode_u_regfile_N277) );
  NOR2X1 U59741 ( .A(n23107), .B(n43223), .Y(n56287) );
  NOR2X1 U59742 ( .A(n44339), .B(n43226), .Y(n56286) );
  NOR2X1 U59743 ( .A(n56287), .B(n56286), .Y(n56289) );
  NOR2X1 U59744 ( .A(n23122), .B(n23121), .Y(n56288) );
  NAND2X1 U59745 ( .A(n56289), .B(n56288), .Y(u_decode_u_regfile_N1165) );
  NOR2X1 U59746 ( .A(n20267), .B(n43223), .Y(n56291) );
  NOR2X1 U59747 ( .A(n44501), .B(n43226), .Y(n56290) );
  NOR2X1 U59748 ( .A(n56291), .B(n56290), .Y(n56293) );
  NOR2X1 U59749 ( .A(n20282), .B(n20281), .Y(n56292) );
  NAND2X1 U59750 ( .A(n56293), .B(n56292), .Y(u_decode_u_regfile_N573) );
  NOR2X1 U59751 ( .A(n18696), .B(n43223), .Y(n56295) );
  NOR2X1 U59752 ( .A(n44576), .B(n43226), .Y(n56294) );
  NOR2X1 U59753 ( .A(n56295), .B(n56294), .Y(n56297) );
  NOR2X1 U59754 ( .A(n18710), .B(n18709), .Y(n56296) );
  NAND2X1 U59755 ( .A(n56297), .B(n56296), .Y(u_decode_u_regfile_N869) );
  NOR2X1 U59756 ( .A(n19875), .B(n43223), .Y(n56299) );
  NOR2X1 U59757 ( .A(n44525), .B(n43226), .Y(n56298) );
  NOR2X1 U59758 ( .A(n56299), .B(n56298), .Y(n56301) );
  NOR2X1 U59759 ( .A(n19890), .B(n19889), .Y(n56300) );
  NAND2X1 U59760 ( .A(n56301), .B(n56300), .Y(u_decode_u_regfile_N647) );
  NOR2X1 U59761 ( .A(n18305), .B(n43223), .Y(n56303) );
  NOR2X1 U59762 ( .A(n44591), .B(n43227), .Y(n56302) );
  NOR2X1 U59763 ( .A(n56303), .B(n56302), .Y(n56305) );
  NOR2X1 U59764 ( .A(n18320), .B(n18319), .Y(n56304) );
  NAND2X1 U59765 ( .A(n56305), .B(n56304), .Y(u_decode_u_regfile_N943) );
  NOR2X1 U59766 ( .A(n22667), .B(n43223), .Y(n56307) );
  NOR2X1 U59767 ( .A(n44363), .B(n43226), .Y(n56306) );
  NOR2X1 U59768 ( .A(n56307), .B(n56306), .Y(n56309) );
  NOR2X1 U59769 ( .A(n22688), .B(n22687), .Y(n56308) );
  NAND2X1 U59770 ( .A(n56309), .B(n56308), .Y(u_decode_u_regfile_N1239) );
  NOR2X1 U59771 ( .A(n21445), .B(n43224), .Y(n56311) );
  NOR2X1 U59772 ( .A(n44441), .B(n43227), .Y(n56310) );
  NOR2X1 U59773 ( .A(n56311), .B(n56310), .Y(n56313) );
  NOR2X1 U59774 ( .A(n21460), .B(n21459), .Y(n56312) );
  NAND2X1 U59775 ( .A(n56313), .B(n56312), .Y(u_decode_u_regfile_N351) );
  MX2X1 U59776 ( .A(u_csr_pc_m_q[29]), .B(opcode_pc_w[29]), .S0(n58128), .Y(
        n8500) );
  NAND2X1 U59777 ( .A(n43288), .B(n56349), .Y(n56315) );
  NAND2X1 U59778 ( .A(n43236), .B(n44024), .Y(n56314) );
  NAND2X1 U59779 ( .A(n56315), .B(n56314), .Y(n56321) );
  INVX1 U59780 ( .A(n56316), .Y(n56330) );
  NAND2X1 U59781 ( .A(n56330), .B(n43239), .Y(n56319) );
  NAND2X1 U59782 ( .A(n44282), .B(n44029), .Y(n56331) );
  NAND2X1 U59783 ( .A(n27477), .B(n56331), .Y(n56317) );
  NAND2X1 U59784 ( .A(u_csr_csr_mepc_q[29]), .B(n56317), .Y(n56318) );
  NAND2X1 U59785 ( .A(n56319), .B(n56318), .Y(n56320) );
  NOR2X1 U59786 ( .A(n56321), .B(n56320), .Y(n56327) );
  NOR2X1 U59787 ( .A(n42952), .B(n37759), .Y(n56325) );
  NAND2X1 U59788 ( .A(n43243), .B(opcode_pc_w[29]), .Y(n56323) );
  NAND2X1 U59789 ( .A(n43248), .B(n56348), .Y(n56322) );
  NAND2X1 U59790 ( .A(n56323), .B(n56322), .Y(n56324) );
  NOR2X1 U59791 ( .A(n56325), .B(n56324), .Y(n56326) );
  NAND2X1 U59792 ( .A(n56327), .B(n56326), .Y(u_csr_csr_mepc_r[29]) );
  NAND2X1 U59793 ( .A(n43291), .B(n56348), .Y(n56329) );
  NAND2X1 U59794 ( .A(n43253), .B(n44027), .Y(n56328) );
  NAND2X1 U59795 ( .A(n56329), .B(n56328), .Y(n56336) );
  NAND2X1 U59796 ( .A(n56330), .B(n43249), .Y(n56334) );
  NAND2X1 U59797 ( .A(n26373), .B(n56331), .Y(n56332) );
  NAND2X1 U59798 ( .A(u_csr_csr_sepc_q[29]), .B(n56332), .Y(n56333) );
  NAND2X1 U59799 ( .A(n56334), .B(n56333), .Y(n56335) );
  NOR2X1 U59800 ( .A(n56336), .B(n56335), .Y(n56342) );
  NOR2X1 U59801 ( .A(n42955), .B(n37759), .Y(n56340) );
  NAND2X1 U59802 ( .A(n43256), .B(opcode_pc_w[29]), .Y(n56338) );
  NAND2X1 U59803 ( .A(n56600), .B(n56349), .Y(n56337) );
  NAND2X1 U59804 ( .A(n56338), .B(n56337), .Y(n56339) );
  NOR2X1 U59805 ( .A(n56340), .B(n56339), .Y(n56341) );
  NAND2X1 U59806 ( .A(n56342), .B(n56341), .Y(u_csr_csr_sepc_r[29]) );
  AND2X1 U59807 ( .A(n28278), .B(n28276), .Y(n56347) );
  NOR2X1 U59808 ( .A(n56343), .B(n43292), .Y(n56345) );
  NOR2X1 U59809 ( .A(n58486), .B(n43295), .Y(n56344) );
  NOR2X1 U59810 ( .A(n56345), .B(n56344), .Y(n56346) );
  NAND2X1 U59811 ( .A(n56347), .B(n56346), .Y(u_csr_N3694) );
  NAND2X1 U59812 ( .A(n43300), .B(n56348), .Y(n56351) );
  NAND2X1 U59813 ( .A(n43303), .B(n56349), .Y(n56350) );
  NAND2X1 U59814 ( .A(n56351), .B(n56350), .Y(net2315) );
  XNOR2X1 U59815 ( .A(n56352), .B(n42414), .Y(u_fetch_N78) );
  NAND2X1 U59816 ( .A(n44833), .B(n44019), .Y(n56362) );
  NAND2X1 U59817 ( .A(n44021), .B(n44845), .Y(n56360) );
  NAND2X1 U59818 ( .A(n44833), .B(n44010), .Y(n56359) );
  NAND2X1 U59819 ( .A(n44013), .B(n44845), .Y(n56357) );
  NAND2X1 U59820 ( .A(n44833), .B(n44002), .Y(n56356) );
  NAND2X1 U59821 ( .A(n44004), .B(n44845), .Y(n56354) );
  NAND2X1 U59822 ( .A(n56354), .B(n56353), .Y(n56355) );
  NAND2X1 U59823 ( .A(n56356), .B(n56355), .Y(n56631) );
  NAND2X1 U59824 ( .A(n56357), .B(n56631), .Y(n56358) );
  NAND2X1 U59825 ( .A(n56359), .B(n56358), .Y(n56703) );
  NAND2X1 U59826 ( .A(n56360), .B(n56703), .Y(n56361) );
  NAND2X1 U59827 ( .A(n56362), .B(n56361), .Y(n56545) );
  INVX1 U59828 ( .A(n56545), .Y(n56364) );
  XNOR2X1 U59829 ( .A(n44837), .B(n56364), .Y(n56363) );
  NAND2X1 U59830 ( .A(n56363), .B(n43375), .Y(n56366) );
  MX2X1 U59831 ( .A(n37555), .B(n42219), .S0(n56364), .Y(n56365) );
  MX2X1 U59832 ( .A(n56366), .B(n56365), .S0(n44029), .Y(u_lsu_mem_addr_r[29])
         );
  NAND2X1 U59833 ( .A(n42253), .B(n56367), .Y(n56369) );
  NAND2X1 U59834 ( .A(n42252), .B(n14), .Y(n56368) );
  NAND2X1 U59835 ( .A(u_mmu_virt_addr_q_29), .B(n57397), .Y(n56370) );
  NAND2X1 U59836 ( .A(n42422), .B(n56370), .Y(n8552) );
  MX2X1 U59837 ( .A(u_mmu_itlb_va_addr_q[29]), .B(u_mmu_virt_addr_q_29), .S0(
        n37548), .Y(n8444) );
  NOR2X1 U59838 ( .A(n43315), .B(n56374), .Y(net2415) );
  INVX1 U59839 ( .A(n56566), .Y(n56371) );
  XNOR2X1 U59840 ( .A(opcode_pc_w[30]), .B(n56371), .Y(n56509) );
  NOR2X1 U59841 ( .A(n43326), .B(n56509), .Y(n56373) );
  NOR2X1 U59842 ( .A(n56373), .B(n56372), .Y(n56378) );
  NOR2X1 U59843 ( .A(n1929), .B(n43322), .Y(n56376) );
  NOR2X1 U59844 ( .A(n43325), .B(n56374), .Y(n56375) );
  NOR2X1 U59845 ( .A(n56376), .B(n56375), .Y(n56377) );
  NAND2X1 U59846 ( .A(n56378), .B(n56377), .Y(u_decode_N320) );
  NAND2X1 U59847 ( .A(n15836), .B(n42451), .Y(n56379) );
  NAND2X1 U59848 ( .A(n15834), .B(n56379), .Y(n56380) );
  NOR2X1 U59849 ( .A(n15881), .B(n56380), .Y(n56382) );
  NOR2X1 U59850 ( .A(n15832), .B(n15882), .Y(n56381) );
  NAND2X1 U59851 ( .A(n56382), .B(n56381), .Y(u_exec_alu_p_w[30]) );
  NOR2X1 U59852 ( .A(n44539), .B(n43231), .Y(n56384) );
  NOR2X1 U59853 ( .A(n44537), .B(n43234), .Y(n56383) );
  NOR2X1 U59854 ( .A(n56384), .B(n56383), .Y(n56386) );
  NOR2X1 U59855 ( .A(n19687), .B(n19686), .Y(n56385) );
  NAND2X1 U59856 ( .A(n56386), .B(n56385), .Y(u_decode_u_regfile_N685) );
  NOR2X1 U59857 ( .A(n44603), .B(n43231), .Y(n56388) );
  NOR2X1 U59858 ( .A(n44600), .B(n43234), .Y(n56387) );
  NOR2X1 U59859 ( .A(n56388), .B(n56387), .Y(n56390) );
  NOR2X1 U59860 ( .A(n18097), .B(n18095), .Y(n56389) );
  NAND2X1 U59861 ( .A(n56390), .B(n56389), .Y(u_decode_u_regfile_N981) );
  NOR2X1 U59862 ( .A(n43229), .B(n57131), .Y(n56392) );
  NOR2X1 U59863 ( .A(n43232), .B(n43386), .Y(n56391) );
  NOR2X1 U59864 ( .A(n56392), .B(n56391), .Y(n56394) );
  NOR2X1 U59865 ( .A(n21257), .B(n21256), .Y(n56393) );
  NAND2X1 U59866 ( .A(n56394), .B(n56393), .Y(u_decode_u_regfile_N389) );
  NOR2X1 U59867 ( .A(n44474), .B(n43231), .Y(n56396) );
  NOR2X1 U59868 ( .A(n44471), .B(n43234), .Y(n56395) );
  NOR2X1 U59869 ( .A(n56396), .B(n56395), .Y(n56398) );
  NOR2X1 U59870 ( .A(n20864), .B(n20863), .Y(n56397) );
  NAND2X1 U59871 ( .A(n56398), .B(n56397), .Y(u_decode_u_regfile_N463) );
  NOR2X1 U59872 ( .A(n44561), .B(n43231), .Y(n56400) );
  NOR2X1 U59873 ( .A(n44558), .B(n43234), .Y(n56399) );
  NOR2X1 U59874 ( .A(n56400), .B(n56399), .Y(n56402) );
  NOR2X1 U59875 ( .A(n19292), .B(n19291), .Y(n56401) );
  NAND2X1 U59876 ( .A(n56402), .B(n56401), .Y(u_decode_u_regfile_N759) );
  NOR2X1 U59877 ( .A(n22425), .B(n43230), .Y(n56404) );
  NOR2X1 U59878 ( .A(n44381), .B(n43234), .Y(n56403) );
  NOR2X1 U59879 ( .A(n56404), .B(n56403), .Y(n56406) );
  NOR2X1 U59880 ( .A(n22434), .B(n22433), .Y(n56405) );
  NAND2X1 U59881 ( .A(n56406), .B(n56405), .Y(u_decode_u_regfile_N167) );
  NOR2X1 U59882 ( .A(n23761), .B(n43230), .Y(n56408) );
  NOR2X1 U59883 ( .A(n44303), .B(n43233), .Y(n56407) );
  NOR2X1 U59884 ( .A(n56408), .B(n56407), .Y(n56410) );
  NOR2X1 U59885 ( .A(n23770), .B(n23769), .Y(n56409) );
  NAND2X1 U59886 ( .A(n56410), .B(n56409), .Y(u_decode_u_regfile_N1055) );
  NOR2X1 U59887 ( .A(n44573), .B(n43230), .Y(n56412) );
  NOR2X1 U59888 ( .A(n44570), .B(n43233), .Y(n56411) );
  NOR2X1 U59889 ( .A(n56412), .B(n56411), .Y(n56414) );
  NOR2X1 U59890 ( .A(n18900), .B(n18899), .Y(n56413) );
  NAND2X1 U59891 ( .A(n56414), .B(n56413), .Y(u_decode_u_regfile_N833) );
  NOR2X1 U59892 ( .A(n43229), .B(n57209), .Y(n56416) );
  NOR2X1 U59893 ( .A(n43232), .B(n43383), .Y(n56415) );
  NOR2X1 U59894 ( .A(n56416), .B(n56415), .Y(n56418) );
  NOR2X1 U59895 ( .A(n20472), .B(n20471), .Y(n56417) );
  NAND2X1 U59896 ( .A(n56418), .B(n56417), .Y(u_decode_u_regfile_N537) );
  NOR2X1 U59897 ( .A(n22033), .B(n43230), .Y(n56420) );
  NOR2X1 U59898 ( .A(n44405), .B(n43233), .Y(n56419) );
  NOR2X1 U59899 ( .A(n56420), .B(n56419), .Y(n56422) );
  NOR2X1 U59900 ( .A(n22042), .B(n22041), .Y(n56421) );
  NAND2X1 U59901 ( .A(n56422), .B(n56421), .Y(u_decode_u_regfile_N241) );
  NOR2X1 U59902 ( .A(n23321), .B(n43230), .Y(n56424) );
  NOR2X1 U59903 ( .A(n44327), .B(n43233), .Y(n56423) );
  NOR2X1 U59904 ( .A(n56424), .B(n56423), .Y(n56426) );
  NOR2X1 U59905 ( .A(n23336), .B(n23335), .Y(n56425) );
  NAND2X1 U59906 ( .A(n56426), .B(n56425), .Y(u_decode_u_regfile_N1129) );
  NOR2X1 U59907 ( .A(n44585), .B(n43230), .Y(n56428) );
  NOR2X1 U59908 ( .A(n44582), .B(n43233), .Y(n56427) );
  NOR2X1 U59909 ( .A(n56428), .B(n56427), .Y(n56430) );
  NOR2X1 U59910 ( .A(n18508), .B(n18507), .Y(n56429) );
  NAND2X1 U59911 ( .A(n56430), .B(n56429), .Y(u_decode_u_regfile_N907) );
  NOR2X1 U59912 ( .A(n21641), .B(n43230), .Y(n56432) );
  NOR2X1 U59913 ( .A(n44429), .B(n43233), .Y(n56431) );
  NOR2X1 U59914 ( .A(n56432), .B(n56431), .Y(n56434) );
  NOR2X1 U59915 ( .A(n21650), .B(n21649), .Y(n56433) );
  NAND2X1 U59916 ( .A(n56434), .B(n56433), .Y(u_decode_u_regfile_N315) );
  NOR2X1 U59917 ( .A(n20071), .B(n43230), .Y(n56436) );
  NOR2X1 U59918 ( .A(n44513), .B(n43233), .Y(n56435) );
  NOR2X1 U59919 ( .A(n56436), .B(n56435), .Y(n56438) );
  NOR2X1 U59920 ( .A(n20080), .B(n20079), .Y(n56437) );
  NAND2X1 U59921 ( .A(n56438), .B(n56437), .Y(u_decode_u_regfile_N611) );
  NOR2X1 U59922 ( .A(n22887), .B(n43230), .Y(n56440) );
  NOR2X1 U59923 ( .A(n44351), .B(n43233), .Y(n56439) );
  NOR2X1 U59924 ( .A(n56440), .B(n56439), .Y(n56442) );
  NOR2X1 U59925 ( .A(n22896), .B(n22895), .Y(n56441) );
  NAND2X1 U59926 ( .A(n56442), .B(n56441), .Y(u_decode_u_regfile_N1203) );
  NOR2X1 U59927 ( .A(n18002), .B(n43230), .Y(n56444) );
  NOR2X1 U59928 ( .A(n44606), .B(n43233), .Y(n56443) );
  NOR2X1 U59929 ( .A(n56444), .B(n56443), .Y(n56446) );
  NOR2X1 U59930 ( .A(n23986), .B(n23985), .Y(n56445) );
  NAND2X1 U59931 ( .A(n56446), .B(n56445), .Y(u_decode_u_regfile_N1018) );
  NOR2X1 U59932 ( .A(n43229), .B(n57144), .Y(n56448) );
  NOR2X1 U59933 ( .A(n43232), .B(n43389), .Y(n56447) );
  NOR2X1 U59934 ( .A(n56448), .B(n56447), .Y(n56450) );
  NOR2X1 U59935 ( .A(n22630), .B(n22629), .Y(n56449) );
  NAND2X1 U59936 ( .A(n56450), .B(n56449), .Y(u_decode_u_regfile_N130) );
  NOR2X1 U59937 ( .A(n21051), .B(n43230), .Y(n56452) );
  NOR2X1 U59938 ( .A(n44459), .B(n43233), .Y(n56451) );
  NOR2X1 U59939 ( .A(n56452), .B(n56451), .Y(n56454) );
  NOR2X1 U59940 ( .A(n21060), .B(n21059), .Y(n56453) );
  NAND2X1 U59941 ( .A(n56454), .B(n56453), .Y(u_decode_u_regfile_N426) );
  NOR2X1 U59942 ( .A(n19481), .B(n43230), .Y(n56456) );
  NOR2X1 U59943 ( .A(n44549), .B(n43233), .Y(n56455) );
  NOR2X1 U59944 ( .A(n56456), .B(n56455), .Y(n56458) );
  NOR2X1 U59945 ( .A(n19490), .B(n19489), .Y(n56457) );
  NAND2X1 U59946 ( .A(n56458), .B(n56457), .Y(u_decode_u_regfile_N722) );
  NOR2X1 U59947 ( .A(n19088), .B(n43229), .Y(n56460) );
  NOR2X1 U59948 ( .A(n44564), .B(n43233), .Y(n56459) );
  NOR2X1 U59949 ( .A(n56460), .B(n56459), .Y(n56462) );
  NOR2X1 U59950 ( .A(n19096), .B(n19095), .Y(n56461) );
  NAND2X1 U59951 ( .A(n56462), .B(n56461), .Y(u_decode_u_regfile_N796) );
  NOR2X1 U59952 ( .A(n23541), .B(n43229), .Y(n56464) );
  NOR2X1 U59953 ( .A(n44315), .B(n43232), .Y(n56463) );
  NOR2X1 U59954 ( .A(n56464), .B(n56463), .Y(n56466) );
  NOR2X1 U59955 ( .A(n23550), .B(n23549), .Y(n56465) );
  NAND2X1 U59956 ( .A(n56466), .B(n56465), .Y(u_decode_u_regfile_N1092) );
  NOR2X1 U59957 ( .A(n22229), .B(n43229), .Y(n56468) );
  NOR2X1 U59958 ( .A(n44393), .B(n43232), .Y(n56467) );
  NOR2X1 U59959 ( .A(n56468), .B(n56467), .Y(n56470) );
  NOR2X1 U59960 ( .A(n22238), .B(n22237), .Y(n56469) );
  NAND2X1 U59961 ( .A(n56470), .B(n56469), .Y(u_decode_u_regfile_N204) );
  NOR2X1 U59962 ( .A(n20659), .B(n43229), .Y(n56472) );
  NOR2X1 U59963 ( .A(n44483), .B(n43232), .Y(n56471) );
  NOR2X1 U59964 ( .A(n56472), .B(n56471), .Y(n56474) );
  NOR2X1 U59965 ( .A(n20668), .B(n20667), .Y(n56473) );
  NAND2X1 U59966 ( .A(n56474), .B(n56473), .Y(u_decode_u_regfile_N500) );
  NOR2X1 U59967 ( .A(n21837), .B(n43229), .Y(n56476) );
  NOR2X1 U59968 ( .A(n44417), .B(n43232), .Y(n56475) );
  NOR2X1 U59969 ( .A(n56476), .B(n56475), .Y(n56478) );
  NOR2X1 U59970 ( .A(n21846), .B(n21845), .Y(n56477) );
  NAND2X1 U59971 ( .A(n56478), .B(n56477), .Y(u_decode_u_regfile_N278) );
  NOR2X1 U59972 ( .A(n23107), .B(n43229), .Y(n56480) );
  NOR2X1 U59973 ( .A(n44339), .B(n43232), .Y(n56479) );
  NOR2X1 U59974 ( .A(n56480), .B(n56479), .Y(n56482) );
  NOR2X1 U59975 ( .A(n23116), .B(n23115), .Y(n56481) );
  NAND2X1 U59976 ( .A(n56482), .B(n56481), .Y(u_decode_u_regfile_N1166) );
  NOR2X1 U59977 ( .A(n20267), .B(n43229), .Y(n56484) );
  NOR2X1 U59978 ( .A(n44501), .B(n43232), .Y(n56483) );
  NOR2X1 U59979 ( .A(n56484), .B(n56483), .Y(n56486) );
  NOR2X1 U59980 ( .A(n20276), .B(n20275), .Y(n56485) );
  NAND2X1 U59981 ( .A(n56486), .B(n56485), .Y(u_decode_u_regfile_N574) );
  NOR2X1 U59982 ( .A(n18696), .B(n43229), .Y(n56488) );
  NOR2X1 U59983 ( .A(n44576), .B(n43232), .Y(n56487) );
  NOR2X1 U59984 ( .A(n56488), .B(n56487), .Y(n56490) );
  NOR2X1 U59985 ( .A(n18704), .B(n18703), .Y(n56489) );
  NAND2X1 U59986 ( .A(n56490), .B(n56489), .Y(u_decode_u_regfile_N870) );
  NOR2X1 U59987 ( .A(n19875), .B(n43229), .Y(n56492) );
  NOR2X1 U59988 ( .A(n44525), .B(n43232), .Y(n56491) );
  NOR2X1 U59989 ( .A(n56492), .B(n56491), .Y(n56494) );
  NOR2X1 U59990 ( .A(n19884), .B(n19883), .Y(n56493) );
  NAND2X1 U59991 ( .A(n56494), .B(n56493), .Y(u_decode_u_regfile_N648) );
  NOR2X1 U59992 ( .A(n18305), .B(n43230), .Y(n56496) );
  NOR2X1 U59993 ( .A(n44591), .B(n43233), .Y(n56495) );
  NOR2X1 U59994 ( .A(n56496), .B(n56495), .Y(n56498) );
  NOR2X1 U59995 ( .A(n18314), .B(n18313), .Y(n56497) );
  NAND2X1 U59996 ( .A(n56498), .B(n56497), .Y(u_decode_u_regfile_N944) );
  NOR2X1 U59997 ( .A(n22667), .B(n43229), .Y(n56500) );
  NOR2X1 U59998 ( .A(n44363), .B(n43232), .Y(n56499) );
  NOR2X1 U59999 ( .A(n56500), .B(n56499), .Y(n56502) );
  NOR2X1 U60000 ( .A(n22676), .B(n22675), .Y(n56501) );
  NAND2X1 U60001 ( .A(n56502), .B(n56501), .Y(u_decode_u_regfile_N1240) );
  NOR2X1 U60002 ( .A(n21445), .B(n43230), .Y(n56504) );
  NOR2X1 U60003 ( .A(n44441), .B(n43233), .Y(n56503) );
  NOR2X1 U60004 ( .A(n56504), .B(n56503), .Y(n56506) );
  NOR2X1 U60005 ( .A(n21454), .B(n21453), .Y(n56505) );
  NAND2X1 U60006 ( .A(n56506), .B(n56505), .Y(u_decode_u_regfile_N352) );
  MX2X1 U60007 ( .A(u_csr_pc_m_q[30]), .B(opcode_pc_w[30]), .S0(n58128), .Y(
        n8499) );
  NAND2X1 U60008 ( .A(n43288), .B(n56542), .Y(n56508) );
  NAND2X1 U60009 ( .A(n43236), .B(n44050), .Y(n56507) );
  NAND2X1 U60010 ( .A(n56508), .B(n56507), .Y(n56514) );
  INVX1 U60011 ( .A(n56509), .Y(n56523) );
  NAND2X1 U60012 ( .A(n56523), .B(n43239), .Y(n56512) );
  NAND2X1 U60013 ( .A(n44282), .B(n44053), .Y(n56524) );
  NAND2X1 U60014 ( .A(n27477), .B(n56524), .Y(n56510) );
  NAND2X1 U60015 ( .A(u_csr_csr_mepc_q[30]), .B(n56510), .Y(n56511) );
  NAND2X1 U60016 ( .A(n56512), .B(n56511), .Y(n56513) );
  NOR2X1 U60017 ( .A(n56514), .B(n56513), .Y(n56520) );
  NOR2X1 U60018 ( .A(n42953), .B(n37760), .Y(n56518) );
  NAND2X1 U60019 ( .A(n43243), .B(opcode_pc_w[30]), .Y(n56516) );
  NAND2X1 U60020 ( .A(n43248), .B(n56541), .Y(n56515) );
  NAND2X1 U60021 ( .A(n56516), .B(n56515), .Y(n56517) );
  NOR2X1 U60022 ( .A(n56518), .B(n56517), .Y(n56519) );
  NAND2X1 U60023 ( .A(n56520), .B(n56519), .Y(u_csr_csr_mepc_r[30]) );
  NAND2X1 U60024 ( .A(n43291), .B(n56541), .Y(n56522) );
  NAND2X1 U60025 ( .A(n43253), .B(n44050), .Y(n56521) );
  NAND2X1 U60026 ( .A(n56522), .B(n56521), .Y(n56529) );
  NAND2X1 U60027 ( .A(n56523), .B(n43249), .Y(n56527) );
  NAND2X1 U60028 ( .A(n26373), .B(n56524), .Y(n56525) );
  NAND2X1 U60029 ( .A(u_csr_csr_sepc_q[30]), .B(n56525), .Y(n56526) );
  NAND2X1 U60030 ( .A(n56527), .B(n56526), .Y(n56528) );
  NOR2X1 U60031 ( .A(n56529), .B(n56528), .Y(n56535) );
  NOR2X1 U60032 ( .A(n42956), .B(n37760), .Y(n56533) );
  NAND2X1 U60033 ( .A(n43256), .B(opcode_pc_w[30]), .Y(n56531) );
  NAND2X1 U60034 ( .A(n56600), .B(n56542), .Y(n56530) );
  NAND2X1 U60035 ( .A(n56531), .B(n56530), .Y(n56532) );
  NOR2X1 U60036 ( .A(n56533), .B(n56532), .Y(n56534) );
  NAND2X1 U60037 ( .A(n56535), .B(n56534), .Y(u_csr_csr_sepc_r[30]) );
  AND2X1 U60038 ( .A(n28270), .B(n28268), .Y(n56540) );
  NOR2X1 U60039 ( .A(n58489), .B(n43292), .Y(n56538) );
  NOR2X1 U60040 ( .A(n56536), .B(n43295), .Y(n56537) );
  NOR2X1 U60041 ( .A(n56538), .B(n56537), .Y(n56539) );
  NAND2X1 U60042 ( .A(n56540), .B(n56539), .Y(u_csr_N3695) );
  NAND2X1 U60043 ( .A(n43300), .B(n56541), .Y(n56544) );
  NAND2X1 U60044 ( .A(n43303), .B(n56542), .Y(n56543) );
  NAND2X1 U60045 ( .A(n56544), .B(n56543), .Y(net2316) );
  INVX1 U60046 ( .A(n16), .Y(n56617) );
  NAND2X1 U60047 ( .A(n42414), .B(n14), .Y(n56616) );
  NAND2X1 U60048 ( .A(n44833), .B(n44027), .Y(n56548) );
  NAND2X1 U60049 ( .A(n44028), .B(n44843), .Y(n56546) );
  NAND2X1 U60050 ( .A(n56546), .B(n56545), .Y(n56547) );
  NAND2X1 U60051 ( .A(n56548), .B(n56547), .Y(n56620) );
  INVX1 U60052 ( .A(n56620), .Y(n56550) );
  XNOR2X1 U60053 ( .A(n42852), .B(n56550), .Y(n56549) );
  NAND2X1 U60054 ( .A(n56549), .B(n43375), .Y(n56552) );
  MX2X1 U60055 ( .A(n37555), .B(n42219), .S0(n56550), .Y(n56551) );
  MX2X1 U60056 ( .A(n56552), .B(n56551), .S0(n44053), .Y(u_lsu_mem_addr_r[30])
         );
  NAND2X1 U60057 ( .A(n42253), .B(n56553), .Y(n56555) );
  NAND2X1 U60058 ( .A(n42252), .B(n16), .Y(n56554) );
  NAND2X1 U60059 ( .A(u_mmu_virt_addr_q_30), .B(n57397), .Y(n56556) );
  NAND2X1 U60060 ( .A(n42421), .B(n56556), .Y(n8553) );
  MX2X1 U60061 ( .A(u_mmu_itlb_va_addr_q[30]), .B(u_mmu_virt_addr_q_30), .S0(
        n37548), .Y(n8427) );
  INVX1 U60062 ( .A(n56557), .Y(n56559) );
  XNOR2X1 U60063 ( .A(n44837), .B(n56559), .Y(n56558) );
  NAND2X1 U60064 ( .A(n56558), .B(n43375), .Y(n56561) );
  MX2X1 U60065 ( .A(n37555), .B(n42219), .S0(n56559), .Y(n56560) );
  MX2X1 U60066 ( .A(n56561), .B(n56560), .S0(n43949), .Y(u_lsu_mem_addr_r[22])
         );
  NOR2X1 U60067 ( .A(n2483), .B(n40673), .Y(n56563) );
  NOR2X1 U60068 ( .A(n8318), .B(n40688), .Y(n56562) );
  NOR2X1 U60069 ( .A(n56563), .B(n56562), .Y(n56565) );
  NAND2X1 U60070 ( .A(n56767), .B(n17), .Y(n56564) );
  NAND2X1 U60071 ( .A(n56565), .B(n56564), .Y(u_mmu_request_addr_w[22]) );
  MX2X1 U60072 ( .A(u_mmu_itlb_va_addr_q[22]), .B(n57388), .S0(n37548), .Y(
        n8436) );
  NOR2X1 U60073 ( .A(n43315), .B(n56570), .Y(net2416) );
  NOR2X1 U60074 ( .A(n58409), .B(n56566), .Y(n56567) );
  XNOR2X1 U60075 ( .A(opcode_pc_w[31]), .B(n56567), .Y(n56577) );
  NOR2X1 U60076 ( .A(n43326), .B(n56577), .Y(n56569) );
  NOR2X1 U60077 ( .A(n56569), .B(n56568), .Y(n56574) );
  NOR2X1 U60078 ( .A(n1930), .B(n43322), .Y(n56572) );
  NOR2X1 U60079 ( .A(n43325), .B(n56570), .Y(n56571) );
  NOR2X1 U60080 ( .A(n56572), .B(n56571), .Y(n56573) );
  NAND2X1 U60081 ( .A(n56574), .B(n56573), .Y(u_decode_N321) );
  MX2X1 U60082 ( .A(u_csr_pc_m_q[31]), .B(opcode_pc_w[31]), .S0(n58128), .Y(
        n8537) );
  NAND2X1 U60083 ( .A(n43288), .B(n56613), .Y(n56576) );
  NAND2X1 U60084 ( .A(n43236), .B(n44057), .Y(n56575) );
  NAND2X1 U60085 ( .A(n56576), .B(n56575), .Y(n56583) );
  INVX1 U60086 ( .A(n56577), .Y(n56591) );
  NAND2X1 U60087 ( .A(n56591), .B(n43239), .Y(n56581) );
  NAND2X1 U60088 ( .A(n44282), .B(n44060), .Y(n56594) );
  NAND2X1 U60089 ( .A(n27477), .B(n56594), .Y(n56579) );
  NAND2X1 U60090 ( .A(u_csr_csr_mepc_q[31]), .B(n56579), .Y(n56580) );
  NAND2X1 U60091 ( .A(n56581), .B(n56580), .Y(n56582) );
  NOR2X1 U60092 ( .A(n56583), .B(n56582), .Y(n56589) );
  NOR2X1 U60093 ( .A(n42952), .B(n37761), .Y(n56587) );
  NAND2X1 U60094 ( .A(n43243), .B(opcode_pc_w[31]), .Y(n56585) );
  NAND2X1 U60095 ( .A(n43248), .B(n56612), .Y(n56584) );
  NAND2X1 U60096 ( .A(n56585), .B(n56584), .Y(n56586) );
  NOR2X1 U60097 ( .A(n56587), .B(n56586), .Y(n56588) );
  NAND2X1 U60098 ( .A(n56589), .B(n56588), .Y(u_csr_csr_mepc_r[31]) );
  NAND2X1 U60099 ( .A(n56591), .B(n43249), .Y(n56593) );
  NAND2X1 U60100 ( .A(n43291), .B(n56612), .Y(n56592) );
  NAND2X1 U60101 ( .A(n56593), .B(n56592), .Y(n56599) );
  NAND2X1 U60102 ( .A(n43253), .B(n44057), .Y(n56597) );
  NAND2X1 U60103 ( .A(n26373), .B(n56594), .Y(n56595) );
  NAND2X1 U60104 ( .A(u_csr_csr_sepc_q[31]), .B(n56595), .Y(n56596) );
  NAND2X1 U60105 ( .A(n56597), .B(n56596), .Y(n56598) );
  NOR2X1 U60106 ( .A(n56599), .B(n56598), .Y(n56606) );
  NOR2X1 U60107 ( .A(n42956), .B(n37761), .Y(n56604) );
  NAND2X1 U60108 ( .A(n43256), .B(opcode_pc_w[31]), .Y(n56602) );
  NAND2X1 U60109 ( .A(n56600), .B(n56613), .Y(n56601) );
  NAND2X1 U60110 ( .A(n56602), .B(n56601), .Y(n56603) );
  NOR2X1 U60111 ( .A(n56604), .B(n56603), .Y(n56605) );
  NAND2X1 U60112 ( .A(n56606), .B(n56605), .Y(u_csr_csr_sepc_r[31]) );
  AND2X1 U60113 ( .A(n28259), .B(n28256), .Y(n56611) );
  NOR2X1 U60114 ( .A(n58490), .B(n43292), .Y(n56609) );
  NOR2X1 U60115 ( .A(n56607), .B(n43295), .Y(n56608) );
  NOR2X1 U60116 ( .A(n56609), .B(n56608), .Y(n56610) );
  NAND2X1 U60117 ( .A(n56611), .B(n56610), .Y(u_csr_N3696) );
  NAND2X1 U60118 ( .A(n43300), .B(n56612), .Y(n56615) );
  NAND2X1 U60119 ( .A(n43303), .B(n56613), .Y(n56614) );
  NAND2X1 U60120 ( .A(n56615), .B(n56614), .Y(net2317) );
  XNOR2X1 U60121 ( .A(n56619), .B(n56618), .Y(u_fetch_N80) );
  NAND2X1 U60122 ( .A(n44833), .B(n44050), .Y(n56623) );
  NAND2X1 U60123 ( .A(n44051), .B(n44843), .Y(n56621) );
  NAND2X1 U60124 ( .A(n56621), .B(n56620), .Y(n56622) );
  XNOR2X1 U60125 ( .A(n42852), .B(n42123), .Y(n56624) );
  NAND2X1 U60126 ( .A(n56624), .B(n43375), .Y(n56626) );
  MX2X1 U60127 ( .A(n37555), .B(n42219), .S0(n42123), .Y(n56625) );
  MX2X1 U60128 ( .A(n56626), .B(n56625), .S0(n44060), .Y(u_lsu_mem_addr_r[31])
         );
  NAND2X1 U60129 ( .A(n42253), .B(n56627), .Y(n56629) );
  NAND2X1 U60130 ( .A(n42252), .B(\mmu_ifetch_pc_w[31] ), .Y(n56628) );
  NAND2X1 U60131 ( .A(u_mmu_virt_addr_q_31), .B(n57397), .Y(n56630) );
  NAND2X1 U60132 ( .A(n42423), .B(n56630), .Y(n8560) );
  MX2X1 U60133 ( .A(u_mmu_itlb_va_addr_q[31]), .B(u_mmu_virt_addr_q_31), .S0(
        n37548), .Y(n8425) );
  INVX1 U60134 ( .A(n56631), .Y(n56633) );
  XNOR2X1 U60135 ( .A(n44837), .B(n56633), .Y(n56632) );
  NAND2X1 U60136 ( .A(n56632), .B(n43375), .Y(n56635) );
  MX2X1 U60137 ( .A(n37555), .B(n42219), .S0(n56633), .Y(n56634) );
  MX2X1 U60138 ( .A(n56635), .B(n56634), .S0(n44013), .Y(u_lsu_mem_addr_r[27])
         );
  NOR2X1 U60139 ( .A(n2785), .B(n40671), .Y(n56637) );
  NOR2X1 U60140 ( .A(n8328), .B(n40686), .Y(n56636) );
  NOR2X1 U60141 ( .A(n56637), .B(n56636), .Y(n56639) );
  NAND2X1 U60142 ( .A(n56767), .B(n19), .Y(n56638) );
  NAND2X1 U60143 ( .A(n56639), .B(n56638), .Y(u_mmu_request_addr_w[27]) );
  MX2X1 U60144 ( .A(u_mmu_itlb_va_addr_q[27]), .B(n57390), .S0(n37548), .Y(
        n8442) );
  INVX1 U60145 ( .A(n56640), .Y(n56642) );
  XNOR2X1 U60146 ( .A(n42852), .B(n56642), .Y(n56641) );
  NAND2X1 U60147 ( .A(n56641), .B(n43375), .Y(n56644) );
  MX2X1 U60148 ( .A(n37555), .B(n42219), .S0(n56642), .Y(n56643) );
  MX2X1 U60149 ( .A(n56644), .B(n56643), .S0(n43996), .Y(u_lsu_mem_addr_r[25])
         );
  NOR2X1 U60150 ( .A(n2817), .B(n40672), .Y(n56646) );
  NOR2X1 U60151 ( .A(n8324), .B(n40687), .Y(n56645) );
  NOR2X1 U60152 ( .A(n56646), .B(n56645), .Y(n56648) );
  NAND2X1 U60153 ( .A(n56767), .B(n23), .Y(n56647) );
  NAND2X1 U60154 ( .A(n56648), .B(n56647), .Y(u_mmu_request_addr_w[25]) );
  MX2X1 U60155 ( .A(u_mmu_itlb_va_addr_q[25]), .B(n57391), .S0(n37548), .Y(
        n8431) );
  INVX1 U60156 ( .A(n56649), .Y(n56651) );
  XNOR2X1 U60157 ( .A(n42852), .B(n56651), .Y(n56650) );
  NAND2X1 U60158 ( .A(n56650), .B(n43375), .Y(n56653) );
  MX2X1 U60159 ( .A(n37555), .B(n42219), .S0(n56651), .Y(n56652) );
  MX2X1 U60160 ( .A(n56653), .B(n56652), .S0(n43908), .Y(u_lsu_mem_addr_r[17])
         );
  NOR2X1 U60161 ( .A(n2882), .B(n40671), .Y(n56655) );
  NOR2X1 U60162 ( .A(n8306), .B(n40686), .Y(n56654) );
  NOR2X1 U60163 ( .A(n56655), .B(n56654), .Y(n56657) );
  NAND2X1 U60164 ( .A(n56767), .B(n6), .Y(n56656) );
  NAND2X1 U60165 ( .A(n56657), .B(n56656), .Y(u_mmu_request_addr_w[17]) );
  INVX1 U60166 ( .A(n56658), .Y(n56660) );
  XNOR2X1 U60167 ( .A(n44837), .B(n56660), .Y(n56659) );
  NAND2X1 U60168 ( .A(n56659), .B(n43375), .Y(n56662) );
  MX2X1 U60169 ( .A(n37555), .B(n42219), .S0(n56660), .Y(n56661) );
  MX2X1 U60170 ( .A(n56662), .B(n56661), .S0(n43931), .Y(u_lsu_mem_addr_r[20])
         );
  NOR2X1 U60171 ( .A(n2383), .B(n40671), .Y(n56664) );
  NOR2X1 U60172 ( .A(n8314), .B(n40686), .Y(n56663) );
  NOR2X1 U60173 ( .A(n56664), .B(n56663), .Y(n56666) );
  NAND2X1 U60174 ( .A(n56767), .B(n7), .Y(n56665) );
  NAND2X1 U60175 ( .A(n56666), .B(n56665), .Y(u_mmu_request_addr_w[20]) );
  INVX1 U60176 ( .A(n56667), .Y(n56669) );
  XNOR2X1 U60177 ( .A(n42852), .B(n56669), .Y(n56668) );
  NAND2X1 U60178 ( .A(n56668), .B(n43375), .Y(n56671) );
  MX2X1 U60179 ( .A(n37555), .B(n42219), .S0(n56669), .Y(n56670) );
  MX2X1 U60180 ( .A(n56671), .B(n56670), .S0(n43902), .Y(u_lsu_mem_addr_r[16])
         );
  NOR2X1 U60181 ( .A(n2516), .B(n40672), .Y(n56673) );
  NOR2X1 U60182 ( .A(n8304), .B(n40687), .Y(n56672) );
  NOR2X1 U60183 ( .A(n56673), .B(n56672), .Y(n56675) );
  NAND2X1 U60184 ( .A(n56767), .B(n8), .Y(n56674) );
  NAND2X1 U60185 ( .A(n56675), .B(n56674), .Y(u_mmu_request_addr_w[16]) );
  INVX1 U60186 ( .A(n56676), .Y(n56678) );
  XNOR2X1 U60187 ( .A(n42852), .B(n56678), .Y(n56677) );
  NAND2X1 U60188 ( .A(n56677), .B(n43374), .Y(n56680) );
  MX2X1 U60189 ( .A(n37555), .B(n42219), .S0(n56678), .Y(n56679) );
  MX2X1 U60190 ( .A(n56680), .B(n56679), .S0(n43988), .Y(u_lsu_mem_addr_r[24])
         );
  NOR2X1 U60191 ( .A(n2850), .B(n40673), .Y(n56682) );
  NOR2X1 U60192 ( .A(n8322), .B(n40688), .Y(n56681) );
  NOR2X1 U60193 ( .A(n56682), .B(n56681), .Y(n56684) );
  NAND2X1 U60194 ( .A(n56767), .B(n11), .Y(n56683) );
  NAND2X1 U60195 ( .A(n56684), .B(n56683), .Y(u_mmu_request_addr_w[24]) );
  MX2X1 U60196 ( .A(u_mmu_itlb_va_addr_q[24]), .B(n57386), .S0(n37548), .Y(
        n8429) );
  INVX1 U60197 ( .A(n56685), .Y(n56687) );
  XNOR2X1 U60198 ( .A(n44838), .B(n56687), .Y(n56686) );
  NAND2X1 U60199 ( .A(n56686), .B(n43374), .Y(n56689) );
  MX2X1 U60200 ( .A(n37555), .B(n42219), .S0(n56687), .Y(n56688) );
  MX2X1 U60201 ( .A(n56689), .B(n56688), .S0(n43939), .Y(u_lsu_mem_addr_r[21])
         );
  NOR2X1 U60202 ( .A(n2549), .B(n40672), .Y(n56691) );
  NOR2X1 U60203 ( .A(n8316), .B(n40687), .Y(n56690) );
  NOR2X1 U60204 ( .A(n56691), .B(n56690), .Y(n56693) );
  NAND2X1 U60205 ( .A(n56767), .B(n12), .Y(n56692) );
  NAND2X1 U60206 ( .A(n56693), .B(n56692), .Y(u_mmu_request_addr_w[21]) );
  INVX1 U60207 ( .A(n56694), .Y(n56696) );
  XNOR2X1 U60208 ( .A(n42852), .B(n56696), .Y(n56695) );
  NAND2X1 U60209 ( .A(n56695), .B(n43374), .Y(n56698) );
  MX2X1 U60210 ( .A(n37555), .B(n42219), .S0(n56696), .Y(n56697) );
  MX2X1 U60211 ( .A(n56698), .B(n56697), .S0(n43978), .Y(u_lsu_mem_addr_r[23])
         );
  NOR2X1 U60212 ( .A(n2451), .B(n40671), .Y(n56700) );
  NOR2X1 U60213 ( .A(n8320), .B(n40686), .Y(n56699) );
  NOR2X1 U60214 ( .A(n56700), .B(n56699), .Y(n56702) );
  NAND2X1 U60215 ( .A(n56767), .B(n15), .Y(n56701) );
  NAND2X1 U60216 ( .A(n56702), .B(n56701), .Y(u_mmu_request_addr_w[23]) );
  MX2X1 U60217 ( .A(u_mmu_itlb_va_addr_q[23]), .B(n57387), .S0(n37548), .Y(
        n8438) );
  INVX1 U60218 ( .A(n56703), .Y(n56705) );
  XNOR2X1 U60219 ( .A(n42851), .B(n56705), .Y(n56704) );
  NAND2X1 U60220 ( .A(n56704), .B(n43374), .Y(n56707) );
  MX2X1 U60221 ( .A(n37555), .B(n42219), .S0(n56705), .Y(n56706) );
  MX2X1 U60222 ( .A(n56707), .B(n56706), .S0(n44021), .Y(u_lsu_mem_addr_r[28])
         );
  NAND2X1 U60223 ( .A(n42253), .B(n56708), .Y(n56710) );
  NAND2X1 U60224 ( .A(n42252), .B(n18), .Y(n56709) );
  NAND2X1 U60225 ( .A(u_mmu_virt_addr_q_28), .B(n57397), .Y(n56711) );
  NAND2X1 U60226 ( .A(n42420), .B(n56711), .Y(n8551) );
  MX2X1 U60227 ( .A(u_mmu_itlb_va_addr_q[28]), .B(u_mmu_virt_addr_q_28), .S0(
        n37548), .Y(n8440) );
  INVX1 U60228 ( .A(n56712), .Y(n56714) );
  XNOR2X1 U60229 ( .A(n42851), .B(n56714), .Y(n56713) );
  NAND2X1 U60230 ( .A(n56713), .B(n43374), .Y(n56716) );
  MX2X1 U60231 ( .A(n37555), .B(n42219), .S0(n56714), .Y(n56715) );
  MX2X1 U60232 ( .A(n56716), .B(n56715), .S0(n43924), .Y(u_lsu_mem_addr_r[19])
         );
  NOR2X1 U60233 ( .A(n2283), .B(n40673), .Y(n56718) );
  NOR2X1 U60234 ( .A(n8310), .B(n40688), .Y(n56717) );
  NOR2X1 U60235 ( .A(n56718), .B(n56717), .Y(n56720) );
  NAND2X1 U60236 ( .A(n56767), .B(n20), .Y(n56719) );
  NAND2X1 U60237 ( .A(n56720), .B(n56719), .Y(u_mmu_request_addr_w[19]) );
  INVX1 U60238 ( .A(n56721), .Y(n56723) );
  XNOR2X1 U60239 ( .A(n44838), .B(n56723), .Y(n56722) );
  NAND2X1 U60240 ( .A(n56722), .B(n43374), .Y(n56725) );
  MX2X1 U60241 ( .A(n37555), .B(n42219), .S0(n56723), .Y(n56724) );
  MX2X1 U60242 ( .A(n56725), .B(n56724), .S0(n43959), .Y(u_lsu_mem_addr_r[12])
         );
  NAND2X1 U60243 ( .A(n29657), .B(n56726), .Y(n17216) );
  NOR2X1 U60244 ( .A(n2683), .B(n40673), .Y(n56728) );
  NOR2X1 U60245 ( .A(n8296), .B(n40688), .Y(n56727) );
  NOR2X1 U60246 ( .A(n56728), .B(n56727), .Y(n56730) );
  NAND2X1 U60247 ( .A(n56767), .B(n21), .Y(n56729) );
  NAND2X1 U60248 ( .A(n56730), .B(n56729), .Y(u_mmu_request_addr_w[12]) );
  INVX1 U60249 ( .A(n56731), .Y(n56733) );
  XNOR2X1 U60250 ( .A(n42852), .B(n56733), .Y(n56732) );
  NAND2X1 U60251 ( .A(n56732), .B(n43374), .Y(n56735) );
  MX2X1 U60252 ( .A(n37555), .B(n42219), .S0(n56733), .Y(n56734) );
  MX2X1 U60253 ( .A(n56735), .B(n56734), .S0(n43895), .Y(u_lsu_mem_addr_r[15])
         );
  NOR2X1 U60254 ( .A(n1869), .B(n40671), .Y(n56737) );
  NOR2X1 U60255 ( .A(n8302), .B(n40686), .Y(n56736) );
  NOR2X1 U60256 ( .A(n56737), .B(n56736), .Y(n56739) );
  NAND2X1 U60257 ( .A(n56767), .B(n22), .Y(n56738) );
  NAND2X1 U60258 ( .A(n56739), .B(n56738), .Y(u_mmu_request_addr_w[15]) );
  INVX1 U60259 ( .A(n56740), .Y(n56742) );
  XNOR2X1 U60260 ( .A(n44837), .B(n56742), .Y(n56741) );
  NAND2X1 U60261 ( .A(n56741), .B(n43374), .Y(n56744) );
  MX2X1 U60262 ( .A(n37555), .B(n42219), .S0(n56742), .Y(n56743) );
  MX2X1 U60263 ( .A(n56744), .B(n56743), .S0(n43886), .Y(u_lsu_mem_addr_r[14])
         );
  NOR2X1 U60264 ( .A(n1797), .B(n40672), .Y(n56746) );
  NOR2X1 U60265 ( .A(n8300), .B(n40687), .Y(n56745) );
  NOR2X1 U60266 ( .A(n56746), .B(n56745), .Y(n56748) );
  NAND2X1 U60267 ( .A(n56767), .B(n24), .Y(n56747) );
  NAND2X1 U60268 ( .A(n56748), .B(n56747), .Y(u_mmu_request_addr_w[14]) );
  INVX1 U60269 ( .A(n56749), .Y(n56751) );
  XNOR2X1 U60270 ( .A(n44838), .B(n56751), .Y(n56750) );
  NAND2X1 U60271 ( .A(n56750), .B(n43374), .Y(n56753) );
  MX2X1 U60272 ( .A(n37555), .B(n42219), .S0(n56751), .Y(n56752) );
  MX2X1 U60273 ( .A(n56753), .B(n56752), .S0(n43915), .Y(u_lsu_mem_addr_r[18])
         );
  NOR2X1 U60274 ( .A(n2650), .B(n40671), .Y(n56755) );
  NOR2X1 U60275 ( .A(n8308), .B(n40686), .Y(n56754) );
  NOR2X1 U60276 ( .A(n56755), .B(n56754), .Y(n56757) );
  NAND2X1 U60277 ( .A(n56767), .B(n10), .Y(n56756) );
  NAND2X1 U60278 ( .A(n56757), .B(n56756), .Y(u_mmu_request_addr_w[18]) );
  INVX1 U60279 ( .A(n56758), .Y(n56760) );
  XNOR2X1 U60280 ( .A(n44837), .B(n56760), .Y(n56759) );
  NAND2X1 U60281 ( .A(n56759), .B(n43374), .Y(n56762) );
  MX2X1 U60282 ( .A(n37555), .B(n42219), .S0(n56760), .Y(n56761) );
  MX2X1 U60283 ( .A(n56762), .B(n56761), .S0(n43875), .Y(u_lsu_mem_addr_r[13])
         );
  NOR2X1 U60284 ( .A(n2753), .B(n40673), .Y(n56766) );
  NOR2X1 U60285 ( .A(n8298), .B(n40688), .Y(n56765) );
  NOR2X1 U60286 ( .A(n56766), .B(n56765), .Y(n56769) );
  NAND2X1 U60287 ( .A(n56767), .B(n9), .Y(n56768) );
  NAND2X1 U60288 ( .A(n56769), .B(n56768), .Y(u_mmu_request_addr_w[13]) );
  NAND2X1 U60289 ( .A(challenge[102]), .B(n44854), .Y(n56770) );
  NAND2X1 U60290 ( .A(n56771), .B(n56770), .Y(n17310) );
  NOR2X1 U60291 ( .A(n1972), .B(n43305), .Y(n56776) );
  NAND2X1 U60292 ( .A(n43307), .B(n56772), .Y(n56775) );
  NAND2X1 U60293 ( .A(n43311), .B(n56773), .Y(n56774) );
  NAND2X1 U60294 ( .A(n56775), .B(n56774), .Y(n56779) );
  NOR2X1 U60295 ( .A(n56776), .B(n56779), .Y(n56778) );
  OR2X1 U60296 ( .A(n1759), .B(n42847), .Y(n56777) );
  NAND2X1 U60297 ( .A(n56778), .B(n56777), .Y(mem_i_pc_o[1]) );
  NOR2X1 U60298 ( .A(n43315), .B(n56781), .Y(net2381) );
  NOR2X1 U60299 ( .A(n1973), .B(n43322), .Y(n56780) );
  NOR2X1 U60300 ( .A(n56780), .B(n56779), .Y(n56786) );
  NOR2X1 U60301 ( .A(n43325), .B(n56781), .Y(n56784) );
  NOR2X1 U60302 ( .A(n56782), .B(n43328), .Y(n56783) );
  NOR2X1 U60303 ( .A(n56784), .B(n56783), .Y(n56785) );
  NAND2X1 U60304 ( .A(n56786), .B(n56785), .Y(u_decode_N291) );
  NOR2X1 U60305 ( .A(n43315), .B(n56789), .Y(net2383) );
  NOR2X1 U60306 ( .A(n2036), .B(n43322), .Y(n56788) );
  NOR2X1 U60307 ( .A(n56788), .B(n56787), .Y(n56794) );
  NOR2X1 U60308 ( .A(n43325), .B(n56789), .Y(n56792) );
  NOR2X1 U60309 ( .A(n43326), .B(n56790), .Y(n56791) );
  NOR2X1 U60310 ( .A(n56792), .B(n56791), .Y(n56793) );
  NAND2X1 U60311 ( .A(n56794), .B(n56793), .Y(u_decode_N293) );
  NAND2X1 U60312 ( .A(n43269), .B(n40393), .Y(n56796) );
  NAND2X1 U60313 ( .A(opcode_pc_w[3]), .B(n56852), .Y(n56795) );
  NAND2X1 U60314 ( .A(n56796), .B(n56795), .Y(n15739) );
  INVX1 U60315 ( .A(n15739), .Y(n73495) );
  NOR2X1 U60316 ( .A(n40674), .B(n73495), .Y(n56800) );
  INVX1 U60317 ( .A(n15463), .Y(n73511) );
  NAND2X1 U60318 ( .A(n56797), .B(n73511), .Y(n56798) );
  NAND2X1 U60319 ( .A(n15668), .B(n56798), .Y(n56799) );
  NOR2X1 U60320 ( .A(n56800), .B(n56799), .Y(n56803) );
  OR2X1 U60321 ( .A(n15701), .B(n15700), .Y(n56801) );
  NOR2X1 U60322 ( .A(n15666), .B(n56801), .Y(n56802) );
  NAND2X1 U60323 ( .A(n56803), .B(n56802), .Y(u_exec_alu_p_w[4]) );
  NOR2X1 U60324 ( .A(n22667), .B(n43262), .Y(n56805) );
  NOR2X1 U60325 ( .A(n44363), .B(n43265), .Y(n56804) );
  NOR2X1 U60326 ( .A(n56805), .B(n56804), .Y(n56807) );
  NOR2X1 U60327 ( .A(n22850), .B(n22849), .Y(n56806) );
  NAND2X1 U60328 ( .A(n56807), .B(n56806), .Y(u_decode_u_regfile_N1214) );
  NOR2X1 U60329 ( .A(n43315), .B(n56811), .Y(net2388) );
  NOR2X1 U60330 ( .A(n43326), .B(n56808), .Y(n56810) );
  NOR2X1 U60331 ( .A(n56810), .B(n56809), .Y(n56815) );
  NOR2X1 U60332 ( .A(n2137), .B(n43322), .Y(n56813) );
  NOR2X1 U60333 ( .A(n43325), .B(n56811), .Y(n56812) );
  NOR2X1 U60334 ( .A(n56813), .B(n56812), .Y(n56814) );
  NAND2X1 U60335 ( .A(n56815), .B(n56814), .Y(u_decode_N298) );
  NAND2X1 U60336 ( .A(n43269), .B(n44038), .Y(n56817) );
  NAND2X1 U60337 ( .A(opcode_pc_w[8]), .B(n40680), .Y(n56816) );
  NAND2X1 U60338 ( .A(n56817), .B(n56816), .Y(n15447) );
  NAND2X1 U60339 ( .A(n43410), .B(n43737), .Y(n56819) );
  INVX1 U60340 ( .A(n58548), .Y(n58554) );
  NAND2X1 U60341 ( .A(n58554), .B(opcode_opcode_w[28]), .Y(n56818) );
  NAND2X1 U60342 ( .A(n56819), .B(n56818), .Y(n17354) );
  INVX1 U60343 ( .A(n15447), .Y(n73494) );
  NAND2X1 U60344 ( .A(n17354), .B(n73494), .Y(n17541) );
  NAND2X1 U60345 ( .A(n43269), .B(n42715), .Y(n56821) );
  NAND2X1 U60346 ( .A(opcode_pc_w[1]), .B(n56852), .Y(n56820) );
  NAND2X1 U60347 ( .A(n56821), .B(n56820), .Y(n16596) );
  NAND2X1 U60348 ( .A(n43269), .B(n43457), .Y(n56823) );
  NAND2X1 U60349 ( .A(opcode_pc_w[2]), .B(n40680), .Y(n56822) );
  NAND2X1 U60350 ( .A(n56823), .B(n56822), .Y(n15919) );
  INVX1 U60351 ( .A(n56824), .Y(n56826) );
  NOR2X1 U60352 ( .A(n56826), .B(n56825), .Y(n56828) );
  NAND2X1 U60353 ( .A(n43410), .B(n43816), .Y(n56827) );
  NAND2X1 U60354 ( .A(n56828), .B(n56827), .Y(n15734) );
  NAND2X1 U60355 ( .A(n43269), .B(n43466), .Y(n56830) );
  NAND2X1 U60356 ( .A(opcode_pc_w[4]), .B(n40679), .Y(n56829) );
  NAND2X1 U60357 ( .A(n56830), .B(n56829), .Y(n15679) );
  NAND2X1 U60358 ( .A(n43410), .B(n39525), .Y(n56833) );
  NAND2X1 U60359 ( .A(n42747), .B(n56831), .Y(n56832) );
  NAND2X1 U60360 ( .A(n56833), .B(n56832), .Y(n15682) );
  NAND2X1 U60361 ( .A(n43269), .B(n39943), .Y(n56835) );
  NAND2X1 U60362 ( .A(opcode_pc_w[5]), .B(n40680), .Y(n56834) );
  NAND2X1 U60363 ( .A(n56835), .B(n56834), .Y(n17094) );
  NAND2X1 U60364 ( .A(n43410), .B(n38611), .Y(n56837) );
  NAND2X1 U60365 ( .A(n58554), .B(opcode_opcode_w[25]), .Y(n56836) );
  NAND2X1 U60366 ( .A(n56837), .B(n56836), .Y(n15633) );
  NAND2X1 U60367 ( .A(n43269), .B(n43843), .Y(n56839) );
  NAND2X1 U60368 ( .A(opcode_pc_w[6]), .B(n56852), .Y(n56838) );
  NAND2X1 U60369 ( .A(n56839), .B(n56838), .Y(n15443) );
  NAND2X1 U60370 ( .A(n43410), .B(n43792), .Y(n56841) );
  NAND2X1 U60371 ( .A(n58554), .B(opcode_opcode_w[26]), .Y(n56840) );
  NAND2X1 U60372 ( .A(n56841), .B(n56840), .Y(n17361) );
  INVX1 U60373 ( .A(n17361), .Y(n73485) );
  NAND2X1 U60374 ( .A(n15443), .B(n73485), .Y(n15567) );
  NAND2X1 U60375 ( .A(n43268), .B(n38383), .Y(n56843) );
  NAND2X1 U60376 ( .A(opcode_pc_w[7]), .B(n40679), .Y(n56842) );
  NAND2X1 U60377 ( .A(n56843), .B(n56842), .Y(n15441) );
  NAND2X1 U60378 ( .A(n43409), .B(n43780), .Y(n56845) );
  NAND2X1 U60379 ( .A(n58554), .B(opcode_opcode_w[27]), .Y(n56844) );
  NAND2X1 U60380 ( .A(n56845), .B(n56844), .Y(n15524) );
  INVX1 U60381 ( .A(n17354), .Y(n73493) );
  NAND2X1 U60382 ( .A(n15447), .B(n73493), .Y(n15476) );
  NAND2X1 U60383 ( .A(n43268), .B(n43853), .Y(n56847) );
  NAND2X1 U60384 ( .A(opcode_pc_w[9]), .B(n56852), .Y(n56846) );
  NAND2X1 U60385 ( .A(n56847), .B(n56846), .Y(n15414) );
  NAND2X1 U60386 ( .A(n43409), .B(n43758), .Y(n56849) );
  NAND2X1 U60387 ( .A(n58554), .B(opcode_opcode_w[29]), .Y(n56848) );
  NAND2X1 U60388 ( .A(n56849), .B(n56848), .Y(n15420) );
  NAND2X1 U60389 ( .A(n43268), .B(n43862), .Y(n56851) );
  NAND2X1 U60390 ( .A(opcode_pc_w[10]), .B(n40679), .Y(n56850) );
  NAND2X1 U60391 ( .A(n56851), .B(n56850), .Y(n15845) );
  NAND2X1 U60392 ( .A(n43409), .B(n43820), .Y(n58561) );
  NAND2X1 U60393 ( .A(n58554), .B(opcode_opcode_w[30]), .Y(n58560) );
  NAND2X1 U60394 ( .A(n58561), .B(n58560), .Y(n330) );
  INVX1 U60395 ( .A(n330), .Y(n73479) );
  NAND2X1 U60396 ( .A(n15845), .B(n73479), .Y(n17203) );
  NAND2X1 U60397 ( .A(n43268), .B(n43965), .Y(n56854) );
  NAND2X1 U60398 ( .A(opcode_pc_w[11]), .B(n56852), .Y(n56853) );
  NAND2X1 U60399 ( .A(n56854), .B(n56853), .Y(n15728) );
  NAND2X1 U60400 ( .A(n43409), .B(n43812), .Y(n56855) );
  NAND2X1 U60401 ( .A(n58554), .B(n44835), .Y(n57001) );
  NAND2X1 U60402 ( .A(n56855), .B(n57001), .Y(n318) );
  NOR2X1 U60403 ( .A(n42940), .B(n58291), .Y(n56857) );
  NOR2X1 U60404 ( .A(n56860), .B(n42937), .Y(n56856) );
  NOR2X1 U60405 ( .A(n56857), .B(n56856), .Y(n56859) );
  NAND2X1 U60406 ( .A(n43268), .B(n43955), .Y(n56858) );
  NAND2X1 U60407 ( .A(n56859), .B(n56858), .Y(n16042) );
  INVX1 U60408 ( .A(n57001), .Y(n56986) );
  NOR2X1 U60409 ( .A(n56860), .B(n42935), .Y(n56861) );
  NOR2X1 U60410 ( .A(n56986), .B(n56861), .Y(n56863) );
  NAND2X1 U60411 ( .A(n43409), .B(n40463), .Y(n56862) );
  NAND2X1 U60412 ( .A(n56863), .B(n56862), .Y(n17017) );
  NOR2X1 U60413 ( .A(n42941), .B(n58298), .Y(n56865) );
  NOR2X1 U60414 ( .A(n56868), .B(n42938), .Y(n56864) );
  NOR2X1 U60415 ( .A(n56865), .B(n56864), .Y(n56867) );
  NAND2X1 U60416 ( .A(n43268), .B(n43872), .Y(n56866) );
  NAND2X1 U60417 ( .A(n56867), .B(n56866), .Y(n15977) );
  NOR2X1 U60418 ( .A(n56868), .B(n42936), .Y(n56869) );
  NOR2X1 U60419 ( .A(n56986), .B(n56869), .Y(n56871) );
  NAND2X1 U60420 ( .A(n43409), .B(n40471), .Y(n56870) );
  NAND2X1 U60421 ( .A(n56871), .B(n56870), .Y(n16952) );
  NOR2X1 U60422 ( .A(n42939), .B(n58305), .Y(n56873) );
  NOR2X1 U60423 ( .A(n56876), .B(n56993), .Y(n56872) );
  NOR2X1 U60424 ( .A(n56873), .B(n56872), .Y(n56875) );
  NAND2X1 U60425 ( .A(n43268), .B(n43882), .Y(n56874) );
  NAND2X1 U60426 ( .A(n56875), .B(n56874), .Y(n15846) );
  NOR2X1 U60427 ( .A(n56876), .B(n56998), .Y(n56877) );
  NOR2X1 U60428 ( .A(n56986), .B(n56877), .Y(n56879) );
  NAND2X1 U60429 ( .A(n43409), .B(n40484), .Y(n56878) );
  NAND2X1 U60430 ( .A(n56879), .B(n56878), .Y(n16891) );
  NOR2X1 U60431 ( .A(n42940), .B(n58312), .Y(n56881) );
  NOR2X1 U60432 ( .A(n42730), .B(n42937), .Y(n56880) );
  NOR2X1 U60433 ( .A(n56881), .B(n56880), .Y(n56883) );
  NAND2X1 U60434 ( .A(n43268), .B(n43892), .Y(n56882) );
  NAND2X1 U60435 ( .A(n56883), .B(n56882), .Y(n15805) );
  NOR2X1 U60436 ( .A(n42732), .B(n42935), .Y(n56884) );
  NOR2X1 U60437 ( .A(n56986), .B(n56884), .Y(n56886) );
  NAND2X1 U60438 ( .A(n43409), .B(n43787), .Y(n56885) );
  NAND2X1 U60439 ( .A(n56886), .B(n56885), .Y(n16844) );
  NOR2X1 U60440 ( .A(n42941), .B(n58319), .Y(n56888) );
  NOR2X1 U60441 ( .A(n42727), .B(n42938), .Y(n56887) );
  NOR2X1 U60442 ( .A(n56888), .B(n56887), .Y(n56890) );
  NAND2X1 U60443 ( .A(n43268), .B(n43899), .Y(n56889) );
  NAND2X1 U60444 ( .A(n56890), .B(n56889), .Y(n16775) );
  NOR2X1 U60445 ( .A(n42725), .B(n42936), .Y(n56891) );
  NOR2X1 U60446 ( .A(n56986), .B(n56891), .Y(n56893) );
  NAND2X1 U60447 ( .A(n43409), .B(n43725), .Y(n56892) );
  NAND2X1 U60448 ( .A(n56893), .B(n56892), .Y(n16792) );
  NOR2X1 U60449 ( .A(n42939), .B(n58324), .Y(n56895) );
  NOR2X1 U60450 ( .A(n42689), .B(n56993), .Y(n56894) );
  NOR2X1 U60451 ( .A(n56895), .B(n56894), .Y(n56897) );
  NAND2X1 U60452 ( .A(n43268), .B(n43906), .Y(n56896) );
  NAND2X1 U60453 ( .A(n56897), .B(n56896), .Y(n16563) );
  NOR2X1 U60454 ( .A(n42689), .B(n56998), .Y(n56898) );
  NOR2X1 U60455 ( .A(n56986), .B(n56898), .Y(n56900) );
  NAND2X1 U60456 ( .A(n43409), .B(n42632), .Y(n56899) );
  NAND2X1 U60457 ( .A(n56900), .B(n56899), .Y(n16739) );
  NOR2X1 U60458 ( .A(n42940), .B(n58331), .Y(n56902) );
  NOR2X1 U60459 ( .A(n42665), .B(n42937), .Y(n56901) );
  NOR2X1 U60460 ( .A(n56902), .B(n56901), .Y(n56904) );
  NAND2X1 U60461 ( .A(n43268), .B(n43912), .Y(n56903) );
  NAND2X1 U60462 ( .A(n56904), .B(n56903), .Y(n16181) );
  NOR2X1 U60463 ( .A(n42663), .B(n42935), .Y(n56905) );
  NOR2X1 U60464 ( .A(n56986), .B(n56905), .Y(n56907) );
  NAND2X1 U60465 ( .A(n43409), .B(n40260), .Y(n56906) );
  NAND2X1 U60466 ( .A(n56907), .B(n56906), .Y(n16685) );
  NOR2X1 U60467 ( .A(n42941), .B(n58338), .Y(n56909) );
  NOR2X1 U60468 ( .A(n42787), .B(n42938), .Y(n56908) );
  NOR2X1 U60469 ( .A(n56909), .B(n56908), .Y(n56911) );
  NAND2X1 U60470 ( .A(n43268), .B(n43921), .Y(n56910) );
  NAND2X1 U60471 ( .A(n56911), .B(n56910), .Y(n15801) );
  NOR2X1 U60472 ( .A(n42786), .B(n42936), .Y(n56912) );
  NOR2X1 U60473 ( .A(n56986), .B(n56912), .Y(n56914) );
  NAND2X1 U60474 ( .A(n43408), .B(n43799), .Y(n56913) );
  NAND2X1 U60475 ( .A(n56914), .B(n56913), .Y(n16557) );
  NOR2X1 U60476 ( .A(n42939), .B(n58344), .Y(n56916) );
  NOR2X1 U60477 ( .A(n39116), .B(n56993), .Y(n56915) );
  NOR2X1 U60478 ( .A(n56916), .B(n56915), .Y(n56918) );
  NAND2X1 U60479 ( .A(n43267), .B(n43929), .Y(n56917) );
  NAND2X1 U60480 ( .A(n56918), .B(n56917), .Y(n16048) );
  NOR2X1 U60481 ( .A(n42739), .B(n56998), .Y(n56919) );
  NOR2X1 U60482 ( .A(n56986), .B(n56919), .Y(n56921) );
  NAND2X1 U60483 ( .A(n43408), .B(n42661), .Y(n56920) );
  NAND2X1 U60484 ( .A(n56921), .B(n56920), .Y(n16504) );
  NOR2X1 U60485 ( .A(n42940), .B(n58349), .Y(n56923) );
  NOR2X1 U60486 ( .A(n42468), .B(n42937), .Y(n56922) );
  NOR2X1 U60487 ( .A(n56923), .B(n56922), .Y(n56925) );
  NAND2X1 U60488 ( .A(n43267), .B(n43936), .Y(n56924) );
  NAND2X1 U60489 ( .A(n56925), .B(n56924), .Y(n16449) );
  NOR2X1 U60490 ( .A(n42468), .B(n42935), .Y(n56926) );
  NOR2X1 U60491 ( .A(n56986), .B(n56926), .Y(n56928) );
  NAND2X1 U60492 ( .A(n43408), .B(n42712), .Y(n56927) );
  NAND2X1 U60493 ( .A(n56928), .B(n56927), .Y(n16450) );
  NOR2X1 U60494 ( .A(n42941), .B(n58356), .Y(n56930) );
  NOR2X1 U60495 ( .A(n39640), .B(n42938), .Y(n56929) );
  NOR2X1 U60496 ( .A(n56930), .B(n56929), .Y(n56932) );
  NAND2X1 U60497 ( .A(n43267), .B(n43945), .Y(n56931) );
  NAND2X1 U60498 ( .A(n56932), .B(n56931), .Y(n16290) );
  NOR2X1 U60499 ( .A(n39640), .B(n42936), .Y(n56933) );
  NOR2X1 U60500 ( .A(n56986), .B(n56933), .Y(n56935) );
  NAND2X1 U60501 ( .A(n43408), .B(n43795), .Y(n56934) );
  NAND2X1 U60502 ( .A(n56935), .B(n56934), .Y(n16396) );
  NOR2X1 U60503 ( .A(n42939), .B(n58363), .Y(n56937) );
  NOR2X1 U60504 ( .A(n42760), .B(n56993), .Y(n56936) );
  NOR2X1 U60505 ( .A(n56937), .B(n56936), .Y(n56939) );
  NAND2X1 U60506 ( .A(n43267), .B(n43975), .Y(n56938) );
  NAND2X1 U60507 ( .A(n56939), .B(n56938), .Y(n15802) );
  NOR2X1 U60508 ( .A(n42760), .B(n56998), .Y(n56940) );
  NOR2X1 U60509 ( .A(n56986), .B(n56940), .Y(n56942) );
  NAND2X1 U60510 ( .A(n43409), .B(n43776), .Y(n56941) );
  NAND2X1 U60511 ( .A(n56942), .B(n56941), .Y(n16338) );
  NOR2X1 U60512 ( .A(n42940), .B(n58370), .Y(n56944) );
  NOR2X1 U60513 ( .A(n42749), .B(n42937), .Y(n56943) );
  NOR2X1 U60514 ( .A(n56944), .B(n56943), .Y(n56946) );
  NAND2X1 U60515 ( .A(n43267), .B(n43985), .Y(n56945) );
  NAND2X1 U60516 ( .A(n56946), .B(n56945), .Y(n16047) );
  NOR2X1 U60517 ( .A(n42749), .B(n42935), .Y(n56947) );
  NOR2X1 U60518 ( .A(n56986), .B(n56947), .Y(n56949) );
  NAND2X1 U60519 ( .A(n43408), .B(n43479), .Y(n56948) );
  NAND2X1 U60520 ( .A(n56949), .B(n56948), .Y(n16278) );
  NOR2X1 U60521 ( .A(n42941), .B(n58377), .Y(n56951) );
  NOR2X1 U60522 ( .A(n58817), .B(n42938), .Y(n56950) );
  NOR2X1 U60523 ( .A(n56951), .B(n56950), .Y(n56953) );
  NAND2X1 U60524 ( .A(n43267), .B(n43994), .Y(n56952) );
  NAND2X1 U60525 ( .A(n56953), .B(n56952), .Y(n16213) );
  NOR2X1 U60526 ( .A(n58817), .B(n42936), .Y(n56954) );
  NOR2X1 U60527 ( .A(n56986), .B(n56954), .Y(n56956) );
  NAND2X1 U60528 ( .A(n43408), .B(n38312), .Y(n56955) );
  NAND2X1 U60529 ( .A(n56956), .B(n56955), .Y(n16214) );
  NOR2X1 U60530 ( .A(n42939), .B(n58382), .Y(n56958) );
  NOR2X1 U60531 ( .A(n73364), .B(n56993), .Y(n56957) );
  NOR2X1 U60532 ( .A(n56958), .B(n56957), .Y(n56960) );
  NAND2X1 U60533 ( .A(n43267), .B(n44002), .Y(n56959) );
  NAND2X1 U60534 ( .A(n56960), .B(n56959), .Y(n16143) );
  NOR2X1 U60535 ( .A(n73364), .B(n56998), .Y(n56961) );
  NOR2X1 U60536 ( .A(n56986), .B(n56961), .Y(n56963) );
  NAND2X1 U60537 ( .A(n43408), .B(n38311), .Y(n56962) );
  NAND2X1 U60538 ( .A(n56963), .B(n56962), .Y(n16144) );
  NOR2X1 U60539 ( .A(n42940), .B(n58389), .Y(n56965) );
  NOR2X1 U60540 ( .A(n58818), .B(n42937), .Y(n56964) );
  NOR2X1 U60541 ( .A(n56965), .B(n56964), .Y(n56967) );
  NAND2X1 U60542 ( .A(n43267), .B(n44010), .Y(n56966) );
  NAND2X1 U60543 ( .A(n56967), .B(n56966), .Y(n16077) );
  NOR2X1 U60544 ( .A(n58818), .B(n42935), .Y(n56968) );
  NOR2X1 U60545 ( .A(n56986), .B(n56968), .Y(n56970) );
  NAND2X1 U60546 ( .A(n43408), .B(n43493), .Y(n56969) );
  NAND2X1 U60547 ( .A(n56970), .B(n56969), .Y(n16078) );
  NOR2X1 U60548 ( .A(n42941), .B(n58396), .Y(n56972) );
  NOR2X1 U60549 ( .A(n58457), .B(n42938), .Y(n56971) );
  NOR2X1 U60550 ( .A(n56972), .B(n56971), .Y(n56974) );
  NAND2X1 U60551 ( .A(n43267), .B(n44019), .Y(n56973) );
  NAND2X1 U60552 ( .A(n56974), .B(n56973), .Y(n16003) );
  NOR2X1 U60553 ( .A(n58457), .B(n42936), .Y(n56975) );
  NOR2X1 U60554 ( .A(n56986), .B(n56975), .Y(n56977) );
  NAND2X1 U60555 ( .A(n43408), .B(n43497), .Y(n56976) );
  NAND2X1 U60556 ( .A(n56977), .B(n56976), .Y(n16004) );
  NOR2X1 U60557 ( .A(n42939), .B(n58403), .Y(n56979) );
  NOR2X1 U60558 ( .A(n73367), .B(n56993), .Y(n56978) );
  NOR2X1 U60559 ( .A(n56979), .B(n56978), .Y(n56981) );
  NAND2X1 U60560 ( .A(n43267), .B(n44027), .Y(n56980) );
  NAND2X1 U60561 ( .A(n56981), .B(n56980), .Y(n15874) );
  NOR2X1 U60562 ( .A(n73367), .B(n56998), .Y(n56982) );
  NOR2X1 U60563 ( .A(n56986), .B(n56982), .Y(n56984) );
  NAND2X1 U60564 ( .A(n43408), .B(n43502), .Y(n56983) );
  NAND2X1 U60565 ( .A(n56984), .B(n56983), .Y(n15875) );
  NOR2X1 U60566 ( .A(n57889), .B(n42935), .Y(n56985) );
  NOR2X1 U60567 ( .A(n56986), .B(n56985), .Y(n56988) );
  NAND2X1 U60568 ( .A(n43408), .B(n39844), .Y(n56987) );
  NAND2X1 U60569 ( .A(n56988), .B(n56987), .Y(n15810) );
  NOR2X1 U60570 ( .A(n42940), .B(n58409), .Y(n56990) );
  NOR2X1 U60571 ( .A(n57889), .B(n42937), .Y(n56989) );
  NOR2X1 U60572 ( .A(n56990), .B(n56989), .Y(n56992) );
  NAND2X1 U60573 ( .A(n43267), .B(n44050), .Y(n56991) );
  NAND2X1 U60574 ( .A(n56992), .B(n56991), .Y(n15862) );
  NOR2X1 U60575 ( .A(n42941), .B(n58416), .Y(n56995) );
  NOR2X1 U60576 ( .A(n44842), .B(n42938), .Y(n56994) );
  NOR2X1 U60577 ( .A(n56995), .B(n56994), .Y(n56997) );
  NAND2X1 U60578 ( .A(n43267), .B(n44057), .Y(n56996) );
  NAND2X1 U60579 ( .A(n56997), .B(n56996), .Y(n58580) );
  INVX1 U60580 ( .A(n58580), .Y(n73438) );
  NOR2X1 U60581 ( .A(n44841), .B(n42936), .Y(n57000) );
  NOR2X1 U60582 ( .A(n39083), .B(n43411), .Y(n56999) );
  NOR2X1 U60583 ( .A(n57000), .B(n56999), .Y(n57002) );
  NAND2X1 U60584 ( .A(n57002), .B(n57001), .Y(n57323) );
  INVX1 U60585 ( .A(n57323), .Y(n73437) );
  XNOR2X1 U60586 ( .A(n73438), .B(n73437), .Y(n58760) );
  INVX1 U60587 ( .A(n15862), .Y(n73439) );
  NOR2X1 U60588 ( .A(n15810), .B(n73439), .Y(n57086) );
  INVX1 U60589 ( .A(n15875), .Y(n73441) );
  NAND2X1 U60590 ( .A(n15874), .B(n73441), .Y(n57085) );
  INVX1 U60591 ( .A(n15874), .Y(n73442) );
  NAND2X1 U60592 ( .A(n15875), .B(n73442), .Y(n57083) );
  INVX1 U60593 ( .A(n16004), .Y(n73443) );
  NAND2X1 U60594 ( .A(n16003), .B(n73443), .Y(n57082) );
  INVX1 U60595 ( .A(n16003), .Y(n73444) );
  NAND2X1 U60596 ( .A(n16004), .B(n73444), .Y(n57080) );
  INVX1 U60597 ( .A(n16078), .Y(n73445) );
  NAND2X1 U60598 ( .A(n16077), .B(n73445), .Y(n57079) );
  INVX1 U60599 ( .A(n16077), .Y(n73446) );
  NAND2X1 U60600 ( .A(n16078), .B(n73446), .Y(n57077) );
  INVX1 U60601 ( .A(n16144), .Y(n73447) );
  NAND2X1 U60602 ( .A(n16143), .B(n73447), .Y(n57076) );
  INVX1 U60603 ( .A(n16143), .Y(n73448) );
  NAND2X1 U60604 ( .A(n16144), .B(n73448), .Y(n57074) );
  INVX1 U60605 ( .A(n16214), .Y(n73449) );
  NAND2X1 U60606 ( .A(n16213), .B(n73449), .Y(n57073) );
  INVX1 U60607 ( .A(n16213), .Y(n73450) );
  NAND2X1 U60608 ( .A(n16214), .B(n73450), .Y(n57071) );
  INVX1 U60609 ( .A(n16278), .Y(n73451) );
  NAND2X1 U60610 ( .A(n16047), .B(n73451), .Y(n57070) );
  INVX1 U60611 ( .A(n16047), .Y(n73452) );
  NAND2X1 U60612 ( .A(n16278), .B(n73452), .Y(n57068) );
  INVX1 U60613 ( .A(n16338), .Y(n73453) );
  NAND2X1 U60614 ( .A(n15802), .B(n73453), .Y(n57067) );
  INVX1 U60615 ( .A(n15802), .Y(n73454) );
  NAND2X1 U60616 ( .A(n16338), .B(n73454), .Y(n57065) );
  INVX1 U60617 ( .A(n16396), .Y(n73455) );
  NAND2X1 U60618 ( .A(n16290), .B(n73455), .Y(n57064) );
  INVX1 U60619 ( .A(n16290), .Y(n73456) );
  NAND2X1 U60620 ( .A(n16396), .B(n73456), .Y(n57062) );
  INVX1 U60621 ( .A(n16450), .Y(n73457) );
  NAND2X1 U60622 ( .A(n16449), .B(n73457), .Y(n57061) );
  INVX1 U60623 ( .A(n16449), .Y(n73458) );
  NAND2X1 U60624 ( .A(n16450), .B(n73458), .Y(n57059) );
  INVX1 U60625 ( .A(n16504), .Y(n73459) );
  NAND2X1 U60626 ( .A(n16048), .B(n73459), .Y(n57058) );
  INVX1 U60627 ( .A(n16048), .Y(n73460) );
  NAND2X1 U60628 ( .A(n16504), .B(n73460), .Y(n57056) );
  INVX1 U60629 ( .A(n16557), .Y(n73461) );
  NAND2X1 U60630 ( .A(n15801), .B(n73461), .Y(n57055) );
  INVX1 U60631 ( .A(n15801), .Y(n73462) );
  NAND2X1 U60632 ( .A(n16557), .B(n73462), .Y(n57053) );
  INVX1 U60633 ( .A(n16685), .Y(n73463) );
  NAND2X1 U60634 ( .A(n16181), .B(n73463), .Y(n57052) );
  INVX1 U60635 ( .A(n16181), .Y(n73464) );
  NAND2X1 U60636 ( .A(n16685), .B(n73464), .Y(n57050) );
  INVX1 U60637 ( .A(n16739), .Y(n73465) );
  NAND2X1 U60638 ( .A(n16563), .B(n73465), .Y(n57049) );
  INVX1 U60639 ( .A(n16563), .Y(n73466) );
  NAND2X1 U60640 ( .A(n16739), .B(n73466), .Y(n57047) );
  INVX1 U60641 ( .A(n16792), .Y(n73467) );
  NAND2X1 U60642 ( .A(n16775), .B(n73467), .Y(n57046) );
  INVX1 U60643 ( .A(n16775), .Y(n73468) );
  NAND2X1 U60644 ( .A(n16792), .B(n73468), .Y(n57044) );
  INVX1 U60645 ( .A(n16844), .Y(n73469) );
  NAND2X1 U60646 ( .A(n15805), .B(n73469), .Y(n57043) );
  INVX1 U60647 ( .A(n15805), .Y(n73470) );
  NAND2X1 U60648 ( .A(n16844), .B(n73470), .Y(n57041) );
  INVX1 U60649 ( .A(n16891), .Y(n73471) );
  NAND2X1 U60650 ( .A(n15846), .B(n73471), .Y(n57040) );
  INVX1 U60651 ( .A(n15846), .Y(n73472) );
  NAND2X1 U60652 ( .A(n16891), .B(n73472), .Y(n57038) );
  INVX1 U60653 ( .A(n16952), .Y(n73473) );
  NAND2X1 U60654 ( .A(n15977), .B(n73473), .Y(n57037) );
  INVX1 U60655 ( .A(n15977), .Y(n73474) );
  NAND2X1 U60656 ( .A(n16952), .B(n73474), .Y(n57035) );
  INVX1 U60657 ( .A(n17017), .Y(n73475) );
  NAND2X1 U60658 ( .A(n16042), .B(n73475), .Y(n57034) );
  INVX1 U60659 ( .A(n16042), .Y(n73476) );
  NAND2X1 U60660 ( .A(n17017), .B(n73476), .Y(n57032) );
  INVX1 U60661 ( .A(n318), .Y(n73477) );
  NAND2X1 U60662 ( .A(n15728), .B(n73477), .Y(n57031) );
  INVX1 U60663 ( .A(n15728), .Y(n73478) );
  NAND2X1 U60664 ( .A(n318), .B(n73478), .Y(n57029) );
  INVX1 U60665 ( .A(n15845), .Y(n73480) );
  NAND2X1 U60666 ( .A(n330), .B(n73480), .Y(n57027) );
  INVX1 U60667 ( .A(n15420), .Y(n73481) );
  NAND2X1 U60668 ( .A(n15414), .B(n73481), .Y(n57026) );
  INVX1 U60669 ( .A(n15414), .Y(n73482) );
  NAND2X1 U60670 ( .A(n15420), .B(n73482), .Y(n57024) );
  INVX1 U60671 ( .A(n15524), .Y(n73483) );
  NAND2X1 U60672 ( .A(n15441), .B(n73483), .Y(n57022) );
  INVX1 U60673 ( .A(n15441), .Y(n73484) );
  NAND2X1 U60674 ( .A(n15524), .B(n73484), .Y(n57020) );
  INVX1 U60675 ( .A(n15443), .Y(n73486) );
  NAND2X1 U60676 ( .A(n17361), .B(n73486), .Y(n57018) );
  INVX1 U60677 ( .A(n15633), .Y(n73487) );
  NAND2X1 U60678 ( .A(n17094), .B(n73487), .Y(n57017) );
  INVX1 U60679 ( .A(n17094), .Y(n73488) );
  NAND2X1 U60680 ( .A(n15633), .B(n73488), .Y(n57015) );
  INVX1 U60681 ( .A(n15682), .Y(n73489) );
  NAND2X1 U60682 ( .A(n15679), .B(n73489), .Y(n57014) );
  INVX1 U60683 ( .A(n15679), .Y(n73490) );
  NAND2X1 U60684 ( .A(n15682), .B(n73490), .Y(n57012) );
  NAND2X1 U60685 ( .A(n15739), .B(n73525), .Y(n57011) );
  NAND2X1 U60686 ( .A(n15742), .B(n73495), .Y(n57009) );
  INVX1 U60687 ( .A(n15734), .Y(n73433) );
  NAND2X1 U60688 ( .A(n15919), .B(n73433), .Y(n57008) );
  INVX1 U60689 ( .A(n15919), .Y(n73491) );
  NAND2X1 U60690 ( .A(n15734), .B(n73491), .Y(n57006) );
  NAND2X1 U60691 ( .A(n16596), .B(n73523), .Y(n57005) );
  INVX1 U60692 ( .A(n16596), .Y(n73492) );
  NAND2X1 U60693 ( .A(n16593), .B(n73492), .Y(n57003) );
  INVX1 U60694 ( .A(n58597), .Y(n58577) );
  NAND2X1 U60695 ( .A(n58577), .B(n57316), .Y(n58659) );
  NAND2X1 U60696 ( .A(n57003), .B(n58659), .Y(n57004) );
  NAND2X1 U60697 ( .A(n57005), .B(n57004), .Y(n58746) );
  NAND2X1 U60698 ( .A(n57006), .B(n58746), .Y(n57007) );
  NAND2X1 U60699 ( .A(n57008), .B(n57007), .Y(n58765) );
  NAND2X1 U60700 ( .A(n57009), .B(n58765), .Y(n57010) );
  NAND2X1 U60701 ( .A(n57011), .B(n57010), .Y(n58772) );
  NAND2X1 U60702 ( .A(n57012), .B(n58772), .Y(n57013) );
  NAND2X1 U60703 ( .A(n57014), .B(n57013), .Y(n58779) );
  NAND2X1 U60704 ( .A(n57015), .B(n58779), .Y(n57016) );
  NAND2X1 U60705 ( .A(n57017), .B(n57016), .Y(n58785) );
  NAND2X1 U60706 ( .A(n57018), .B(n58785), .Y(n57019) );
  NAND2X1 U60707 ( .A(n57019), .B(n15567), .Y(n58791) );
  NAND2X1 U60708 ( .A(n57020), .B(n58791), .Y(n57021) );
  NAND2X1 U60709 ( .A(n57022), .B(n57021), .Y(n58798) );
  NAND2X1 U60710 ( .A(n58798), .B(n17541), .Y(n57023) );
  NAND2X1 U60711 ( .A(n57023), .B(n15476), .Y(n58808) );
  NAND2X1 U60712 ( .A(n57024), .B(n58808), .Y(n57025) );
  NAND2X1 U60713 ( .A(n57026), .B(n57025), .Y(n58573) );
  NAND2X1 U60714 ( .A(n57027), .B(n58573), .Y(n57028) );
  NAND2X1 U60715 ( .A(n57028), .B(n17203), .Y(n58581) );
  NAND2X1 U60716 ( .A(n57029), .B(n58581), .Y(n57030) );
  NAND2X1 U60717 ( .A(n57031), .B(n57030), .Y(n58589) );
  NAND2X1 U60718 ( .A(n57032), .B(n58589), .Y(n57033) );
  NAND2X1 U60719 ( .A(n57034), .B(n57033), .Y(n58600) );
  NAND2X1 U60720 ( .A(n57035), .B(n58600), .Y(n57036) );
  NAND2X1 U60721 ( .A(n57037), .B(n57036), .Y(n58611) );
  NAND2X1 U60722 ( .A(n57038), .B(n58611), .Y(n57039) );
  NAND2X1 U60723 ( .A(n57040), .B(n57039), .Y(n58614) );
  NAND2X1 U60724 ( .A(n57041), .B(n58614), .Y(n57042) );
  NAND2X1 U60725 ( .A(n57043), .B(n57042), .Y(n58622) );
  NAND2X1 U60726 ( .A(n57044), .B(n58622), .Y(n57045) );
  NAND2X1 U60727 ( .A(n57046), .B(n57045), .Y(n58630) );
  NAND2X1 U60728 ( .A(n57047), .B(n58630), .Y(n57048) );
  NAND2X1 U60729 ( .A(n57049), .B(n57048), .Y(n58638) );
  NAND2X1 U60730 ( .A(n57050), .B(n58638), .Y(n57051) );
  NAND2X1 U60731 ( .A(n57052), .B(n57051), .Y(n58646) );
  NAND2X1 U60732 ( .A(n57053), .B(n58646), .Y(n57054) );
  NAND2X1 U60733 ( .A(n57055), .B(n57054), .Y(n58662) );
  NAND2X1 U60734 ( .A(n57056), .B(n58662), .Y(n57057) );
  NAND2X1 U60735 ( .A(n57058), .B(n57057), .Y(n58670) );
  NAND2X1 U60736 ( .A(n57059), .B(n58670), .Y(n57060) );
  NAND2X1 U60737 ( .A(n57061), .B(n57060), .Y(n58678) );
  NAND2X1 U60738 ( .A(n57062), .B(n58678), .Y(n57063) );
  NAND2X1 U60739 ( .A(n57064), .B(n57063), .Y(n58686) );
  NAND2X1 U60740 ( .A(n57065), .B(n58686), .Y(n57066) );
  NAND2X1 U60741 ( .A(n57067), .B(n57066), .Y(n58694) );
  NAND2X1 U60742 ( .A(n57068), .B(n58694), .Y(n57069) );
  NAND2X1 U60743 ( .A(n57070), .B(n57069), .Y(n58702) );
  NAND2X1 U60744 ( .A(n57071), .B(n58702), .Y(n57072) );
  NAND2X1 U60745 ( .A(n57073), .B(n57072), .Y(n58710) );
  NAND2X1 U60746 ( .A(n57074), .B(n58710), .Y(n57075) );
  NAND2X1 U60747 ( .A(n57076), .B(n57075), .Y(n58718) );
  NAND2X1 U60748 ( .A(n57077), .B(n58718), .Y(n57078) );
  NAND2X1 U60749 ( .A(n57079), .B(n57078), .Y(n58726) );
  NAND2X1 U60750 ( .A(n57080), .B(n58726), .Y(n57081) );
  NAND2X1 U60751 ( .A(n57082), .B(n57081), .Y(n58735) );
  NAND2X1 U60752 ( .A(n57083), .B(n58735), .Y(n57084) );
  NAND2X1 U60753 ( .A(n57085), .B(n57084), .Y(n58750) );
  NOR2X1 U60754 ( .A(n57086), .B(n58750), .Y(n57088) );
  INVX1 U60755 ( .A(n15810), .Y(n73440) );
  NOR2X1 U60756 ( .A(n15862), .B(n73440), .Y(n57087) );
  INVX1 U60757 ( .A(n57318), .Y(n57319) );
  INVX1 U60758 ( .A(n58544), .Y(n57334) );
  INVX1 U60759 ( .A(n57089), .Y(n57093) );
  NOR2X1 U60760 ( .A(opcode_instr_w_16), .B(n42609), .Y(n57090) );
  NOR2X1 U60761 ( .A(opcode_instr_w_17), .B(n57090), .Y(n57091) );
  NOR2X1 U60762 ( .A(opcode_instr_w[11]), .B(n57091), .Y(n57092) );
  NOR2X1 U60763 ( .A(n57093), .B(n57092), .Y(n57103) );
  NAND2X1 U60764 ( .A(n17896), .B(n57094), .Y(n57101) );
  NAND2X1 U60765 ( .A(opcode_instr_w[8]), .B(n57095), .Y(n57097) );
  NAND2X1 U60766 ( .A(n57097), .B(n57096), .Y(n57098) );
  NAND2X1 U60767 ( .A(n57099), .B(n57098), .Y(n57100) );
  AND2X1 U60768 ( .A(n57101), .B(n57100), .Y(n57102) );
  NAND2X1 U60769 ( .A(n57103), .B(n57102), .Y(n57326) );
  NOR2X1 U60770 ( .A(n57334), .B(n57326), .Y(n57104) );
  NAND2X1 U60771 ( .A(n57104), .B(n58543), .Y(n58802) );
  NOR2X1 U60772 ( .A(n57319), .B(n43436), .Y(n57106) );
  NAND2X1 U60773 ( .A(n15815), .B(n15779), .Y(n57105) );
  NOR2X1 U60774 ( .A(n57106), .B(n57105), .Y(n57110) );
  NOR2X1 U60775 ( .A(n43414), .B(n37340), .Y(n57107) );
  OR2X1 U60776 ( .A(n15813), .B(n57107), .Y(n57108) );
  NOR2X1 U60777 ( .A(n15777), .B(n57108), .Y(n57109) );
  NAND2X1 U60778 ( .A(n57110), .B(n57109), .Y(u_exec_alu_p_w[31]) );
  NOR2X1 U60779 ( .A(n44539), .B(n43281), .Y(n57112) );
  NOR2X1 U60780 ( .A(n44537), .B(n43282), .Y(n57111) );
  NOR2X1 U60781 ( .A(n57112), .B(n57111), .Y(n57114) );
  NOR2X1 U60782 ( .A(n19679), .B(n19676), .Y(n57113) );
  NAND2X1 U60783 ( .A(n57114), .B(n57113), .Y(u_decode_u_regfile_N686) );
  NOR2X1 U60784 ( .A(n19088), .B(n43281), .Y(n57116) );
  NOR2X1 U60785 ( .A(n44564), .B(n43284), .Y(n57115) );
  NOR2X1 U60786 ( .A(n57116), .B(n57115), .Y(n57118) );
  NOR2X1 U60787 ( .A(n19089), .B(n19087), .Y(n57117) );
  NAND2X1 U60788 ( .A(n57118), .B(n57117), .Y(u_decode_u_regfile_N797) );
  NOR2X1 U60789 ( .A(n23541), .B(n43281), .Y(n57120) );
  NOR2X1 U60790 ( .A(n44315), .B(n43284), .Y(n57119) );
  NOR2X1 U60791 ( .A(n57120), .B(n57119), .Y(n57122) );
  NOR2X1 U60792 ( .A(n23542), .B(n23539), .Y(n57121) );
  NAND2X1 U60793 ( .A(n57122), .B(n57121), .Y(u_decode_u_regfile_N1093) );
  NOR2X1 U60794 ( .A(n22229), .B(n43281), .Y(n57124) );
  NOR2X1 U60795 ( .A(n44393), .B(n43284), .Y(n57123) );
  NOR2X1 U60796 ( .A(n57124), .B(n57123), .Y(n57126) );
  NOR2X1 U60797 ( .A(n22230), .B(n22227), .Y(n57125) );
  NAND2X1 U60798 ( .A(n57126), .B(n57125), .Y(u_decode_u_regfile_N205) );
  NOR2X1 U60799 ( .A(n20659), .B(n43281), .Y(n57128) );
  NOR2X1 U60800 ( .A(n44483), .B(n43284), .Y(n57127) );
  NOR2X1 U60801 ( .A(n57128), .B(n57127), .Y(n57130) );
  NOR2X1 U60802 ( .A(n20660), .B(n20657), .Y(n57129) );
  NAND2X1 U60803 ( .A(n57130), .B(n57129), .Y(u_decode_u_regfile_N501) );
  NOR2X1 U60804 ( .A(n43279), .B(n43271), .Y(n57133) );
  NOR2X1 U60805 ( .A(n43282), .B(n43386), .Y(n57132) );
  NOR2X1 U60806 ( .A(n57133), .B(n57132), .Y(n57135) );
  NOR2X1 U60807 ( .A(n21249), .B(n21246), .Y(n57134) );
  NAND2X1 U60808 ( .A(n57135), .B(n57134), .Y(u_decode_u_regfile_N390) );
  NOR2X1 U60809 ( .A(n44603), .B(n43280), .Y(n57137) );
  NOR2X1 U60810 ( .A(n44600), .B(n43283), .Y(n57136) );
  NOR2X1 U60811 ( .A(n57137), .B(n57136), .Y(n57139) );
  NOR2X1 U60812 ( .A(n18089), .B(n18086), .Y(n57138) );
  NAND2X1 U60813 ( .A(n57139), .B(n57138), .Y(u_decode_u_regfile_N982) );
  NOR2X1 U60814 ( .A(n19481), .B(n43280), .Y(n57141) );
  NOR2X1 U60815 ( .A(n44549), .B(n43283), .Y(n57140) );
  NOR2X1 U60816 ( .A(n57141), .B(n57140), .Y(n57143) );
  NOR2X1 U60817 ( .A(n19482), .B(n19479), .Y(n57142) );
  NAND2X1 U60818 ( .A(n57143), .B(n57142), .Y(u_decode_u_regfile_N723) );
  NOR2X1 U60819 ( .A(n43279), .B(n57144), .Y(n57146) );
  NOR2X1 U60820 ( .A(n43282), .B(n43389), .Y(n57145) );
  NOR2X1 U60821 ( .A(n57146), .B(n57145), .Y(n57148) );
  NOR2X1 U60822 ( .A(n22622), .B(n22619), .Y(n57147) );
  NAND2X1 U60823 ( .A(n57148), .B(n57147), .Y(u_decode_u_regfile_N131) );
  NOR2X1 U60824 ( .A(n21051), .B(n43280), .Y(n57150) );
  NOR2X1 U60825 ( .A(n44459), .B(n43283), .Y(n57149) );
  NOR2X1 U60826 ( .A(n57150), .B(n57149), .Y(n57152) );
  NOR2X1 U60827 ( .A(n21052), .B(n21049), .Y(n57151) );
  NAND2X1 U60828 ( .A(n57152), .B(n57151), .Y(u_decode_u_regfile_N427) );
  NOR2X1 U60829 ( .A(n18002), .B(n43280), .Y(n57154) );
  NOR2X1 U60830 ( .A(n44606), .B(n43283), .Y(n57153) );
  NOR2X1 U60831 ( .A(n57154), .B(n57153), .Y(n57156) );
  NOR2X1 U60832 ( .A(n23980), .B(n23979), .Y(n57155) );
  NAND2X1 U60833 ( .A(n57156), .B(n57155), .Y(u_decode_u_regfile_N1019) );
  NOR2X1 U60834 ( .A(n23321), .B(n43280), .Y(n57158) );
  NOR2X1 U60835 ( .A(n44327), .B(n43283), .Y(n57157) );
  NOR2X1 U60836 ( .A(n57158), .B(n57157), .Y(n57160) );
  NOR2X1 U60837 ( .A(n23322), .B(n23319), .Y(n57159) );
  NAND2X1 U60838 ( .A(n57160), .B(n57159), .Y(u_decode_u_regfile_N1130) );
  NOR2X1 U60839 ( .A(n22033), .B(n43280), .Y(n57162) );
  NOR2X1 U60840 ( .A(n44405), .B(n43283), .Y(n57161) );
  NOR2X1 U60841 ( .A(n57162), .B(n57161), .Y(n57164) );
  NOR2X1 U60842 ( .A(n22034), .B(n22031), .Y(n57163) );
  NAND2X1 U60843 ( .A(n57164), .B(n57163), .Y(u_decode_u_regfile_N242) );
  NOR2X1 U60844 ( .A(n18696), .B(n43280), .Y(n57166) );
  NOR2X1 U60845 ( .A(n44576), .B(n43283), .Y(n57165) );
  NOR2X1 U60846 ( .A(n57166), .B(n57165), .Y(n57168) );
  NOR2X1 U60847 ( .A(n18697), .B(n18695), .Y(n57167) );
  NAND2X1 U60848 ( .A(n57168), .B(n57167), .Y(u_decode_u_regfile_N871) );
  NOR2X1 U60849 ( .A(n23761), .B(n43280), .Y(n57170) );
  NOR2X1 U60850 ( .A(n44303), .B(n43283), .Y(n57169) );
  NOR2X1 U60851 ( .A(n57170), .B(n57169), .Y(n57172) );
  NOR2X1 U60852 ( .A(n23762), .B(n23759), .Y(n57171) );
  NAND2X1 U60853 ( .A(n57172), .B(n57171), .Y(u_decode_u_regfile_N1056) );
  NOR2X1 U60854 ( .A(n23107), .B(n43280), .Y(n57174) );
  NOR2X1 U60855 ( .A(n44339), .B(n43283), .Y(n57173) );
  NOR2X1 U60856 ( .A(n57174), .B(n57173), .Y(n57176) );
  NOR2X1 U60857 ( .A(n23108), .B(n23105), .Y(n57175) );
  NAND2X1 U60858 ( .A(n57176), .B(n57175), .Y(u_decode_u_regfile_N1167) );
  NOR2X1 U60859 ( .A(n22425), .B(n43280), .Y(n57178) );
  NOR2X1 U60860 ( .A(n44381), .B(n43283), .Y(n57177) );
  NOR2X1 U60861 ( .A(n57178), .B(n57177), .Y(n57180) );
  NOR2X1 U60862 ( .A(n22426), .B(n22423), .Y(n57179) );
  NAND2X1 U60863 ( .A(n57180), .B(n57179), .Y(u_decode_u_regfile_N168) );
  NOR2X1 U60864 ( .A(n20267), .B(n43280), .Y(n57182) );
  NOR2X1 U60865 ( .A(n44501), .B(n43283), .Y(n57181) );
  NOR2X1 U60866 ( .A(n57182), .B(n57181), .Y(n57184) );
  NOR2X1 U60867 ( .A(n20268), .B(n20265), .Y(n57183) );
  NAND2X1 U60868 ( .A(n57184), .B(n57183), .Y(u_decode_u_regfile_N575) );
  NOR2X1 U60869 ( .A(n21641), .B(n43280), .Y(n57186) );
  NOR2X1 U60870 ( .A(n44429), .B(n43283), .Y(n57185) );
  NOR2X1 U60871 ( .A(n57186), .B(n57185), .Y(n57188) );
  NOR2X1 U60872 ( .A(n21642), .B(n21639), .Y(n57187) );
  NAND2X1 U60873 ( .A(n57188), .B(n57187), .Y(u_decode_u_regfile_N316) );
  NOR2X1 U60874 ( .A(n22887), .B(n43280), .Y(n57190) );
  NOR2X1 U60875 ( .A(n44351), .B(n43283), .Y(n57189) );
  NOR2X1 U60876 ( .A(n57190), .B(n57189), .Y(n57192) );
  NOR2X1 U60877 ( .A(n22888), .B(n22885), .Y(n57191) );
  NAND2X1 U60878 ( .A(n57192), .B(n57191), .Y(u_decode_u_regfile_N1204) );
  NOR2X1 U60879 ( .A(n44573), .B(n43279), .Y(n57194) );
  NOR2X1 U60880 ( .A(n44570), .B(n43282), .Y(n57193) );
  NOR2X1 U60881 ( .A(n57194), .B(n57193), .Y(n57196) );
  NOR2X1 U60882 ( .A(n18893), .B(n18891), .Y(n57195) );
  NAND2X1 U60883 ( .A(n57196), .B(n57195), .Y(u_decode_u_regfile_N834) );
  NOR2X1 U60884 ( .A(n44474), .B(n43279), .Y(n57198) );
  NOR2X1 U60885 ( .A(n44471), .B(n43282), .Y(n57197) );
  NOR2X1 U60886 ( .A(n57198), .B(n57197), .Y(n57200) );
  NOR2X1 U60887 ( .A(n20856), .B(n20853), .Y(n57199) );
  NAND2X1 U60888 ( .A(n57200), .B(n57199), .Y(u_decode_u_regfile_N464) );
  NOR2X1 U60889 ( .A(n19875), .B(n43279), .Y(n57202) );
  NOR2X1 U60890 ( .A(n44525), .B(n43282), .Y(n57201) );
  NOR2X1 U60891 ( .A(n57202), .B(n57201), .Y(n57204) );
  NOR2X1 U60892 ( .A(n19876), .B(n19873), .Y(n57203) );
  NAND2X1 U60893 ( .A(n57204), .B(n57203), .Y(u_decode_u_regfile_N649) );
  NOR2X1 U60894 ( .A(n20071), .B(n43279), .Y(n57206) );
  NOR2X1 U60895 ( .A(n44513), .B(n43282), .Y(n57205) );
  NOR2X1 U60896 ( .A(n57206), .B(n57205), .Y(n57208) );
  NOR2X1 U60897 ( .A(n20072), .B(n20069), .Y(n57207) );
  NAND2X1 U60898 ( .A(n57208), .B(n57207), .Y(u_decode_u_regfile_N612) );
  NOR2X1 U60899 ( .A(n43279), .B(n57209), .Y(n57211) );
  NOR2X1 U60900 ( .A(n43282), .B(n43383), .Y(n57210) );
  NOR2X1 U60901 ( .A(n57211), .B(n57210), .Y(n57213) );
  NOR2X1 U60902 ( .A(n20464), .B(n20461), .Y(n57212) );
  NAND2X1 U60903 ( .A(n57213), .B(n57212), .Y(u_decode_u_regfile_N538) );
  NOR2X1 U60904 ( .A(n21837), .B(n43279), .Y(n57215) );
  NOR2X1 U60905 ( .A(n44417), .B(n43282), .Y(n57214) );
  NOR2X1 U60906 ( .A(n57215), .B(n57214), .Y(n57217) );
  NOR2X1 U60907 ( .A(n21838), .B(n21835), .Y(n57216) );
  NAND2X1 U60908 ( .A(n57217), .B(n57216), .Y(u_decode_u_regfile_N279) );
  NOR2X1 U60909 ( .A(n18305), .B(n43279), .Y(n57219) );
  NOR2X1 U60910 ( .A(n44591), .B(n43282), .Y(n57218) );
  NOR2X1 U60911 ( .A(n57219), .B(n57218), .Y(n57221) );
  NOR2X1 U60912 ( .A(n18306), .B(n18303), .Y(n57220) );
  NAND2X1 U60913 ( .A(n57221), .B(n57220), .Y(u_decode_u_regfile_N945) );
  NOR2X1 U60914 ( .A(n44585), .B(n43279), .Y(n57223) );
  NOR2X1 U60915 ( .A(n44582), .B(n43282), .Y(n57222) );
  NOR2X1 U60916 ( .A(n57223), .B(n57222), .Y(n57225) );
  NOR2X1 U60917 ( .A(n18501), .B(n18499), .Y(n57224) );
  NAND2X1 U60918 ( .A(n57225), .B(n57224), .Y(u_decode_u_regfile_N908) );
  NOR2X1 U60919 ( .A(n44561), .B(n43279), .Y(n57227) );
  NOR2X1 U60920 ( .A(n44558), .B(n43282), .Y(n57226) );
  NOR2X1 U60921 ( .A(n57227), .B(n57226), .Y(n57229) );
  NOR2X1 U60922 ( .A(n19285), .B(n19283), .Y(n57228) );
  NAND2X1 U60923 ( .A(n57229), .B(n57228), .Y(u_decode_u_regfile_N760) );
  NOR2X1 U60924 ( .A(n21445), .B(n43279), .Y(n57231) );
  NOR2X1 U60925 ( .A(n44441), .B(n43282), .Y(n57230) );
  NOR2X1 U60926 ( .A(n57231), .B(n57230), .Y(n57233) );
  NOR2X1 U60927 ( .A(n21446), .B(n21443), .Y(n57232) );
  NAND2X1 U60928 ( .A(n57233), .B(n57232), .Y(u_decode_u_regfile_N353) );
  NOR2X1 U60929 ( .A(n22667), .B(n43280), .Y(n57236) );
  NOR2X1 U60930 ( .A(n44363), .B(n43283), .Y(n57235) );
  NOR2X1 U60931 ( .A(n57236), .B(n57235), .Y(n57238) );
  NOR2X1 U60932 ( .A(n22668), .B(n22665), .Y(n57237) );
  NAND2X1 U60933 ( .A(n57238), .B(n57237), .Y(u_decode_u_regfile_N1241) );
  NOR2X1 U60934 ( .A(n57563), .B(n57405), .Y(u_decode_N761) );
  NOR2X1 U60935 ( .A(n57563), .B(n57414), .Y(u_decode_N760) );
  NAND2X1 U60936 ( .A(n43013), .B(n42873), .Y(n57239) );
  NAND2X1 U60937 ( .A(u_csr_N184), .B(n57239), .Y(n57255) );
  NOR2X1 U60938 ( .A(n57255), .B(n57240), .Y(n57246) );
  NAND2X1 U60939 ( .A(u_csr_N184), .B(n57241), .Y(n57244) );
  NAND2X1 U60940 ( .A(n27560), .B(n26906), .Y(n57242) );
  NAND2X1 U60941 ( .A(u_csr_csr_mepc_q[0]), .B(n57242), .Y(n57243) );
  NAND2X1 U60942 ( .A(n57244), .B(n57243), .Y(n57245) );
  NOR2X1 U60943 ( .A(n57246), .B(n57245), .Y(n57253) );
  NOR2X1 U60944 ( .A(n42952), .B(n37747), .Y(n57251) );
  INVX1 U60945 ( .A(n26127), .Y(n73521) );
  NAND2X1 U60946 ( .A(n73521), .B(n42442), .Y(n58277) );
  INVX1 U60947 ( .A(n58277), .Y(n58451) );
  NAND2X1 U60948 ( .A(n58451), .B(n57247), .Y(n57249) );
  NAND2X1 U60949 ( .A(n43288), .B(n57273), .Y(n57248) );
  NAND2X1 U60950 ( .A(n57249), .B(n57248), .Y(n57250) );
  NOR2X1 U60951 ( .A(n57251), .B(n57250), .Y(n57252) );
  NAND2X1 U60952 ( .A(n57253), .B(n57252), .Y(u_csr_csr_mepc_r[0]) );
  NOR2X1 U60953 ( .A(n8848), .B(n57254), .Y(n57260) );
  INVX1 U60954 ( .A(n57255), .Y(n57274) );
  NAND2X1 U60955 ( .A(n43291), .B(n57274), .Y(n57258) );
  NAND2X1 U60956 ( .A(u_csr_N184), .B(n57256), .Y(n57257) );
  NAND2X1 U60957 ( .A(n57258), .B(n57257), .Y(n57259) );
  NOR2X1 U60958 ( .A(n57260), .B(n57259), .Y(n57266) );
  NOR2X1 U60959 ( .A(n58274), .B(n58277), .Y(n57262) );
  NOR2X1 U60960 ( .A(n42957), .B(n37747), .Y(n57261) );
  NOR2X1 U60961 ( .A(n57262), .B(n57261), .Y(n57264) );
  NAND2X1 U60962 ( .A(n26905), .B(u_csr_csr_sepc_q[0]), .Y(n57263) );
  AND2X1 U60963 ( .A(n57264), .B(n57263), .Y(n57265) );
  NAND2X1 U60964 ( .A(n57266), .B(n57265), .Y(u_csr_csr_sepc_r[0]) );
  AND2X1 U60965 ( .A(n28512), .B(n28508), .Y(n57270) );
  NOR2X1 U60966 ( .A(n58456), .B(n43293), .Y(n57268) );
  NOR2X1 U60967 ( .A(n58455), .B(n43296), .Y(n57267) );
  NOR2X1 U60968 ( .A(n57268), .B(n57267), .Y(n57269) );
  NAND2X1 U60969 ( .A(n57270), .B(n57269), .Y(u_csr_N3665) );
  NAND2X1 U60970 ( .A(n43300), .B(n57274), .Y(n57272) );
  NAND2X1 U60971 ( .A(n43303), .B(n57273), .Y(n57271) );
  NAND2X1 U60972 ( .A(n57272), .B(n57271), .Y(net2281) );
  NOR2X1 U60973 ( .A(n1940), .B(n43306), .Y(n57277) );
  NAND2X1 U60974 ( .A(n43308), .B(n57273), .Y(n57276) );
  NAND2X1 U60975 ( .A(n57274), .B(n43313), .Y(n57275) );
  NAND2X1 U60976 ( .A(n57276), .B(n57275), .Y(n57281) );
  NOR2X1 U60977 ( .A(n57277), .B(n57281), .Y(n57279) );
  OR2X1 U60978 ( .A(n1758), .B(n42847), .Y(n57278) );
  NAND2X1 U60979 ( .A(n57279), .B(n57278), .Y(mem_i_pc_o[0]) );
  NOR2X1 U60980 ( .A(n43315), .B(n57283), .Y(net2380) );
  NOR2X1 U60981 ( .A(n1941), .B(n43322), .Y(n57282) );
  NOR2X1 U60982 ( .A(n57282), .B(n57281), .Y(n57288) );
  NOR2X1 U60983 ( .A(n43325), .B(n57283), .Y(n57286) );
  NOR2X1 U60984 ( .A(n57284), .B(n43328), .Y(n57285) );
  NOR2X1 U60985 ( .A(n57286), .B(n57285), .Y(n57287) );
  NAND2X1 U60986 ( .A(n57288), .B(n57287), .Y(u_decode_N290) );
  NAND2X1 U60987 ( .A(n58597), .B(n42942), .Y(n57289) );
  NAND2X1 U60988 ( .A(n15945), .B(n57289), .Y(n57290) );
  NOR2X1 U60989 ( .A(n15948), .B(n57290), .Y(n57293) );
  OR2X1 U60990 ( .A(n15896), .B(n15938), .Y(n57291) );
  NOR2X1 U60991 ( .A(n15897), .B(n57291), .Y(n57292) );
  NAND2X1 U60992 ( .A(n57293), .B(n57292), .Y(u_exec_alu_p_w[2]) );
  NOR2X1 U60993 ( .A(n22667), .B(n43330), .Y(n57295) );
  NOR2X1 U60994 ( .A(n44363), .B(n43333), .Y(n57294) );
  NOR2X1 U60995 ( .A(n57295), .B(n57294), .Y(n57297) );
  NOR2X1 U60996 ( .A(n22862), .B(n22861), .Y(n57296) );
  NAND2X1 U60997 ( .A(n57297), .B(n57296), .Y(u_decode_u_regfile_N1212) );
  NAND2X1 U60998 ( .A(n15682), .B(n15734), .Y(n15737) );
  NOR2X1 U60999 ( .A(n15465), .B(n43422), .Y(n57298) );
  OR2X1 U61000 ( .A(n15749), .B(n57298), .Y(n361) );
  INVX1 U61001 ( .A(n15505), .Y(n73570) );
  NAND2X1 U61002 ( .A(n42948), .B(n73570), .Y(n15722) );
  NAND2X1 U61003 ( .A(n43419), .B(n73570), .Y(n15747) );
  NAND2X1 U61004 ( .A(n42451), .B(n73570), .Y(n15723) );
  NAND2X1 U61005 ( .A(n43424), .B(n73570), .Y(n15649) );
  INVX1 U61006 ( .A(n15723), .Y(n57299) );
  NAND2X1 U61007 ( .A(n15443), .B(n57299), .Y(n57302) );
  INVX1 U61008 ( .A(n15747), .Y(n57300) );
  NAND2X1 U61009 ( .A(n15441), .B(n57300), .Y(n57301) );
  NAND2X1 U61010 ( .A(n57302), .B(n57301), .Y(n57307) );
  INVX1 U61011 ( .A(n15722), .Y(n57303) );
  NAND2X1 U61012 ( .A(n17094), .B(n57303), .Y(n57305) );
  NAND2X1 U61013 ( .A(n58597), .B(n42972), .Y(n57304) );
  NAND2X1 U61014 ( .A(n57305), .B(n57304), .Y(n57306) );
  NOR2X1 U61015 ( .A(n57307), .B(n57306), .Y(n57311) );
  NOR2X1 U61016 ( .A(n15649), .B(n73490), .Y(n57308) );
  OR2X1 U61017 ( .A(n17883), .B(n57308), .Y(n57309) );
  NOR2X1 U61018 ( .A(n17425), .B(n57309), .Y(n57310) );
  NAND2X1 U61019 ( .A(n57311), .B(n57310), .Y(n57345) );
  INVX1 U61020 ( .A(n15495), .Y(n57312) );
  NAND2X1 U61021 ( .A(n15736), .B(n57312), .Y(n57313) );
  NAND2X1 U61022 ( .A(n17880), .B(n57313), .Y(n57315) );
  NAND2X1 U61023 ( .A(n17808), .B(n17809), .Y(n57314) );
  NOR2X1 U61024 ( .A(n57315), .B(n57314), .Y(n57343) );
  NAND2X1 U61025 ( .A(n58597), .B(n57316), .Y(n58658) );
  NOR2X1 U61026 ( .A(n42968), .B(n58658), .Y(n57341) );
  INVX1 U61027 ( .A(n57333), .Y(n57317) );
  NOR2X1 U61028 ( .A(n57334), .B(n57317), .Y(n57330) );
  NAND2X1 U61029 ( .A(n73437), .B(n57318), .Y(n57322) );
  NAND2X1 U61030 ( .A(n57319), .B(n57323), .Y(n57320) );
  NAND2X1 U61031 ( .A(n57320), .B(n58580), .Y(n57321) );
  NAND2X1 U61032 ( .A(n57322), .B(n57321), .Y(n57328) );
  NAND2X1 U61033 ( .A(n17446), .B(n73438), .Y(n57325) );
  NAND2X1 U61034 ( .A(n17444), .B(n57323), .Y(n57324) );
  NAND2X1 U61035 ( .A(n57325), .B(n57324), .Y(n57327) );
  INVX1 U61036 ( .A(n57326), .Y(n73513) );
  MX2X1 U61037 ( .A(n57328), .B(n57327), .S0(n73513), .Y(n57329) );
  NAND2X1 U61038 ( .A(n57330), .B(n57329), .Y(n57339) );
  NAND2X1 U61039 ( .A(n57331), .B(n58597), .Y(n57332) );
  NAND2X1 U61040 ( .A(n57332), .B(n58659), .Y(n57337) );
  NAND2X1 U61041 ( .A(n57334), .B(n58543), .Y(n58805) );
  INVX1 U61042 ( .A(n58805), .Y(n58801) );
  NOR2X1 U61043 ( .A(n43427), .B(n43434), .Y(n57335) );
  NAND2X1 U61044 ( .A(n57334), .B(n57333), .Y(n58759) );
  NAND2X1 U61045 ( .A(n57335), .B(n58759), .Y(n57336) );
  NAND2X1 U61046 ( .A(n57337), .B(n57336), .Y(n57338) );
  NAND2X1 U61047 ( .A(n57339), .B(n57338), .Y(n57340) );
  NOR2X1 U61048 ( .A(n57341), .B(n57340), .Y(n57342) );
  NAND2X1 U61049 ( .A(n57343), .B(n57342), .Y(n57344) );
  OR2X1 U61050 ( .A(n57345), .B(n57344), .Y(u_exec_alu_p_w[0]) );
  NOR2X1 U61051 ( .A(n18002), .B(n43451), .Y(n57347) );
  NOR2X1 U61052 ( .A(n44606), .B(n43336), .Y(n57346) );
  NOR2X1 U61053 ( .A(n57347), .B(n57346), .Y(n57349) );
  NOR2X1 U61054 ( .A(n18081), .B(n18079), .Y(n57348) );
  NAND2X1 U61055 ( .A(n57349), .B(n57348), .Y(u_decode_u_regfile_N988) );
  INVX1 U61056 ( .A(n57350), .Y(n57352) );
  NAND2X1 U61057 ( .A(n57352), .B(n42608), .Y(n57357) );
  NOR2X1 U61058 ( .A(n57353), .B(n57362), .Y(n57356) );
  NAND2X1 U61059 ( .A(opcode_instr_w_36), .B(n57365), .Y(n57354) );
  NAND2X1 U61060 ( .A(n57354), .B(n58812), .Y(n57355) );
  NAND2X1 U61061 ( .A(n57356), .B(n57355), .Y(n72740) );
  NAND2X1 U61062 ( .A(n57357), .B(n72740), .Y(u_lsu_N226) );
  NOR2X1 U61063 ( .A(n73430), .B(n57364), .Y(n57358) );
  NAND2X1 U61064 ( .A(n42608), .B(n57358), .Y(n72739) );
  NAND2X1 U61065 ( .A(n72739), .B(n72740), .Y(u_lsu_N227) );
  NOR2X1 U61066 ( .A(n73431), .B(n57362), .Y(n57359) );
  NAND2X1 U61067 ( .A(opcode_instr_w_36), .B(n57560), .Y(n57367) );
  NAND2X1 U61068 ( .A(n57367), .B(n57360), .Y(n57361) );
  NAND2X1 U61069 ( .A(n42318), .B(n57361), .Y(n72756) );
  NOR2X1 U61070 ( .A(n57362), .B(n58812), .Y(n57363) );
  NAND2X1 U61071 ( .A(n57363), .B(n57560), .Y(n72796) );
  NAND2X1 U61072 ( .A(n72756), .B(n72796), .Y(u_lsu_N228) );
  NOR2X1 U61073 ( .A(n57365), .B(n57364), .Y(n57366) );
  NAND2X1 U61074 ( .A(n57366), .B(n42608), .Y(n72736) );
  INVX1 U61075 ( .A(n72796), .Y(n72816) );
  INVX1 U61076 ( .A(n57367), .Y(n57368) );
  NAND2X1 U61077 ( .A(n57368), .B(n42318), .Y(n72797) );
  INVX1 U61078 ( .A(n72797), .Y(n57369) );
  NOR2X1 U61079 ( .A(n72816), .B(n57369), .Y(n57370) );
  NAND2X1 U61080 ( .A(n72736), .B(n57370), .Y(u_lsu_N229) );
  NAND2X1 U61081 ( .A(n42441), .B(n58194), .Y(n57372) );
  NAND2X1 U61082 ( .A(u_mmu_store_q[0]), .B(n57377), .Y(n57371) );
  NAND2X1 U61083 ( .A(n57372), .B(n57371), .Y(n8542) );
  NAND2X1 U61084 ( .A(n42441), .B(n37328), .Y(n57374) );
  NAND2X1 U61085 ( .A(u_mmu_store_q[1]), .B(n57377), .Y(n57373) );
  NAND2X1 U61086 ( .A(n57374), .B(n57373), .Y(n8541) );
  NAND2X1 U61087 ( .A(n42441), .B(n37327), .Y(n57376) );
  NAND2X1 U61088 ( .A(u_mmu_store_q[2]), .B(n57377), .Y(n57375) );
  NAND2X1 U61089 ( .A(n57376), .B(n57375), .Y(n8540) );
  NAND2X1 U61090 ( .A(n42441), .B(n58184), .Y(n57379) );
  NAND2X1 U61091 ( .A(u_mmu_store_q[3]), .B(n57377), .Y(n57378) );
  NAND2X1 U61092 ( .A(n57379), .B(n57378), .Y(n8539) );
  NOR2X1 U61093 ( .A(n28797), .B(n43380), .Y(n57383) );
  INVX1 U61094 ( .A(n28765), .Y(n57916) );
  NOR2X1 U61095 ( .A(n57380), .B(n57916), .Y(n57381) );
  NAND2X1 U61096 ( .A(n57381), .B(n37550), .Y(n57382) );
  NAND2X1 U61097 ( .A(n57383), .B(n57382), .Y(n8555) );
  NAND2X1 U61098 ( .A(u_mmu_dtlb_req_q), .B(n37547), .Y(n28953) );
  INVX1 U61099 ( .A(n28953), .Y(n73429) );
  NOR2X1 U61100 ( .A(u_mmu_dtlb_valid_q), .B(n73429), .Y(n57384) );
  NOR2X1 U61101 ( .A(n57385), .B(n57384), .Y(n8504) );
  MX2X1 U61102 ( .A(u_mmu_dtlb_va_addr_q[24]), .B(n57386), .S0(n73429), .Y(
        n8428) );
  MX2X1 U61103 ( .A(u_mmu_dtlb_va_addr_q[30]), .B(u_mmu_virt_addr_q_30), .S0(
        n73429), .Y(n8426) );
  MX2X1 U61104 ( .A(u_mmu_dtlb_va_addr_q[28]), .B(u_mmu_virt_addr_q_28), .S0(
        n73429), .Y(n8439) );
  MX2X1 U61105 ( .A(u_mmu_dtlb_va_addr_q[23]), .B(n57387), .S0(n73429), .Y(
        n8437) );
  MX2X1 U61106 ( .A(u_mmu_dtlb_va_addr_q[22]), .B(n57388), .S0(n73429), .Y(
        n8435) );
  MX2X1 U61107 ( .A(u_mmu_dtlb_va_addr_q[21]), .B(u_mmu_virt_addr_q[21]), .S0(
        n73429), .Y(n8434) );
  MX2X1 U61108 ( .A(u_mmu_dtlb_va_addr_q[26]), .B(n57389), .S0(n73429), .Y(
        n8432) );
  MX2X1 U61109 ( .A(u_mmu_dtlb_va_addr_q[27]), .B(n57390), .S0(n73429), .Y(
        n8445) );
  NAND2X1 U61110 ( .A(n73429), .B(n57391), .Y(n57392) );
  NAND2X1 U61111 ( .A(n28982), .B(n57392), .Y(n8430) );
  MX2X1 U61112 ( .A(u_mmu_dtlb_va_addr_q[31]), .B(u_mmu_virt_addr_q_31), .S0(
        n73429), .Y(n8424) );
  NAND2X1 U61113 ( .A(u_mmu_virt_addr_q_29), .B(n73429), .Y(n57393) );
  NAND2X1 U61114 ( .A(n28996), .B(n57393), .Y(n8423) );
  INVX1 U61115 ( .A(n57394), .Y(n57396) );
  NAND2X1 U61116 ( .A(n57396), .B(n57395), .Y(n57899) );
  NAND2X1 U61117 ( .A(n57899), .B(n57397), .Y(n57960) );
  NAND2X1 U61118 ( .A(mem_d_accept_i), .B(n44257), .Y(n57398) );
  INVX1 U61119 ( .A(n24488), .Y(n57399) );
  NOR2X1 U61120 ( .A(n24384), .B(n57399), .Y(n57403) );
  NOR2X1 U61121 ( .A(n57401), .B(n57400), .Y(n57402) );
  NAND2X1 U61122 ( .A(n57403), .B(n57402), .Y(n24406) );
  NOR2X1 U61123 ( .A(n24406), .B(n57404), .Y(u_decode_N789) );
  NOR2X1 U61124 ( .A(n24406), .B(n57405), .Y(u_decode_N787) );
  NOR2X1 U61125 ( .A(n24406), .B(n57406), .Y(u_decode_N790) );
  NOR2X1 U61126 ( .A(n24406), .B(n57407), .Y(u_decode_N788) );
  NOR2X1 U61127 ( .A(n1891), .B(n58822), .Y(n57408) );
  NAND2X1 U61128 ( .A(n57408), .B(n58165), .Y(n57409) );
  NAND2X1 U61129 ( .A(n42439), .B(n57409), .Y(n28813) );
  NOR2X1 U61130 ( .A(n24406), .B(n58129), .Y(u_decode_N786) );
  INVX1 U61131 ( .A(n24406), .Y(n57410) );
  NAND2X1 U61132 ( .A(n57411), .B(n57410), .Y(n57412) );
  NOR2X1 U61133 ( .A(n57413), .B(n57412), .Y(u_decode_N785) );
  NOR2X1 U61134 ( .A(n24406), .B(n57414), .Y(u_decode_N784) );
  NOR2X1 U61135 ( .A(n24406), .B(n57415), .Y(u_decode_N783) );
  INVX1 U61136 ( .A(n57416), .Y(n57421) );
  NOR2X1 U61137 ( .A(opcode_opcode_w[9]), .B(n57429), .Y(n57418) );
  NAND2X1 U61138 ( .A(n61174), .B(n57417), .Y(n59119) );
  OR2X1 U61139 ( .A(n1837), .B(n72732), .Y(n57628) );
  NAND2X1 U61140 ( .A(n42439), .B(n57628), .Y(n57547) );
  NAND2X1 U61141 ( .A(n57547), .B(n28813), .Y(n73374) );
  NAND2X1 U61142 ( .A(n57418), .B(n58521), .Y(n57520) );
  NOR2X1 U61143 ( .A(n57419), .B(n57520), .Y(n57420) );
  NOR2X1 U61144 ( .A(n57421), .B(n57420), .Y(n57422) );
  NOR2X1 U61145 ( .A(n24164), .B(n57422), .Y(u_decode_scoreboard_r[3]) );
  INVX1 U61146 ( .A(n57423), .Y(n57425) );
  NOR2X1 U61147 ( .A(n58525), .B(n57520), .Y(n57424) );
  NOR2X1 U61148 ( .A(n57425), .B(n57424), .Y(n57426) );
  NOR2X1 U61149 ( .A(n24278), .B(n57426), .Y(u_decode_scoreboard_r[19]) );
  NOR2X1 U61150 ( .A(n27326), .B(n57427), .Y(u_csr_N3471) );
  NOR2X1 U61151 ( .A(u_csr_writeback_idx_q[3]), .B(n37592), .Y(n57428) );
  NAND2X1 U61152 ( .A(n37332), .B(n37589), .Y(n58518) );
  NAND2X1 U61153 ( .A(n57428), .B(n58518), .Y(n58520) );
  NOR2X1 U61154 ( .A(n24136), .B(n58520), .Y(n57435) );
  NOR2X1 U61155 ( .A(n57429), .B(n57436), .Y(n57430) );
  NAND2X1 U61156 ( .A(n42460), .B(n57438), .Y(n57432) );
  NAND2X1 U61157 ( .A(n57432), .B(n57431), .Y(n57433) );
  NAND2X1 U61158 ( .A(n24243), .B(n57433), .Y(n57434) );
  NOR2X1 U61159 ( .A(n57435), .B(n57434), .Y(u_decode_scoreboard_r[23]) );
  NOR2X1 U61160 ( .A(n24154), .B(n58520), .Y(n57443) );
  NOR2X1 U61161 ( .A(opcode_opcode_w[8]), .B(n57436), .Y(n57437) );
  NAND2X1 U61162 ( .A(n42606), .B(n57438), .Y(n57440) );
  NAND2X1 U61163 ( .A(n57440), .B(n57439), .Y(n57441) );
  NAND2X1 U61164 ( .A(n24260), .B(n57441), .Y(n57442) );
  NOR2X1 U61165 ( .A(n57443), .B(n57442), .Y(u_decode_scoreboard_r[21]) );
  NOR2X1 U61166 ( .A(n37351), .B(n37592), .Y(n57444) );
  NAND2X1 U61167 ( .A(n57444), .B(n58518), .Y(n24180) );
  NOR2X1 U61168 ( .A(n24145), .B(n24180), .Y(n57449) );
  NAND2X1 U61169 ( .A(u_decode_scoreboard_q[30]), .B(n24188), .Y(n57446) );
  NAND2X1 U61170 ( .A(n42460), .B(n57493), .Y(n57445) );
  NAND2X1 U61171 ( .A(n57446), .B(n57445), .Y(n57447) );
  NAND2X1 U61172 ( .A(n24184), .B(n57447), .Y(n57448) );
  NOR2X1 U61173 ( .A(n57449), .B(n57448), .Y(u_decode_scoreboard_r[30]) );
  NOR2X1 U61174 ( .A(u_csr_writeback_idx_q[4]), .B(n37351), .Y(n57450) );
  NAND2X1 U61175 ( .A(n57450), .B(n58518), .Y(n58519) );
  NOR2X1 U61176 ( .A(n24162), .B(n58519), .Y(n57455) );
  NAND2X1 U61177 ( .A(n42606), .B(n57456), .Y(n57452) );
  NAND2X1 U61178 ( .A(n57452), .B(n57451), .Y(n57453) );
  NAND2X1 U61179 ( .A(n24341), .B(n57453), .Y(n57454) );
  NOR2X1 U61180 ( .A(n57455), .B(n57454), .Y(u_decode_scoreboard_r[12]) );
  NOR2X1 U61181 ( .A(n24145), .B(n58519), .Y(n57461) );
  NAND2X1 U61182 ( .A(n42460), .B(n57456), .Y(n57458) );
  NAND2X1 U61183 ( .A(n57458), .B(n57457), .Y(n57459) );
  NAND2X1 U61184 ( .A(n24323), .B(n57459), .Y(n57460) );
  NOR2X1 U61185 ( .A(n57461), .B(n57460), .Y(u_decode_scoreboard_r[14]) );
  NOR2X1 U61186 ( .A(n24136), .B(n58519), .Y(n57466) );
  NAND2X1 U61187 ( .A(n42460), .B(n57472), .Y(n57463) );
  NAND2X1 U61188 ( .A(n57463), .B(n57462), .Y(n57464) );
  NAND2X1 U61189 ( .A(n24312), .B(n57464), .Y(n57465) );
  NOR2X1 U61190 ( .A(n57466), .B(n57465), .Y(u_decode_scoreboard_r[15]) );
  NOR2X1 U61191 ( .A(n24154), .B(n24180), .Y(n57471) );
  NAND2X1 U61192 ( .A(n42606), .B(n58531), .Y(n57468) );
  NAND2X1 U61193 ( .A(n57468), .B(n57467), .Y(n57469) );
  NAND2X1 U61194 ( .A(n24200), .B(n57469), .Y(n57470) );
  NOR2X1 U61195 ( .A(n57471), .B(n57470), .Y(u_decode_scoreboard_r[29]) );
  NOR2X1 U61196 ( .A(n24154), .B(n58519), .Y(n57477) );
  NAND2X1 U61197 ( .A(n42606), .B(n57472), .Y(n57474) );
  NAND2X1 U61198 ( .A(n57474), .B(n57473), .Y(n57475) );
  NAND2X1 U61199 ( .A(n24333), .B(n57475), .Y(n57476) );
  NOR2X1 U61200 ( .A(n57477), .B(n57476), .Y(u_decode_scoreboard_r[13]) );
  INVX1 U61201 ( .A(n57478), .Y(n57481) );
  NOR2X1 U61202 ( .A(n57479), .B(n57520), .Y(n57480) );
  NOR2X1 U61203 ( .A(n57481), .B(n57480), .Y(n57482) );
  NOR2X1 U61204 ( .A(n24212), .B(n57482), .Y(u_decode_scoreboard_r[27]) );
  NAND2X1 U61205 ( .A(n73526), .B(n40841), .Y(n24153) );
  NAND2X1 U61206 ( .A(n37351), .B(n37592), .Y(n24135) );
  NOR2X1 U61207 ( .A(n24154), .B(n24135), .Y(n57487) );
  NAND2X1 U61208 ( .A(u_decode_scoreboard_q[5]), .B(n24153), .Y(n57484) );
  NAND2X1 U61209 ( .A(n42606), .B(n58527), .Y(n57483) );
  NAND2X1 U61210 ( .A(n57484), .B(n57483), .Y(n57485) );
  NAND2X1 U61211 ( .A(n24149), .B(n57485), .Y(n57486) );
  NOR2X1 U61212 ( .A(n57487), .B(n57486), .Y(u_decode_scoreboard_r[5]) );
  NAND2X1 U61213 ( .A(n73526), .B(n57534), .Y(n24161) );
  NOR2X1 U61214 ( .A(n24162), .B(n24135), .Y(n57492) );
  NAND2X1 U61215 ( .A(u_decode_scoreboard_q[4]), .B(n24161), .Y(n57489) );
  NAND2X1 U61216 ( .A(n42606), .B(n57535), .Y(n57488) );
  NAND2X1 U61217 ( .A(n57489), .B(n57488), .Y(n57490) );
  NAND2X1 U61218 ( .A(n24158), .B(n57490), .Y(n57491) );
  NOR2X1 U61219 ( .A(n57492), .B(n57491), .Y(u_decode_scoreboard_r[4]) );
  NAND2X1 U61220 ( .A(n73526), .B(n36009), .Y(n24210) );
  NOR2X1 U61221 ( .A(n24162), .B(n24180), .Y(n57498) );
  NAND2X1 U61222 ( .A(u_decode_scoreboard_q[28]), .B(n24210), .Y(n57495) );
  NAND2X1 U61223 ( .A(n42606), .B(n57493), .Y(n57494) );
  NAND2X1 U61224 ( .A(n57495), .B(n57494), .Y(n57496) );
  NAND2X1 U61225 ( .A(n24207), .B(n57496), .Y(n57497) );
  NOR2X1 U61226 ( .A(n57498), .B(n57497), .Y(u_decode_scoreboard_r[28]) );
  INVX1 U61227 ( .A(n57499), .Y(n73421) );
  NAND2X1 U61228 ( .A(n73421), .B(n73526), .Y(n24270) );
  NOR2X1 U61229 ( .A(n24162), .B(n58520), .Y(n57504) );
  NAND2X1 U61230 ( .A(u_decode_scoreboard_q[20]), .B(n24270), .Y(n57501) );
  NAND2X1 U61231 ( .A(n42606), .B(n57541), .Y(n57500) );
  NAND2X1 U61232 ( .A(n57501), .B(n57500), .Y(n57502) );
  NAND2X1 U61233 ( .A(n24267), .B(n57502), .Y(n57503) );
  NOR2X1 U61234 ( .A(n57504), .B(n57503), .Y(u_decode_scoreboard_r[20]) );
  NOR2X1 U61235 ( .A(n57505), .B(n57520), .Y(n57507) );
  INVX1 U61236 ( .A(n24196), .Y(n525) );
  NOR2X1 U61237 ( .A(n525), .B(n37752), .Y(n57506) );
  NOR2X1 U61238 ( .A(n57507), .B(n57506), .Y(n57508) );
  NOR2X1 U61239 ( .A(n24190), .B(n57508), .Y(u_decode_scoreboard_r[2]) );
  NAND2X1 U61240 ( .A(n36009), .B(n57519), .Y(n24224) );
  NOR2X1 U61241 ( .A(n58529), .B(n57520), .Y(n57510) );
  INVX1 U61242 ( .A(n24224), .Y(n543) );
  NOR2X1 U61243 ( .A(n543), .B(n37753), .Y(n57509) );
  NOR2X1 U61244 ( .A(n57510), .B(n57509), .Y(n57511) );
  NOR2X1 U61245 ( .A(n24219), .B(n57511), .Y(u_decode_scoreboard_r[26]) );
  NAND2X1 U61246 ( .A(n40937), .B(n57519), .Y(n24353) );
  NOR2X1 U61247 ( .A(n58537), .B(n57520), .Y(n57513) );
  INVX1 U61248 ( .A(n24353), .Y(n493) );
  NOR2X1 U61249 ( .A(n493), .B(n37754), .Y(n57512) );
  NOR2X1 U61250 ( .A(n57513), .B(n57512), .Y(n57514) );
  NOR2X1 U61251 ( .A(n24347), .B(n57514), .Y(u_decode_scoreboard_r[11]) );
  NAND2X1 U61252 ( .A(n57515), .B(n57519), .Y(n24361) );
  NOR2X1 U61253 ( .A(n58534), .B(n57520), .Y(n57517) );
  INVX1 U61254 ( .A(n24361), .Y(n501) );
  NOR2X1 U61255 ( .A(n501), .B(n37755), .Y(n57516) );
  NOR2X1 U61256 ( .A(n57517), .B(n57516), .Y(n57518) );
  NOR2X1 U61257 ( .A(n24355), .B(n57518), .Y(u_decode_scoreboard_r[10]) );
  NAND2X1 U61258 ( .A(n73421), .B(n57519), .Y(n24290) );
  NOR2X1 U61259 ( .A(n58523), .B(n57520), .Y(n57522) );
  INVX1 U61260 ( .A(n24290), .Y(n539) );
  NOR2X1 U61261 ( .A(n539), .B(n37756), .Y(n57521) );
  NOR2X1 U61262 ( .A(n57522), .B(n57521), .Y(n57523) );
  NOR2X1 U61263 ( .A(n24285), .B(n57523), .Y(u_decode_scoreboard_r[18]) );
  NOR2X1 U61264 ( .A(n24136), .B(n24135), .Y(n57528) );
  NAND2X1 U61265 ( .A(n24134), .B(u_decode_scoreboard_q[7]), .Y(n57525) );
  NAND2X1 U61266 ( .A(n42460), .B(n58527), .Y(n57524) );
  NAND2X1 U61267 ( .A(n57525), .B(n57524), .Y(n57526) );
  NAND2X1 U61268 ( .A(n24129), .B(n57526), .Y(n57527) );
  NOR2X1 U61269 ( .A(n57528), .B(n57527), .Y(u_decode_scoreboard_r[7]) );
  NOR2X1 U61270 ( .A(n24136), .B(n24180), .Y(n57533) );
  NAND2X1 U61271 ( .A(n24179), .B(u_decode_scoreboard_q[31]), .Y(n57530) );
  NAND2X1 U61272 ( .A(n42460), .B(n58531), .Y(n57529) );
  NAND2X1 U61273 ( .A(n57530), .B(n57529), .Y(n57531) );
  NAND2X1 U61274 ( .A(n24175), .B(n57531), .Y(n57532) );
  NOR2X1 U61275 ( .A(n57533), .B(n57532), .Y(u_decode_scoreboard_r[31]) );
  NAND2X1 U61276 ( .A(n73427), .B(n57534), .Y(n24144) );
  NOR2X1 U61277 ( .A(n24145), .B(n24135), .Y(n57540) );
  NAND2X1 U61278 ( .A(u_decode_scoreboard_q[6]), .B(n24144), .Y(n57537) );
  NAND2X1 U61279 ( .A(n42460), .B(n57535), .Y(n57536) );
  NAND2X1 U61280 ( .A(n57537), .B(n57536), .Y(n57538) );
  NAND2X1 U61281 ( .A(n24140), .B(n57538), .Y(n57539) );
  NOR2X1 U61282 ( .A(n57540), .B(n57539), .Y(u_decode_scoreboard_r[6]) );
  NAND2X1 U61283 ( .A(n73421), .B(n73427), .Y(n24256) );
  NOR2X1 U61284 ( .A(n24145), .B(n58520), .Y(n57546) );
  NAND2X1 U61285 ( .A(u_decode_scoreboard_q[22]), .B(n24256), .Y(n57543) );
  NAND2X1 U61286 ( .A(n42460), .B(n57541), .Y(n57542) );
  NAND2X1 U61287 ( .A(n57543), .B(n57542), .Y(n57544) );
  NAND2X1 U61288 ( .A(n24252), .B(n57544), .Y(n57545) );
  NOR2X1 U61289 ( .A(n57546), .B(n57545), .Y(u_decode_scoreboard_r[22]) );
  INVX1 U61290 ( .A(n57547), .Y(n36344) );
  INVX1 U61291 ( .A(mem_i_inst_i[15]), .Y(n57548) );
  NOR2X1 U61292 ( .A(n57548), .B(n43405), .Y(net2352) );
  NOR2X1 U61293 ( .A(n8801), .B(n57549), .Y(n57551) );
  NOR2X1 U61294 ( .A(n57600), .B(n57548), .Y(n57550) );
  NOR2X1 U61295 ( .A(n57551), .B(n57550), .Y(n24518) );
  NOR2X1 U61296 ( .A(n24518), .B(n42934), .Y(u_decode_N337) );
  NAND2X1 U61297 ( .A(n44060), .B(n44084), .Y(n73338) );
  NAND2X1 U61298 ( .A(n44280), .B(n73338), .Y(n57552) );
  NAND2X1 U61299 ( .A(u_csr_csr_satp_q_31_), .B(n57552), .Y(n57555) );
  INVX1 U61300 ( .A(n57553), .Y(n73539) );
  NAND2X1 U61301 ( .A(n42304), .B(n44057), .Y(n57554) );
  NAND2X1 U61302 ( .A(n57555), .B(n57554), .Y(u_csr_csr_satp_r[31]) );
  NAND2X1 U61303 ( .A(n57558), .B(n58126), .Y(n57556) );
  NAND2X1 U61304 ( .A(n57557), .B(n57556), .Y(n8561) );
  NOR2X1 U61305 ( .A(n37413), .B(n57558), .Y(u_fetch_N15) );
  NOR2X1 U61306 ( .A(n57559), .B(n42933), .Y(n36342) );
  INVX1 U61307 ( .A(n15219), .Y(n73532) );
  NOR2X1 U61308 ( .A(n73532), .B(n57560), .Y(u_lsu_N98) );
  NOR2X1 U61309 ( .A(n15219), .B(n57560), .Y(u_lsu_N99) );
  NOR2X1 U61310 ( .A(n24429), .B(n73533), .Y(n57562) );
  NOR2X1 U61311 ( .A(n57562), .B(n57561), .Y(n57573) );
  INVX1 U61312 ( .A(n57563), .Y(n57565) );
  NAND2X1 U61313 ( .A(n24397), .B(n73537), .Y(n57564) );
  NAND2X1 U61314 ( .A(n57565), .B(n57564), .Y(n57571) );
  INVX1 U61315 ( .A(n24381), .Y(n57566) );
  NAND2X1 U61316 ( .A(n57567), .B(n57566), .Y(n57569) );
  INVX1 U61317 ( .A(n24389), .Y(n57568) );
  NAND2X1 U61318 ( .A(n57569), .B(n57568), .Y(n57570) );
  NAND2X1 U61319 ( .A(n57571), .B(n57570), .Y(n57572) );
  NOR2X1 U61320 ( .A(n57573), .B(n57572), .Y(n57576) );
  OR2X1 U61321 ( .A(n24412), .B(n24411), .Y(n57574) );
  NOR2X1 U61322 ( .A(n24376), .B(n57574), .Y(n57575) );
  NAND2X1 U61323 ( .A(n57576), .B(n57575), .Y(n57591) );
  NAND2X1 U61324 ( .A(n24407), .B(n57593), .Y(n57578) );
  NAND2X1 U61325 ( .A(n24403), .B(n24379), .Y(n57577) );
  NOR2X1 U61326 ( .A(n57578), .B(n57577), .Y(n57589) );
  NAND2X1 U61327 ( .A(n24384), .B(n57579), .Y(n57584) );
  NOR2X1 U61328 ( .A(n24473), .B(n57580), .Y(n57582) );
  NAND2X1 U61329 ( .A(n57582), .B(n57581), .Y(n57583) );
  NOR2X1 U61330 ( .A(n57584), .B(n57583), .Y(n57587) );
  NAND2X1 U61331 ( .A(n57585), .B(n57595), .Y(n57586) );
  NOR2X1 U61332 ( .A(n57587), .B(n57586), .Y(n57588) );
  NAND2X1 U61333 ( .A(n57589), .B(n57588), .Y(n57590) );
  NOR2X1 U61334 ( .A(n57591), .B(n57590), .Y(u_decode_N793) );
  NAND2X1 U61335 ( .A(n57593), .B(n57592), .Y(n57594) );
  NOR2X1 U61336 ( .A(n57595), .B(n57594), .Y(u_decode_N791) );
  NOR2X1 U61337 ( .A(n28235), .B(n42607), .Y(n57597) );
  NOR2X1 U61338 ( .A(n44639), .B(n28252), .Y(n57596) );
  NAND2X1 U61339 ( .A(n57597), .B(n57596), .Y(u_csr_N3697) );
  INVX1 U61340 ( .A(mem_i_inst_i[18]), .Y(n57598) );
  NOR2X1 U61341 ( .A(n57598), .B(n43404), .Y(net2360) );
  NOR2X1 U61342 ( .A(n8801), .B(n57599), .Y(n57602) );
  NOR2X1 U61343 ( .A(n57600), .B(n57598), .Y(n57601) );
  NOR2X1 U61344 ( .A(n57602), .B(n57601), .Y(n24522) );
  NOR2X1 U61345 ( .A(n24522), .B(n42934), .Y(u_decode_N340) );
  NOR2X1 U61346 ( .A(n43338), .B(n73368), .Y(n57603) );
  NOR2X1 U61347 ( .A(n525), .B(n57603), .Y(n36240) );
  NAND2X1 U61348 ( .A(n57605), .B(n57604), .Y(n57606) );
  NAND2X1 U61349 ( .A(n24117), .B(n57606), .Y(n36238) );
  INVX1 U61350 ( .A(n24161), .Y(n527) );
  NOR2X1 U61351 ( .A(n43344), .B(n42777), .Y(n57607) );
  NOR2X1 U61352 ( .A(n527), .B(n57607), .Y(n36221) );
  NAND2X1 U61353 ( .A(n57609), .B(n57608), .Y(n57610) );
  NAND2X1 U61354 ( .A(n24306), .B(n57610), .Y(n36219) );
  NOR2X1 U61355 ( .A(n43345), .B(n38710), .Y(n57611) );
  NOR2X1 U61356 ( .A(n543), .B(n57611), .Y(n36217) );
  NOR2X1 U61357 ( .A(n40447), .B(n43350), .Y(n57612) );
  NOR2X1 U61358 ( .A(n493), .B(n57612), .Y(n36212) );
  INVX1 U61359 ( .A(n24144), .Y(n529) );
  NOR2X1 U61360 ( .A(n43351), .B(n40514), .Y(n57614) );
  NOR2X1 U61361 ( .A(n529), .B(n57614), .Y(n36202) );
  NOR2X1 U61362 ( .A(n43354), .B(n42781), .Y(n57616) );
  NOR2X1 U61363 ( .A(n501), .B(n57616), .Y(n36200) );
  INVX1 U61364 ( .A(n24270), .Y(n531) );
  NOR2X1 U61365 ( .A(n43360), .B(n57617), .Y(n57618) );
  NOR2X1 U61366 ( .A(n531), .B(n57618), .Y(n36180) );
  INVX1 U61367 ( .A(n24256), .Y(n535) );
  NOR2X1 U61368 ( .A(n43361), .B(n57619), .Y(n57620) );
  NOR2X1 U61369 ( .A(n535), .B(n57620), .Y(n36178) );
  INVX1 U61370 ( .A(n24210), .Y(n547) );
  NOR2X1 U61371 ( .A(n38411), .B(n38844), .Y(n57622) );
  NOR2X1 U61372 ( .A(n547), .B(n57622), .Y(n36006) );
  NOR2X1 U61373 ( .A(n43365), .B(n38085), .Y(n57623) );
  NOR2X1 U61374 ( .A(n539), .B(n57623), .Y(n36002) );
  NAND2X1 U61375 ( .A(n42896), .B(n43370), .Y(n57624) );
  NAND2X1 U61376 ( .A(u_decode_scoreboard_q[7]), .B(n57624), .Y(n35991) );
  NAND2X1 U61377 ( .A(n36609), .B(n57625), .Y(n57626) );
  NAND2X1 U61378 ( .A(u_decode_scoreboard_q[31]), .B(n57626), .Y(n35989) );
  INVX1 U61379 ( .A(n24153), .Y(n571) );
  NOR2X1 U61380 ( .A(n43372), .B(n39318), .Y(n57627) );
  NOR2X1 U61381 ( .A(n571), .B(n57627), .Y(n35983) );
  INVX1 U61382 ( .A(u_csr_N3161), .Y(n73569) );
  INVX1 U61383 ( .A(mem_d_data_rd_i[0]), .Y(n73554) );
  NAND2X1 U61384 ( .A(n57630), .B(n57629), .Y(n57849) );
  INVX1 U61385 ( .A(n57849), .Y(n57631) );
  NAND2X1 U61386 ( .A(n57863), .B(n57631), .Y(n35030) );
  INVX1 U61387 ( .A(n57632), .Y(n57633) );
  INVX1 U61388 ( .A(n57864), .Y(n57855) );
  NOR2X1 U61389 ( .A(n57633), .B(n57855), .Y(n57634) );
  NAND2X1 U61390 ( .A(n57635), .B(n57634), .Y(n35031) );
  INVX1 U61391 ( .A(n57636), .Y(n57638) );
  NOR2X1 U61392 ( .A(n57638), .B(n57637), .Y(n34491) );
  INVX1 U61393 ( .A(n57639), .Y(n57642) );
  INVX1 U61394 ( .A(n57640), .Y(n57641) );
  NOR2X1 U61395 ( .A(n57642), .B(n57641), .Y(n34492) );
  NAND2X1 U61396 ( .A(n57828), .B(n57808), .Y(n57819) );
  INVX1 U61397 ( .A(n57819), .Y(n57643) );
  NAND2X1 U61398 ( .A(n57809), .B(n57643), .Y(n34087) );
  NAND2X1 U61399 ( .A(n43484), .B(n43994), .Y(n68150) );
  INVX1 U61400 ( .A(n68150), .Y(n68425) );
  NOR2X1 U61401 ( .A(n43991), .B(n43482), .Y(n57644) );
  NOR2X1 U61402 ( .A(n68425), .B(n57644), .Y(n57646) );
  NAND2X1 U61403 ( .A(n57793), .B(n57684), .Y(n57645) );
  NOR2X1 U61404 ( .A(n57646), .B(n57645), .Y(n57649) );
  INVX1 U61405 ( .A(n57790), .Y(n57647) );
  NOR2X1 U61406 ( .A(n57647), .B(n42127), .Y(n57648) );
  NAND2X1 U61407 ( .A(n57649), .B(n57648), .Y(n33270) );
  NAND2X1 U61408 ( .A(n43493), .B(n44010), .Y(n57702) );
  INVX1 U61409 ( .A(n57702), .Y(n69790) );
  NAND2X1 U61410 ( .A(n44013), .B(n43495), .Y(n57710) );
  INVX1 U61411 ( .A(n57710), .Y(n57650) );
  NOR2X1 U61412 ( .A(n69790), .B(n57650), .Y(n57652) );
  XNOR2X1 U61413 ( .A(n43766), .B(n43470), .Y(n57651) );
  NOR2X1 U61414 ( .A(n57652), .B(n57651), .Y(n57654) );
  XNOR2X1 U61415 ( .A(n39945), .B(n43747), .Y(n57653) );
  NAND2X1 U61416 ( .A(n57654), .B(n57653), .Y(n33271) );
  NAND2X1 U61417 ( .A(n43797), .B(n43945), .Y(n57656) );
  NAND2X1 U61418 ( .A(n40444), .B(n43936), .Y(n57655) );
  NAND2X1 U61419 ( .A(n57656), .B(n57655), .Y(n31393) );
  NAND2X1 U61420 ( .A(n43481), .B(n43985), .Y(n57658) );
  NAND2X1 U61421 ( .A(n43778), .B(n43975), .Y(n57657) );
  NAND2X1 U61422 ( .A(n57658), .B(n57657), .Y(n31408) );
  NAND2X1 U61423 ( .A(n40460), .B(n43955), .Y(n57660) );
  NAND2X1 U61424 ( .A(n43813), .B(n43965), .Y(n57659) );
  NAND2X1 U61425 ( .A(n57660), .B(n57659), .Y(n31391) );
  INVX1 U61426 ( .A(n57661), .Y(n73434) );
  NAND2X1 U61427 ( .A(n42649), .B(n43929), .Y(n57866) );
  NAND2X1 U61428 ( .A(n40538), .B(n43912), .Y(n57663) );
  NAND2X1 U61429 ( .A(n57663), .B(n57662), .Y(n57850) );
  INVX1 U61430 ( .A(n57850), .Y(n57664) );
  NAND2X1 U61431 ( .A(n57866), .B(n57664), .Y(n32467) );
  NAND2X1 U61432 ( .A(n43794), .B(n43843), .Y(n57766) );
  NOR2X1 U61433 ( .A(n42194), .B(n57665), .Y(n57666) );
  NAND2X1 U61434 ( .A(n57766), .B(n57666), .Y(n32468) );
  NAND2X1 U61435 ( .A(n40477), .B(n43872), .Y(n57812) );
  INVX1 U61436 ( .A(n57812), .Y(n57667) );
  NOR2X1 U61437 ( .A(n57887), .B(n57667), .Y(n32335) );
  NAND2X1 U61438 ( .A(n43783), .B(n38378), .Y(n57754) );
  NAND2X1 U61439 ( .A(n42701), .B(n43920), .Y(n57867) );
  INVX1 U61440 ( .A(n57867), .Y(n57668) );
  NOR2X1 U61441 ( .A(n42195), .B(n57668), .Y(n57669) );
  NAND2X1 U61442 ( .A(n57754), .B(n57669), .Y(n32199) );
  INVX1 U61443 ( .A(n57697), .Y(n57686) );
  NOR2X1 U61444 ( .A(n57686), .B(n57670), .Y(n57671) );
  NAND2X1 U61445 ( .A(n57695), .B(n57671), .Y(n31786) );
  NAND2X1 U61446 ( .A(n43755), .B(n43462), .Y(n57674) );
  NAND2X1 U61447 ( .A(n57674), .B(n62655), .Y(n57675) );
  NAND2X1 U61448 ( .A(n41732), .B(n57675), .Y(n31787) );
  NOR2X1 U61449 ( .A(n57676), .B(n42192), .Y(n31653) );
  INVX1 U61450 ( .A(n57678), .Y(n57884) );
  NOR2X1 U61451 ( .A(n58158), .B(n57884), .Y(n57679) );
  NAND2X1 U61452 ( .A(n57680), .B(n57679), .Y(n31465) );
  NAND2X1 U61453 ( .A(n44020), .B(n44028), .Y(n57682) );
  NAND2X1 U61454 ( .A(n43497), .B(n43502), .Y(n57681) );
  NAND2X1 U61455 ( .A(n57682), .B(n57681), .Y(n57683) );
  NAND2X1 U61456 ( .A(n44812), .B(n57683), .Y(n31450) );
  NAND2X1 U61457 ( .A(n57684), .B(n44816), .Y(n57685) );
  NOR2X1 U61458 ( .A(n57686), .B(n57685), .Y(n57690) );
  NOR2X1 U61459 ( .A(n43504), .B(n44019), .Y(n57688) );
  NOR2X1 U61460 ( .A(n43498), .B(n44027), .Y(n57687) );
  NOR2X1 U61461 ( .A(n57688), .B(n57687), .Y(n57689) );
  NAND2X1 U61462 ( .A(n57690), .B(n57689), .Y(n31451) );
  NAND2X1 U61463 ( .A(n43497), .B(n44019), .Y(n70345) );
  NOR2X1 U61464 ( .A(n44024), .B(n70345), .Y(n57691) );
  NAND2X1 U61465 ( .A(n57691), .B(n43504), .Y(n57694) );
  NAND2X1 U61466 ( .A(n43500), .B(n44027), .Y(n70991) );
  NOR2X1 U61467 ( .A(n43496), .B(n70991), .Y(n57692) );
  NAND2X1 U61468 ( .A(n57692), .B(n44021), .Y(n57693) );
  NAND2X1 U61469 ( .A(n57694), .B(n57693), .Y(n31445) );
  NAND2X1 U61470 ( .A(n43495), .B(n44010), .Y(n57696) );
  NAND2X1 U61471 ( .A(n57696), .B(n57695), .Y(n57700) );
  NAND2X1 U61472 ( .A(n44013), .B(n43493), .Y(n57698) );
  NAND2X1 U61473 ( .A(n57698), .B(n57697), .Y(n57699) );
  MX2X1 U61474 ( .A(n57700), .B(n57699), .S0(n44813), .Y(n31144) );
  NAND2X1 U61475 ( .A(n44004), .B(n43489), .Y(n57701) );
  NOR2X1 U61476 ( .A(n57702), .B(n57701), .Y(n57703) );
  NOR2X1 U61477 ( .A(n31144), .B(n57703), .Y(n31423) );
  NAND2X1 U61478 ( .A(n43999), .B(n44010), .Y(n57705) );
  NAND2X1 U61479 ( .A(n43495), .B(n43489), .Y(n57704) );
  NAND2X1 U61480 ( .A(n57705), .B(n57704), .Y(n57709) );
  NAND2X1 U61481 ( .A(n44013), .B(n44006), .Y(n57707) );
  NAND2X1 U61482 ( .A(n43493), .B(n38310), .Y(n57706) );
  NAND2X1 U61483 ( .A(n57707), .B(n57706), .Y(n57708) );
  MX2X1 U61484 ( .A(n57709), .B(n57708), .S0(n44813), .Y(n57712) );
  NAND2X1 U61485 ( .A(n43999), .B(n43486), .Y(n69400) );
  NOR2X1 U61486 ( .A(n69400), .B(n57710), .Y(n57711) );
  NOR2X1 U61487 ( .A(n57712), .B(n57711), .Y(n31424) );
  NAND2X1 U61488 ( .A(n57714), .B(n57713), .Y(n57715) );
  NAND2X1 U61489 ( .A(n44812), .B(n57715), .Y(n31411) );
  NOR2X1 U61490 ( .A(n44813), .B(n57716), .Y(n57722) );
  INVX1 U61491 ( .A(n57717), .Y(n57720) );
  INVX1 U61492 ( .A(n57718), .Y(n57719) );
  NOR2X1 U61493 ( .A(n57720), .B(n57719), .Y(n57721) );
  NAND2X1 U61494 ( .A(n57722), .B(n57721), .Y(n31412) );
  NOR2X1 U61495 ( .A(n68150), .B(n43479), .Y(n57723) );
  NAND2X1 U61496 ( .A(n57723), .B(n43988), .Y(n57726) );
  NAND2X1 U61497 ( .A(n43477), .B(n43985), .Y(n67698) );
  NOR2X1 U61498 ( .A(n43991), .B(n67698), .Y(n57724) );
  NAND2X1 U61499 ( .A(n57724), .B(n43485), .Y(n57725) );
  NAND2X1 U61500 ( .A(n57726), .B(n57725), .Y(n31409) );
  NOR2X1 U61501 ( .A(n43977), .B(n43949), .Y(n57728) );
  NOR2X1 U61502 ( .A(n43774), .B(n43796), .Y(n57727) );
  NOR2X1 U61503 ( .A(n57728), .B(n57727), .Y(n57729) );
  NOR2X1 U61504 ( .A(n44812), .B(n57729), .Y(n31400) );
  INVX1 U61505 ( .A(n57730), .Y(n57731) );
  NOR2X1 U61506 ( .A(n57731), .B(n44818), .Y(n31401) );
  NAND2X1 U61507 ( .A(n43774), .B(n43975), .Y(n67688) );
  INVX1 U61508 ( .A(n67688), .Y(n67479) );
  NAND2X1 U61509 ( .A(n43797), .B(n67479), .Y(n57732) );
  NOR2X1 U61510 ( .A(n43942), .B(n57732), .Y(n57735) );
  NAND2X1 U61511 ( .A(n43796), .B(n43945), .Y(n66456) );
  NAND2X1 U61512 ( .A(n43778), .B(n43978), .Y(n57733) );
  NOR2X1 U61513 ( .A(n66456), .B(n57733), .Y(n57734) );
  NOR2X1 U61514 ( .A(n57735), .B(n57734), .Y(n31395) );
  NOR2X1 U61515 ( .A(n43968), .B(n43866), .Y(n57737) );
  NOR2X1 U61516 ( .A(n43810), .B(n43821), .Y(n57736) );
  NOR2X1 U61517 ( .A(n57737), .B(n57736), .Y(n57738) );
  NOR2X1 U61518 ( .A(n44812), .B(n57738), .Y(n31383) );
  NOR2X1 U61519 ( .A(n42084), .B(n44818), .Y(n31384) );
  NAND2X1 U61520 ( .A(n43822), .B(n41895), .Y(n57739) );
  NOR2X1 U61521 ( .A(n43861), .B(n57739), .Y(n57742) );
  NAND2X1 U61522 ( .A(n43821), .B(n43862), .Y(n60153) );
  NAND2X1 U61523 ( .A(n43813), .B(n43967), .Y(n57740) );
  NOR2X1 U61524 ( .A(n60153), .B(n57740), .Y(n57741) );
  NOR2X1 U61525 ( .A(n57742), .B(n57741), .Y(n31378) );
  NOR2X1 U61526 ( .A(n42195), .B(n42196), .Y(n57743) );
  NOR2X1 U61527 ( .A(n44812), .B(n57743), .Y(n31371) );
  NOR2X1 U61528 ( .A(n41732), .B(n44815), .Y(n31372) );
  NOR2X1 U61529 ( .A(n43855), .B(n44041), .Y(n57745) );
  NOR2X1 U61530 ( .A(n43759), .B(n43738), .Y(n57744) );
  NOR2X1 U61531 ( .A(n57745), .B(n57744), .Y(n57746) );
  NOR2X1 U61532 ( .A(n44812), .B(n57746), .Y(n31363) );
  NOR2X1 U61533 ( .A(n44036), .B(n43853), .Y(n57748) );
  NOR2X1 U61534 ( .A(n43761), .B(n43740), .Y(n57747) );
  NOR2X1 U61535 ( .A(n57748), .B(n57747), .Y(n57749) );
  NOR2X1 U61536 ( .A(n57749), .B(n44818), .Y(n31364) );
  NAND2X1 U61537 ( .A(n41878), .B(n43740), .Y(n57750) );
  NOR2X1 U61538 ( .A(n44036), .B(n57750), .Y(n57753) );
  NAND2X1 U61539 ( .A(n43736), .B(n44038), .Y(n60497) );
  NAND2X1 U61540 ( .A(n43855), .B(n43760), .Y(n57751) );
  NOR2X1 U61541 ( .A(n60497), .B(n57751), .Y(n57752) );
  NOR2X1 U61542 ( .A(n57753), .B(n57752), .Y(n31358) );
  INVX1 U61543 ( .A(n57754), .Y(n57755) );
  NOR2X1 U61544 ( .A(n42194), .B(n57755), .Y(n57756) );
  NOR2X1 U61545 ( .A(n44812), .B(n57756), .Y(n31351) );
  INVX1 U61546 ( .A(n57757), .Y(n57758) );
  NOR2X1 U61547 ( .A(n57758), .B(n44817), .Y(n31352) );
  NOR2X1 U61548 ( .A(n38387), .B(n43847), .Y(n57760) );
  NOR2X1 U61549 ( .A(n43781), .B(n43791), .Y(n57759) );
  NOR2X1 U61550 ( .A(n57760), .B(n57759), .Y(n57761) );
  NOR2X1 U61551 ( .A(n44812), .B(n57761), .Y(n31343) );
  NOR2X1 U61552 ( .A(n42069), .B(n44817), .Y(n31344) );
  NAND2X1 U61553 ( .A(n43794), .B(n41857), .Y(n57762) );
  NOR2X1 U61554 ( .A(n43841), .B(n57762), .Y(n57765) );
  NAND2X1 U61555 ( .A(n43792), .B(n43843), .Y(n61374) );
  NAND2X1 U61556 ( .A(n43784), .B(n38387), .Y(n57763) );
  NOR2X1 U61557 ( .A(n61374), .B(n57763), .Y(n57764) );
  NOR2X1 U61558 ( .A(n57765), .B(n57764), .Y(n31338) );
  NOR2X1 U61559 ( .A(n44812), .B(n57767), .Y(n31330) );
  NOR2X1 U61560 ( .A(n42068), .B(n44816), .Y(n31331) );
  NOR2X1 U61561 ( .A(n39525), .B(n43744), .Y(n57769) );
  NOR2X1 U61562 ( .A(n39945), .B(n43470), .Y(n57768) );
  NOR2X1 U61563 ( .A(n57769), .B(n57768), .Y(n57770) );
  NOR2X1 U61564 ( .A(n44813), .B(n57770), .Y(n31322) );
  INVX1 U61565 ( .A(n57771), .Y(n57772) );
  NOR2X1 U61566 ( .A(n57772), .B(n44816), .Y(n31323) );
  NAND2X1 U61567 ( .A(n41837), .B(n43470), .Y(n57773) );
  NOR2X1 U61568 ( .A(n43764), .B(n57773), .Y(n57776) );
  NAND2X1 U61569 ( .A(n43764), .B(n43466), .Y(n61661) );
  NAND2X1 U61570 ( .A(n43746), .B(n39946), .Y(n57774) );
  NOR2X1 U61571 ( .A(n61661), .B(n57774), .Y(n57775) );
  NOR2X1 U61572 ( .A(n57776), .B(n57775), .Y(n31317) );
  NOR2X1 U61573 ( .A(n43816), .B(n43805), .Y(n57778) );
  NOR2X1 U61574 ( .A(n40627), .B(n43476), .Y(n57777) );
  NOR2X1 U61575 ( .A(n57778), .B(n57777), .Y(n57779) );
  NOR2X1 U61576 ( .A(n44812), .B(n57779), .Y(n31308) );
  NOR2X1 U61577 ( .A(n43818), .B(n43808), .Y(n57781) );
  NOR2X1 U61578 ( .A(n43472), .B(n43458), .Y(n57780) );
  NOR2X1 U61579 ( .A(n57781), .B(n57780), .Y(n57782) );
  NOR2X1 U61580 ( .A(n57782), .B(n44817), .Y(n31309) );
  NAND2X1 U61581 ( .A(n41836), .B(n43817), .Y(n57783) );
  NOR2X1 U61582 ( .A(n43457), .B(n57783), .Y(n57786) );
  NAND2X1 U61583 ( .A(n38106), .B(n43457), .Y(n62014) );
  NAND2X1 U61584 ( .A(n43807), .B(n43475), .Y(n57784) );
  NOR2X1 U61585 ( .A(n62014), .B(n57784), .Y(n57785) );
  NOR2X1 U61586 ( .A(n57786), .B(n57785), .Y(n31303) );
  NOR2X1 U61587 ( .A(n42192), .B(n42186), .Y(n57787) );
  NOR2X1 U61588 ( .A(n31289), .B(n57787), .Y(n57789) );
  NOR2X1 U61589 ( .A(n43769), .B(n43467), .Y(n57788) );
  NOR2X1 U61590 ( .A(n57789), .B(n57788), .Y(n57791) );
  NAND2X1 U61591 ( .A(n57791), .B(n57790), .Y(n57792) );
  NAND2X1 U61592 ( .A(n44811), .B(n57792), .Y(n31282) );
  NAND2X1 U61593 ( .A(n43768), .B(n43466), .Y(n57794) );
  NAND2X1 U61594 ( .A(n57795), .B(n57794), .Y(n57796) );
  NAND2X1 U61595 ( .A(n44814), .B(n57796), .Y(n31283) );
  NAND2X1 U61596 ( .A(n44814), .B(n31391), .Y(n31266) );
  NOR2X1 U61597 ( .A(n73434), .B(n44815), .Y(n31264) );
  NAND2X1 U61598 ( .A(n57798), .B(n57797), .Y(n57799) );
  NAND2X1 U61599 ( .A(n44811), .B(n57799), .Y(n31252) );
  NOR2X1 U61600 ( .A(n44812), .B(n57800), .Y(n57803) );
  NAND2X1 U61601 ( .A(n57803), .B(n57802), .Y(n31253) );
  NAND2X1 U61602 ( .A(n40461), .B(n43955), .Y(n59840) );
  NOR2X1 U61603 ( .A(n59840), .B(n40470), .Y(n57804) );
  NAND2X1 U61604 ( .A(n57804), .B(n43875), .Y(n57807) );
  NAND2X1 U61605 ( .A(n43869), .B(n40470), .Y(n59664) );
  NOR2X1 U61606 ( .A(n59664), .B(n40461), .Y(n57805) );
  NAND2X1 U61607 ( .A(n57805), .B(n43958), .Y(n57806) );
  NAND2X1 U61608 ( .A(n57807), .B(n57806), .Y(n31250) );
  NAND2X1 U61609 ( .A(n57809), .B(n57808), .Y(n57810) );
  NAND2X1 U61610 ( .A(n44811), .B(n57810), .Y(n31244) );
  NAND2X1 U61611 ( .A(n57812), .B(n57811), .Y(n57813) );
  NAND2X1 U61612 ( .A(n44814), .B(n57813), .Y(n31245) );
  NOR2X1 U61613 ( .A(n44815), .B(n57814), .Y(n57818) );
  NOR2X1 U61614 ( .A(n43885), .B(n43788), .Y(n57816) );
  NOR2X1 U61615 ( .A(n43894), .B(n40483), .Y(n57815) );
  NOR2X1 U61616 ( .A(n57816), .B(n57815), .Y(n57817) );
  NAND2X1 U61617 ( .A(n57818), .B(n57817), .Y(n31230) );
  NOR2X1 U61618 ( .A(n44812), .B(n57819), .Y(n57823) );
  NOR2X1 U61619 ( .A(n43790), .B(n43882), .Y(n57821) );
  NOR2X1 U61620 ( .A(n43722), .B(n43892), .Y(n57820) );
  NOR2X1 U61621 ( .A(n57821), .B(n57820), .Y(n57822) );
  NAND2X1 U61622 ( .A(n57823), .B(n57822), .Y(n31231) );
  NAND2X1 U61623 ( .A(n43879), .B(n40486), .Y(n59959) );
  NOR2X1 U61624 ( .A(n43787), .B(n59959), .Y(n57824) );
  NAND2X1 U61625 ( .A(n57824), .B(n43895), .Y(n57827) );
  NAND2X1 U61626 ( .A(n43889), .B(n43788), .Y(n60711) );
  NOR2X1 U61627 ( .A(n40482), .B(n60711), .Y(n57825) );
  NAND2X1 U61628 ( .A(n57825), .B(n43885), .Y(n57826) );
  NAND2X1 U61629 ( .A(n57827), .B(n57826), .Y(n31228) );
  NAND2X1 U61630 ( .A(n57838), .B(n57828), .Y(n57829) );
  NAND2X1 U61631 ( .A(n44811), .B(n57829), .Y(n31222) );
  NAND2X1 U61632 ( .A(n57831), .B(n57830), .Y(n57832) );
  NAND2X1 U61633 ( .A(n44815), .B(n57832), .Y(n31223) );
  NOR2X1 U61634 ( .A(n57833), .B(n44818), .Y(n57837) );
  NAND2X1 U61635 ( .A(n43908), .B(n43901), .Y(n58905) );
  INVX1 U61636 ( .A(n58905), .Y(n58912) );
  NOR2X1 U61637 ( .A(n58912), .B(n43724), .Y(n57835) );
  NOR2X1 U61638 ( .A(n43901), .B(n42644), .Y(n57834) );
  NOR2X1 U61639 ( .A(n57835), .B(n57834), .Y(n57836) );
  NAND2X1 U61640 ( .A(n57837), .B(n57836), .Y(n31208) );
  NAND2X1 U61641 ( .A(n57838), .B(n44815), .Y(n57839) );
  NOR2X1 U61642 ( .A(n57840), .B(n57839), .Y(n57844) );
  NOR2X1 U61643 ( .A(n42634), .B(n43899), .Y(n57842) );
  NOR2X1 U61644 ( .A(n43727), .B(n43906), .Y(n57841) );
  NOR2X1 U61645 ( .A(n57842), .B(n57841), .Y(n57843) );
  NAND2X1 U61646 ( .A(n57844), .B(n57843), .Y(n31209) );
  NAND2X1 U61647 ( .A(n43903), .B(n42636), .Y(n63611) );
  NOR2X1 U61648 ( .A(n43725), .B(n63611), .Y(n57845) );
  NAND2X1 U61649 ( .A(n57845), .B(n43901), .Y(n57848) );
  NAND2X1 U61650 ( .A(n43724), .B(n43898), .Y(n62511) );
  NOR2X1 U61651 ( .A(n42632), .B(n62511), .Y(n57846) );
  NAND2X1 U61652 ( .A(n57846), .B(n43908), .Y(n57847) );
  NAND2X1 U61653 ( .A(n57848), .B(n57847), .Y(n31206) );
  NAND2X1 U61654 ( .A(n44811), .B(n57849), .Y(n31200) );
  NAND2X1 U61655 ( .A(n44815), .B(n57850), .Y(n31201) );
  NAND2X1 U61656 ( .A(n57852), .B(n57851), .Y(n57853) );
  NAND2X1 U61657 ( .A(n44811), .B(n57853), .Y(n31186) );
  NOR2X1 U61658 ( .A(n44813), .B(n57854), .Y(n57858) );
  NOR2X1 U61659 ( .A(n57856), .B(n57855), .Y(n57857) );
  NAND2X1 U61660 ( .A(n57858), .B(n57857), .Y(n31187) );
  NAND2X1 U61661 ( .A(n40260), .B(n43912), .Y(n63872) );
  NOR2X1 U61662 ( .A(n63872), .B(n43798), .Y(n57859) );
  NAND2X1 U61663 ( .A(n57859), .B(n43923), .Y(n57862) );
  NAND2X1 U61664 ( .A(n43920), .B(n43798), .Y(n64351) );
  NOR2X1 U61665 ( .A(n64351), .B(n40259), .Y(n57860) );
  NAND2X1 U61666 ( .A(n57860), .B(n43915), .Y(n57861) );
  NAND2X1 U61667 ( .A(n57862), .B(n57861), .Y(n31184) );
  NAND2X1 U61668 ( .A(n57864), .B(n57863), .Y(n57865) );
  NAND2X1 U61669 ( .A(n44811), .B(n57865), .Y(n31178) );
  NAND2X1 U61670 ( .A(n57867), .B(n57866), .Y(n57868) );
  NAND2X1 U61671 ( .A(n44815), .B(n57868), .Y(n31179) );
  NAND2X1 U61672 ( .A(n57870), .B(n57869), .Y(n57871) );
  NAND2X1 U61673 ( .A(n44811), .B(n57871), .Y(n31164) );
  NOR2X1 U61674 ( .A(n44813), .B(n57872), .Y(n57877) );
  INVX1 U61675 ( .A(n57873), .Y(n57875) );
  NOR2X1 U61676 ( .A(n57875), .B(n57874), .Y(n57876) );
  NAND2X1 U61677 ( .A(n57877), .B(n57876), .Y(n31165) );
  NAND2X1 U61678 ( .A(n42661), .B(n43929), .Y(n65135) );
  NOR2X1 U61679 ( .A(n65135), .B(n42711), .Y(n57878) );
  NAND2X1 U61680 ( .A(n57878), .B(n43939), .Y(n57881) );
  NAND2X1 U61681 ( .A(n42711), .B(n43936), .Y(n65815) );
  NOR2X1 U61682 ( .A(n65815), .B(n42661), .Y(n57879) );
  NAND2X1 U61683 ( .A(n57879), .B(n43930), .Y(n57880) );
  NAND2X1 U61684 ( .A(n57881), .B(n57880), .Y(n31162) );
  INVX1 U61685 ( .A(n31393), .Y(n57882) );
  NOR2X1 U61686 ( .A(n44813), .B(n57882), .Y(n31158) );
  NAND2X1 U61687 ( .A(n44811), .B(n57883), .Y(n31156) );
  NAND2X1 U61688 ( .A(n44811), .B(n31152), .Y(n31151) );
  NAND2X1 U61689 ( .A(n44811), .B(n41532), .Y(n31138) );
  NOR2X1 U61690 ( .A(n44813), .B(n57884), .Y(n57886) );
  NAND2X1 U61691 ( .A(n43485), .B(n43994), .Y(n57885) );
  NAND2X1 U61692 ( .A(n57886), .B(n57885), .Y(n31139) );
  NOR2X1 U61693 ( .A(n57887), .B(n42127), .Y(n57888) );
  NOR2X1 U61694 ( .A(n44813), .B(n57888), .Y(n31129) );
  NAND2X1 U61695 ( .A(n58426), .B(n58817), .Y(n29787) );
  NAND2X1 U61696 ( .A(opcode_pc_w[5]), .B(opcode_opcode_w[25]), .Y(n29788) );
  NAND2X1 U61697 ( .A(n58431), .B(n73364), .Y(n29766) );
  NAND2X1 U61698 ( .A(opcode_pc_w[6]), .B(opcode_opcode_w[26]), .Y(n29767) );
  NAND2X1 U61699 ( .A(n58436), .B(n58818), .Y(n29745) );
  NAND2X1 U61700 ( .A(opcode_pc_w[7]), .B(opcode_opcode_w[27]), .Y(n29746) );
  NAND2X1 U61701 ( .A(n58441), .B(n58457), .Y(n29724) );
  NAND2X1 U61702 ( .A(opcode_pc_w[8]), .B(opcode_opcode_w[28]), .Y(n29725) );
  NAND2X1 U61703 ( .A(n58446), .B(n73367), .Y(n29703) );
  NAND2X1 U61704 ( .A(opcode_pc_w[9]), .B(opcode_opcode_w[29]), .Y(n29704) );
  NAND2X1 U61705 ( .A(n58280), .B(n57889), .Y(n29941) );
  NAND2X1 U61706 ( .A(n58344), .B(n44844), .Y(n30623) );
  NAND2X1 U61707 ( .A(opcode_pc_w[20]), .B(n44835), .Y(n30621) );
  NAND2X1 U61708 ( .A(n44833), .B(n57890), .Y(n30710) );
  NAND2X1 U61709 ( .A(n58370), .B(n44843), .Y(n30574) );
  NAND2X1 U61710 ( .A(opcode_pc_w[24]), .B(n44835), .Y(n30572) );
  NAND2X1 U61711 ( .A(n58349), .B(n44842), .Y(n30606) );
  NAND2X1 U61712 ( .A(opcode_pc_w[21]), .B(n44835), .Y(n30607) );
  NAND2X1 U61713 ( .A(n58356), .B(n44843), .Y(n30481) );
  NAND2X1 U61714 ( .A(opcode_pc_w[22]), .B(n44835), .Y(n30482) );
  NAND2X1 U61715 ( .A(n58363), .B(n44842), .Y(n30525) );
  NAND2X1 U61716 ( .A(opcode_pc_w[23]), .B(n44835), .Y(n30526) );
  NAND2X1 U61717 ( .A(n58382), .B(n44842), .Y(n30548) );
  NAND2X1 U61718 ( .A(n58377), .B(n44844), .Y(n30329) );
  NAND2X1 U61719 ( .A(opcode_pc_w[25]), .B(n44835), .Y(n30330) );
  INVX1 U61720 ( .A(n57891), .Y(n30429) );
  INVX1 U61721 ( .A(n57892), .Y(n30436) );
  NAND2X1 U61722 ( .A(n57893), .B(n44265), .Y(n58122) );
  INVX1 U61723 ( .A(n58122), .Y(n57991) );
  NAND2X1 U61724 ( .A(n57894), .B(n57991), .Y(n30131) );
  NAND2X1 U61725 ( .A(n57895), .B(n44265), .Y(n58121) );
  INVX1 U61726 ( .A(n58121), .Y(n57993) );
  NAND2X1 U61727 ( .A(mmu_lsu_addr_w[0]), .B(n57993), .Y(n30132) );
  XNOR2X1 U61728 ( .A(n57896), .B(opcode_opcode_w[30]), .Y(n57897) );
  NOR2X1 U61729 ( .A(n43377), .B(n57897), .Y(n57898) );
  XNOR2X1 U61730 ( .A(n43866), .B(n57898), .Y(u_lsu_mem_addr_r[10]) );
  NOR2X1 U61731 ( .A(n2350), .B(n58121), .Y(n30129) );
  NOR2X1 U61732 ( .A(n2351), .B(n58122), .Y(n30130) );
  INVX1 U61733 ( .A(n57899), .Y(n58123) );
  NAND2X1 U61734 ( .A(n43381), .B(u_mmu_request_addr_w[20]), .Y(n57900) );
  NAND2X1 U61735 ( .A(n42421), .B(n57900), .Y(U1_U7_Z_10) );
  MX2X1 U61736 ( .A(n57960), .B(challenge[5]), .S0(n44855), .Y(n17213) );
  NAND2X1 U61737 ( .A(arb_mmu_addr_w[10]), .B(n44257), .Y(n30128) );
  INVX1 U61738 ( .A(n57901), .Y(n57904) );
  XNOR2X1 U61739 ( .A(n44838), .B(n57904), .Y(n57903) );
  NAND2X1 U61740 ( .A(n57903), .B(n43375), .Y(n57906) );
  MX2X1 U61741 ( .A(n37555), .B(n42219), .S0(n57904), .Y(n57905) );
  MX2X1 U61742 ( .A(n57906), .B(n57905), .S0(n43968), .Y(u_lsu_mem_addr_r[11])
         );
  NOR2X1 U61743 ( .A(n2251), .B(n58121), .Y(n30125) );
  NOR2X1 U61744 ( .A(n2252), .B(n58122), .Y(n30126) );
  NAND2X1 U61745 ( .A(n43382), .B(u_mmu_request_addr_w[21]), .Y(n57907) );
  NAND2X1 U61746 ( .A(n42423), .B(n57907), .Y(U1_U7_Z_11) );
  NAND2X1 U61747 ( .A(arb_mmu_addr_w[11]), .B(n44257), .Y(n30124) );
  NAND2X1 U61748 ( .A(n58451), .B(n73539), .Y(n57909) );
  NAND2X1 U61749 ( .A(n27100), .B(n57910), .Y(n57908) );
  NAND2X1 U61750 ( .A(n57909), .B(n57908), .Y(u_csr_csr_satp_r[0]) );
  NAND2X1 U61751 ( .A(n43382), .B(mem_d_data_rd_i[10]), .Y(n57912) );
  NAND2X1 U61752 ( .A(n43380), .B(n57910), .Y(n57911) );
  NAND2X1 U61753 ( .A(n57912), .B(n57911), .Y(U1_U6_Z_12) );
  NOR2X1 U61754 ( .A(n3044), .B(n44262), .Y(n57914) );
  NOR2X1 U61755 ( .A(n8296), .B(n40675), .Y(n57913) );
  NOR2X1 U61756 ( .A(n57914), .B(n57913), .Y(n30117) );
  NAND2X1 U61757 ( .A(n44073), .B(n44261), .Y(n29961) );
  NOR2X1 U61758 ( .A(n73554), .B(n57915), .Y(n57917) );
  NAND2X1 U61759 ( .A(n57917), .B(n57916), .Y(n57921) );
  NOR2X1 U61760 ( .A(n73554), .B(n57918), .Y(n57920) );
  NOR2X1 U61761 ( .A(mem_d_error_i), .B(n28796), .Y(n57919) );
  NAND2X1 U61762 ( .A(n57920), .B(n57919), .Y(n57922) );
  INVX1 U61763 ( .A(n57922), .Y(n58001) );
  NAND2X1 U61764 ( .A(n58001), .B(u_mmu_request_addr_w[12]), .Y(n57924) );
  NAND2X1 U61765 ( .A(mem_d_data_rd_i[10]), .B(n42977), .Y(n57923) );
  NAND2X1 U61766 ( .A(n57924), .B(n57923), .Y(u_mmu_N239) );
  NOR2X1 U61767 ( .A(n2685), .B(n42975), .Y(n57926) );
  NOR2X1 U61768 ( .A(n2683), .B(n40692), .Y(n57925) );
  NOR2X1 U61769 ( .A(n57926), .B(n57925), .Y(n30118) );
  NAND2X1 U61770 ( .A(n58001), .B(u_mmu_request_addr_w[13]), .Y(n57928) );
  NAND2X1 U61771 ( .A(mem_d_data_rd_i[11]), .B(n42978), .Y(n57927) );
  NAND2X1 U61772 ( .A(n57928), .B(n57927), .Y(u_mmu_N240) );
  NOR2X1 U61773 ( .A(n2753), .B(n40693), .Y(n30114) );
  NAND2X1 U61774 ( .A(n73509), .B(n73539), .Y(n57930) );
  NAND2X1 U61775 ( .A(n27064), .B(n73417), .Y(n57929) );
  NAND2X1 U61776 ( .A(n57930), .B(n57929), .Y(u_csr_csr_satp_r[1]) );
  NAND2X1 U61777 ( .A(n43382), .B(mem_d_data_rd_i[11]), .Y(n57932) );
  NAND2X1 U61778 ( .A(n43380), .B(n73417), .Y(n57931) );
  NAND2X1 U61779 ( .A(n57932), .B(n57931), .Y(U1_U6_Z_13) );
  NOR2X1 U61780 ( .A(n3045), .B(n44264), .Y(n57934) );
  NOR2X1 U61781 ( .A(n8298), .B(n40676), .Y(n57933) );
  NOR2X1 U61782 ( .A(n57934), .B(n57933), .Y(n30111) );
  NOR2X1 U61783 ( .A(n8300), .B(n40677), .Y(n30109) );
  NAND2X1 U61784 ( .A(n58452), .B(n73539), .Y(n57936) );
  NAND2X1 U61785 ( .A(n27031), .B(n57937), .Y(n57935) );
  NAND2X1 U61786 ( .A(n57936), .B(n57935), .Y(u_csr_csr_satp_r[2]) );
  NAND2X1 U61787 ( .A(n43382), .B(mem_d_data_rd_i[12]), .Y(n57939) );
  NAND2X1 U61788 ( .A(n43379), .B(n57937), .Y(n57938) );
  NAND2X1 U61789 ( .A(n57939), .B(n57938), .Y(U1_U6_Z_14) );
  NOR2X1 U61790 ( .A(n3046), .B(n44263), .Y(n30110) );
  NAND2X1 U61791 ( .A(n58001), .B(u_mmu_request_addr_w[14]), .Y(n57941) );
  NAND2X1 U61792 ( .A(mem_d_data_rd_i[12]), .B(n42979), .Y(n57940) );
  NAND2X1 U61793 ( .A(n57941), .B(n57940), .Y(u_mmu_N241) );
  NOR2X1 U61794 ( .A(n2154), .B(n42976), .Y(n57943) );
  NOR2X1 U61795 ( .A(n1797), .B(n40694), .Y(n57942) );
  NOR2X1 U61796 ( .A(n57943), .B(n57942), .Y(n30106) );
  NAND2X1 U61797 ( .A(n58453), .B(n73539), .Y(n57945) );
  NAND2X1 U61798 ( .A(n27022), .B(n57946), .Y(n57944) );
  NAND2X1 U61799 ( .A(n57945), .B(n57944), .Y(u_csr_csr_satp_r[3]) );
  NAND2X1 U61800 ( .A(n43382), .B(mem_d_data_rd_i[13]), .Y(n57948) );
  NAND2X1 U61801 ( .A(n43379), .B(n57946), .Y(n57947) );
  NAND2X1 U61802 ( .A(n57948), .B(n57947), .Y(U1_U6_Z_15) );
  NOR2X1 U61803 ( .A(n3047), .B(n44265), .Y(n57950) );
  NOR2X1 U61804 ( .A(n8302), .B(n40675), .Y(n57949) );
  NOR2X1 U61805 ( .A(n57950), .B(n57949), .Y(n30099) );
  NAND2X1 U61806 ( .A(n58001), .B(u_mmu_request_addr_w[15]), .Y(n57952) );
  NAND2X1 U61807 ( .A(mem_d_data_rd_i[13]), .B(n42978), .Y(n57951) );
  NAND2X1 U61808 ( .A(n57952), .B(n57951), .Y(u_mmu_N242) );
  NOR2X1 U61809 ( .A(n2158), .B(n42974), .Y(n57954) );
  NOR2X1 U61810 ( .A(n1869), .B(n40692), .Y(n57953) );
  NOR2X1 U61811 ( .A(n57954), .B(n57953), .Y(n30100) );
  NOR2X1 U61812 ( .A(n8304), .B(n40676), .Y(n30097) );
  NAND2X1 U61813 ( .A(n58454), .B(n73539), .Y(n57956) );
  NAND2X1 U61814 ( .A(n27018), .B(n57957), .Y(n57955) );
  NAND2X1 U61815 ( .A(n57956), .B(n57955), .Y(u_csr_csr_satp_r[4]) );
  NAND2X1 U61816 ( .A(n43382), .B(mem_d_data_rd_i[14]), .Y(n57959) );
  NAND2X1 U61817 ( .A(n43379), .B(n57957), .Y(n57958) );
  NAND2X1 U61818 ( .A(n57959), .B(n57958), .Y(U1_U6_Z_16) );
  MX2X1 U61819 ( .A(n57960), .B(challenge[6]), .S0(n44855), .Y(n17214) );
  NOR2X1 U61820 ( .A(n3048), .B(n44265), .Y(n30098) );
  NAND2X1 U61821 ( .A(n58001), .B(u_mmu_request_addr_w[16]), .Y(n57962) );
  NAND2X1 U61822 ( .A(mem_d_data_rd_i[14]), .B(n42979), .Y(n57961) );
  NAND2X1 U61823 ( .A(n57962), .B(n57961), .Y(u_mmu_N243) );
  NOR2X1 U61824 ( .A(n2516), .B(n40693), .Y(n30096) );
  NAND2X1 U61825 ( .A(n39945), .B(n44083), .Y(n73345) );
  NAND2X1 U61826 ( .A(n44280), .B(n73345), .Y(n57963) );
  NAND2X1 U61827 ( .A(n57963), .B(n73416), .Y(n57965) );
  NAND2X1 U61828 ( .A(n42304), .B(n39937), .Y(n57964) );
  NAND2X1 U61829 ( .A(n57965), .B(n57964), .Y(u_csr_csr_satp_r[5]) );
  NAND2X1 U61830 ( .A(n43382), .B(mem_d_data_rd_i[15]), .Y(n57967) );
  NAND2X1 U61831 ( .A(n43379), .B(n73416), .Y(n57966) );
  NAND2X1 U61832 ( .A(n57967), .B(n57966), .Y(U1_U6_Z_17) );
  NOR2X1 U61833 ( .A(n3049), .B(n44265), .Y(n57969) );
  NOR2X1 U61834 ( .A(n8306), .B(n40677), .Y(n57968) );
  NOR2X1 U61835 ( .A(n57969), .B(n57968), .Y(n30087) );
  NAND2X1 U61836 ( .A(n58001), .B(u_mmu_request_addr_w[17]), .Y(n57971) );
  NAND2X1 U61837 ( .A(mem_d_data_rd_i[15]), .B(n42978), .Y(n57970) );
  NAND2X1 U61838 ( .A(n57971), .B(n57970), .Y(u_mmu_N244) );
  NOR2X1 U61839 ( .A(n2884), .B(n42976), .Y(n57973) );
  NOR2X1 U61840 ( .A(n2882), .B(n40694), .Y(n57972) );
  NOR2X1 U61841 ( .A(n57973), .B(n57972), .Y(n30088) );
  NOR2X1 U61842 ( .A(n8308), .B(n40675), .Y(n30085) );
  NAND2X1 U61843 ( .A(n43845), .B(n44083), .Y(n73170) );
  NAND2X1 U61844 ( .A(n44280), .B(n73170), .Y(n57974) );
  NAND2X1 U61845 ( .A(n57974), .B(n57977), .Y(n57976) );
  NAND2X1 U61846 ( .A(n42304), .B(n43843), .Y(n57975) );
  NAND2X1 U61847 ( .A(n57976), .B(n57975), .Y(u_csr_csr_satp_r[6]) );
  NAND2X1 U61848 ( .A(n43382), .B(mem_d_data_rd_i[16]), .Y(n57979) );
  NAND2X1 U61849 ( .A(n43379), .B(n57977), .Y(n57978) );
  NAND2X1 U61850 ( .A(n57979), .B(n57978), .Y(U1_U6_Z_18) );
  NOR2X1 U61851 ( .A(n3050), .B(n44264), .Y(n30086) );
  NAND2X1 U61852 ( .A(n58001), .B(u_mmu_request_addr_w[18]), .Y(n57981) );
  NAND2X1 U61853 ( .A(n42977), .B(mem_d_data_rd_i[16]), .Y(n57980) );
  NAND2X1 U61854 ( .A(n57981), .B(n57980), .Y(u_mmu_N245) );
  NOR2X1 U61855 ( .A(n2651), .B(n42976), .Y(n57983) );
  NOR2X1 U61856 ( .A(n2650), .B(n40692), .Y(n57982) );
  NOR2X1 U61857 ( .A(n57983), .B(n57982), .Y(n30082) );
  NOR2X1 U61858 ( .A(n8310), .B(n40676), .Y(n30079) );
  NAND2X1 U61859 ( .A(n38386), .B(n44083), .Y(n73352) );
  NAND2X1 U61860 ( .A(n44279), .B(n73352), .Y(n57984) );
  NAND2X1 U61861 ( .A(n57984), .B(n73415), .Y(n57986) );
  NAND2X1 U61862 ( .A(n43836), .B(n38384), .Y(n57985) );
  NAND2X1 U61863 ( .A(n57986), .B(n57985), .Y(u_csr_csr_satp_r[7]) );
  NAND2X1 U61864 ( .A(n43382), .B(mem_d_data_rd_i[17]), .Y(n57988) );
  NAND2X1 U61865 ( .A(n43379), .B(n73415), .Y(n57987) );
  NAND2X1 U61866 ( .A(n57988), .B(n57987), .Y(U1_U6_Z_19) );
  NOR2X1 U61867 ( .A(n3051), .B(n44264), .Y(n30080) );
  NAND2X1 U61868 ( .A(n58001), .B(u_mmu_request_addr_w[19]), .Y(n57990) );
  NAND2X1 U61869 ( .A(n42977), .B(mem_d_data_rd_i[17]), .Y(n57989) );
  NAND2X1 U61870 ( .A(n57990), .B(n57989), .Y(u_mmu_N246) );
  NOR2X1 U61871 ( .A(n2283), .B(n40693), .Y(n30078) );
  NAND2X1 U61872 ( .A(n57992), .B(n57991), .Y(n30073) );
  NAND2X1 U61873 ( .A(mmu_lsu_addr_w[1]), .B(n57993), .Y(n30074) );
  NOR2X1 U61874 ( .A(n8314), .B(n40677), .Y(n30071) );
  NAND2X1 U61875 ( .A(n44040), .B(n44083), .Y(n73359) );
  NAND2X1 U61876 ( .A(n44279), .B(n73359), .Y(n57994) );
  NAND2X1 U61877 ( .A(n57994), .B(n73414), .Y(n57996) );
  NAND2X1 U61878 ( .A(n43836), .B(n44038), .Y(n57995) );
  NAND2X1 U61879 ( .A(n57996), .B(n57995), .Y(u_csr_csr_satp_r[8]) );
  NAND2X1 U61880 ( .A(n43382), .B(mem_d_data_rd_i[18]), .Y(n57998) );
  NAND2X1 U61881 ( .A(n43379), .B(n73414), .Y(n57997) );
  NAND2X1 U61882 ( .A(n57998), .B(n57997), .Y(U1_U6_Z_20) );
  NOR2X1 U61883 ( .A(n3052), .B(n44264), .Y(n30072) );
  NAND2X1 U61884 ( .A(n58001), .B(u_mmu_request_addr_w[20]), .Y(n58000) );
  NAND2X1 U61885 ( .A(n42977), .B(mem_d_data_rd_i[18]), .Y(n57999) );
  NAND2X1 U61886 ( .A(n58000), .B(n57999), .Y(u_mmu_N247) );
  NOR2X1 U61887 ( .A(n2383), .B(n40694), .Y(n30070) );
  NAND2X1 U61888 ( .A(n58001), .B(u_mmu_request_addr_w[21]), .Y(n58003) );
  NAND2X1 U61889 ( .A(n42977), .B(mem_d_data_rd_i[19]), .Y(n58002) );
  NAND2X1 U61890 ( .A(n58003), .B(n58002), .Y(u_mmu_N248) );
  NOR2X1 U61891 ( .A(n2549), .B(n40692), .Y(n30064) );
  NAND2X1 U61892 ( .A(n43855), .B(n44083), .Y(n73179) );
  NAND2X1 U61893 ( .A(n44279), .B(n73179), .Y(n58004) );
  NAND2X1 U61894 ( .A(n58004), .B(n73413), .Y(n58006) );
  NAND2X1 U61895 ( .A(n43836), .B(n43853), .Y(n58005) );
  NAND2X1 U61896 ( .A(n58006), .B(n58005), .Y(u_csr_csr_satp_r[9]) );
  NAND2X1 U61897 ( .A(n43382), .B(mem_d_data_rd_i[19]), .Y(n58008) );
  NAND2X1 U61898 ( .A(n43379), .B(n73413), .Y(n58007) );
  NAND2X1 U61899 ( .A(n58008), .B(n58007), .Y(U1_U6_Z_21) );
  NOR2X1 U61900 ( .A(n3053), .B(n44264), .Y(n58010) );
  NOR2X1 U61901 ( .A(n8316), .B(n40675), .Y(n58009) );
  NOR2X1 U61902 ( .A(n58010), .B(n58009), .Y(n30061) );
  NAND2X1 U61903 ( .A(n43864), .B(n44083), .Y(n73186) );
  NAND2X1 U61904 ( .A(n44279), .B(n73186), .Y(n58011) );
  NAND2X1 U61905 ( .A(n58011), .B(n58014), .Y(n58013) );
  NAND2X1 U61906 ( .A(n43836), .B(n43862), .Y(n58012) );
  NAND2X1 U61907 ( .A(n58013), .B(n58012), .Y(u_csr_csr_satp_r[10]) );
  NAND2X1 U61908 ( .A(n43381), .B(mem_d_data_rd_i[20]), .Y(n58016) );
  NAND2X1 U61909 ( .A(n43379), .B(n58014), .Y(n58015) );
  NAND2X1 U61910 ( .A(n58016), .B(n58015), .Y(U1_U6_Z_22) );
  NOR2X1 U61911 ( .A(n3054), .B(n44265), .Y(n58018) );
  NOR2X1 U61912 ( .A(n8318), .B(n40676), .Y(n58017) );
  NOR2X1 U61913 ( .A(n58018), .B(n58017), .Y(n30055) );
  NOR2X1 U61914 ( .A(n2483), .B(n40693), .Y(n58019) );
  NOR2X1 U61915 ( .A(n30057), .B(n58019), .Y(n30056) );
  NOR2X1 U61916 ( .A(n8320), .B(n40677), .Y(n30053) );
  NAND2X1 U61917 ( .A(n43967), .B(n44083), .Y(n73274) );
  NAND2X1 U61918 ( .A(n44279), .B(n73274), .Y(n58020) );
  NAND2X1 U61919 ( .A(n58020), .B(n73412), .Y(n58022) );
  NAND2X1 U61920 ( .A(n43836), .B(n43965), .Y(n58021) );
  NAND2X1 U61921 ( .A(n58022), .B(n58021), .Y(u_csr_csr_satp_r[11]) );
  NAND2X1 U61922 ( .A(n43381), .B(mem_d_data_rd_i[21]), .Y(n58024) );
  NAND2X1 U61923 ( .A(n43379), .B(n73412), .Y(n58023) );
  NAND2X1 U61924 ( .A(n58024), .B(n58023), .Y(U1_U6_Z_23) );
  NOR2X1 U61925 ( .A(n3055), .B(n44264), .Y(n30054) );
  NOR2X1 U61926 ( .A(n2451), .B(n40694), .Y(n58025) );
  NOR2X1 U61927 ( .A(n30051), .B(n58025), .Y(n30050) );
  NOR2X1 U61928 ( .A(n8322), .B(n40675), .Y(n30047) );
  NAND2X1 U61929 ( .A(n44279), .B(n73267), .Y(n58026) );
  NAND2X1 U61930 ( .A(n58026), .B(n73411), .Y(n58028) );
  NAND2X1 U61931 ( .A(n43836), .B(n43955), .Y(n58027) );
  NAND2X1 U61932 ( .A(n58028), .B(n58027), .Y(u_csr_csr_satp_r[12]) );
  NAND2X1 U61933 ( .A(mem_d_data_rd_i[22]), .B(n58123), .Y(n58030) );
  NAND2X1 U61934 ( .A(n43379), .B(n73411), .Y(n58029) );
  NAND2X1 U61935 ( .A(n58030), .B(n58029), .Y(U1_U6_Z_24) );
  NOR2X1 U61936 ( .A(n3056), .B(n44264), .Y(n30048) );
  NOR2X1 U61937 ( .A(n2850), .B(n40692), .Y(n58031) );
  NOR2X1 U61938 ( .A(n30045), .B(n58031), .Y(n30044) );
  NOR2X1 U61939 ( .A(n8324), .B(n40676), .Y(n30041) );
  NAND2X1 U61940 ( .A(n44279), .B(n73193), .Y(n58032) );
  NAND2X1 U61941 ( .A(n58032), .B(n58035), .Y(n58034) );
  NAND2X1 U61942 ( .A(n43836), .B(n43872), .Y(n58033) );
  NAND2X1 U61943 ( .A(n58034), .B(n58033), .Y(u_csr_csr_satp_r[13]) );
  NAND2X1 U61944 ( .A(mem_d_data_rd_i[23]), .B(n58123), .Y(n58037) );
  NAND2X1 U61945 ( .A(n43378), .B(n58035), .Y(n58036) );
  NAND2X1 U61946 ( .A(n58037), .B(n58036), .Y(U1_U6_Z_25) );
  NOR2X1 U61947 ( .A(n3057), .B(n44265), .Y(n30042) );
  NOR2X1 U61948 ( .A(n2817), .B(n40693), .Y(n30040) );
  NOR2X1 U61949 ( .A(n2617), .B(n40694), .Y(n30034) );
  NAND2X1 U61950 ( .A(n44279), .B(n73200), .Y(n58038) );
  NAND2X1 U61951 ( .A(n58038), .B(n58041), .Y(n58040) );
  NAND2X1 U61952 ( .A(n43836), .B(n43882), .Y(n58039) );
  NAND2X1 U61953 ( .A(n58040), .B(n58039), .Y(u_csr_csr_satp_r[14]) );
  NAND2X1 U61954 ( .A(n43381), .B(mem_d_data_rd_i[24]), .Y(n58043) );
  NAND2X1 U61955 ( .A(n43378), .B(n58041), .Y(n58042) );
  NAND2X1 U61956 ( .A(n58043), .B(n58042), .Y(U1_U6_Z_26) );
  NOR2X1 U61957 ( .A(n3058), .B(n44263), .Y(n58045) );
  NOR2X1 U61958 ( .A(n8326), .B(n40677), .Y(n58044) );
  NOR2X1 U61959 ( .A(n58045), .B(n58044), .Y(n30031) );
  NOR2X1 U61960 ( .A(n2785), .B(n40692), .Y(n30028) );
  NAND2X1 U61961 ( .A(n44279), .B(n73207), .Y(n58046) );
  NAND2X1 U61962 ( .A(n58046), .B(n58049), .Y(n58048) );
  NAND2X1 U61963 ( .A(n43836), .B(n43892), .Y(n58047) );
  NAND2X1 U61964 ( .A(n58048), .B(n58047), .Y(u_csr_csr_satp_r[15]) );
  NAND2X1 U61965 ( .A(n43381), .B(mem_d_data_rd_i[25]), .Y(n58051) );
  NAND2X1 U61966 ( .A(n43378), .B(n58049), .Y(n58050) );
  NAND2X1 U61967 ( .A(n58051), .B(n58050), .Y(U1_U6_Z_27) );
  NOR2X1 U61968 ( .A(n3059), .B(n44263), .Y(n58053) );
  NOR2X1 U61969 ( .A(n8328), .B(n40675), .Y(n58052) );
  NOR2X1 U61970 ( .A(n58053), .B(n58052), .Y(n30025) );
  NOR2X1 U61971 ( .A(n8330), .B(n40676), .Y(n30023) );
  NAND2X1 U61972 ( .A(n44279), .B(n73214), .Y(n58054) );
  NAND2X1 U61973 ( .A(n58054), .B(n73410), .Y(n58056) );
  NAND2X1 U61974 ( .A(n43836), .B(n43898), .Y(n58055) );
  NAND2X1 U61975 ( .A(n58056), .B(n58055), .Y(u_csr_csr_satp_r[16]) );
  NAND2X1 U61976 ( .A(mem_d_data_rd_i[26]), .B(n58123), .Y(n58058) );
  NAND2X1 U61977 ( .A(n43378), .B(n73410), .Y(n58057) );
  NAND2X1 U61978 ( .A(n58058), .B(n58057), .Y(U1_U6_Z_28) );
  NOR2X1 U61979 ( .A(n3060), .B(n44263), .Y(n30024) );
  NOR2X1 U61980 ( .A(n1870), .B(n40693), .Y(n58059) );
  NOR2X1 U61981 ( .A(n30021), .B(n58059), .Y(n30020) );
  NOR2X1 U61982 ( .A(n8332), .B(n40677), .Y(n30017) );
  NAND2X1 U61983 ( .A(n44279), .B(n73222), .Y(n58060) );
  NAND2X1 U61984 ( .A(n58060), .B(n73409), .Y(n58062) );
  NAND2X1 U61985 ( .A(n43836), .B(n43906), .Y(n58061) );
  NAND2X1 U61986 ( .A(n58062), .B(n58061), .Y(u_csr_csr_satp_r[17]) );
  NAND2X1 U61987 ( .A(mem_d_data_rd_i[27]), .B(n58123), .Y(n58064) );
  NAND2X1 U61988 ( .A(n43378), .B(n73409), .Y(n58063) );
  NAND2X1 U61989 ( .A(n58064), .B(n58063), .Y(U1_U6_Z_29) );
  NOR2X1 U61990 ( .A(n3061), .B(n44263), .Y(n30018) );
  NOR2X1 U61991 ( .A(n1801), .B(n40694), .Y(n30016) );
  XOR2X1 U61992 ( .A(n58066), .B(n58065), .Y(n58067) );
  NOR2X1 U61993 ( .A(n43377), .B(n58067), .Y(n58068) );
  XOR2X1 U61994 ( .A(n43458), .B(n58068), .Y(u_lsu_mem_addr_r[2]) );
  NOR2X1 U61995 ( .A(n1861), .B(n58121), .Y(n30011) );
  NOR2X1 U61996 ( .A(n1862), .B(n58122), .Y(n30012) );
  NAND2X1 U61997 ( .A(n43381), .B(u_mmu_request_addr_w[12]), .Y(n58070) );
  NAND2X1 U61998 ( .A(n43378), .B(u_mmu_request_addr_w[22]), .Y(n58069) );
  NAND2X1 U61999 ( .A(n58070), .B(n58069), .Y(U1_U7_Z_2) );
  NAND2X1 U62000 ( .A(arb_mmu_addr_w[2]), .B(n44257), .Y(n30010) );
  NOR2X1 U62001 ( .A(n8336), .B(n40675), .Y(n30007) );
  NAND2X1 U62002 ( .A(n44279), .B(n73230), .Y(n58071) );
  NAND2X1 U62003 ( .A(n58071), .B(n58074), .Y(n58073) );
  NAND2X1 U62004 ( .A(n43836), .B(n43911), .Y(n58072) );
  NAND2X1 U62005 ( .A(n58073), .B(n58072), .Y(u_csr_csr_satp_r[18]) );
  NAND2X1 U62006 ( .A(mem_d_data_rd_i[28]), .B(n58123), .Y(n58076) );
  NAND2X1 U62007 ( .A(n43378), .B(n58074), .Y(n58075) );
  NAND2X1 U62008 ( .A(n58076), .B(n58075), .Y(U1_U6_Z_30) );
  NOR2X1 U62009 ( .A(n3062), .B(n44262), .Y(n30008) );
  NOR2X1 U62010 ( .A(n1871), .B(n40692), .Y(n58077) );
  NOR2X1 U62011 ( .A(n30005), .B(n58077), .Y(n30004) );
  NOR2X1 U62012 ( .A(n1872), .B(n40693), .Y(n29998) );
  NAND2X1 U62013 ( .A(n44278), .B(n73238), .Y(n58079) );
  NAND2X1 U62014 ( .A(n58079), .B(n73408), .Y(n58081) );
  NAND2X1 U62015 ( .A(n43835), .B(n43920), .Y(n58080) );
  NAND2X1 U62016 ( .A(n58081), .B(n58080), .Y(u_csr_csr_satp_r[19]) );
  NAND2X1 U62017 ( .A(mem_d_data_rd_i[29]), .B(n58123), .Y(n58083) );
  NAND2X1 U62018 ( .A(n43378), .B(n73408), .Y(n58082) );
  NAND2X1 U62019 ( .A(n58083), .B(n58082), .Y(U1_U6_Z_31) );
  NOR2X1 U62020 ( .A(n3063), .B(n44262), .Y(n58086) );
  NOR2X1 U62021 ( .A(n8338), .B(n40676), .Y(n58085) );
  NOR2X1 U62022 ( .A(n58086), .B(n58085), .Y(n29995) );
  XNOR2X1 U62023 ( .A(n58088), .B(n58087), .Y(n58089) );
  NOR2X1 U62024 ( .A(n43377), .B(n58089), .Y(n58090) );
  XNOR2X1 U62025 ( .A(n43476), .B(n58090), .Y(u_lsu_mem_addr_r[3]) );
  NOR2X1 U62026 ( .A(n1863), .B(n58121), .Y(n29993) );
  NOR2X1 U62027 ( .A(n1864), .B(n58122), .Y(n29994) );
  NAND2X1 U62028 ( .A(n43381), .B(u_mmu_request_addr_w[13]), .Y(n58092) );
  NAND2X1 U62029 ( .A(n43378), .B(u_mmu_request_addr_w[23]), .Y(n58091) );
  NAND2X1 U62030 ( .A(n58092), .B(n58091), .Y(U1_U7_Z_3) );
  NAND2X1 U62031 ( .A(arb_mmu_addr_w[3]), .B(n44257), .Y(n29992) );
  XOR2X1 U62032 ( .A(n58094), .B(n58093), .Y(n58095) );
  NOR2X1 U62033 ( .A(n43377), .B(n58095), .Y(n58096) );
  XOR2X1 U62034 ( .A(n43467), .B(n58096), .Y(u_lsu_mem_addr_r[4]) );
  NOR2X1 U62035 ( .A(n1865), .B(n58121), .Y(n29989) );
  NOR2X1 U62036 ( .A(n1866), .B(n58122), .Y(n29990) );
  NAND2X1 U62037 ( .A(n43381), .B(u_mmu_request_addr_w[14]), .Y(n58098) );
  NAND2X1 U62038 ( .A(n43378), .B(u_mmu_request_addr_w[24]), .Y(n58097) );
  NAND2X1 U62039 ( .A(n58098), .B(n58097), .Y(U1_U7_Z_4) );
  NAND2X1 U62040 ( .A(arb_mmu_addr_w[4]), .B(n44257), .Y(n29988) );
  XNOR2X1 U62041 ( .A(n58099), .B(opcode_opcode_w[25]), .Y(n58100) );
  NOR2X1 U62042 ( .A(n43376), .B(n58100), .Y(n58101) );
  XNOR2X1 U62043 ( .A(n39944), .B(n58101), .Y(u_lsu_mem_addr_r[5]) );
  NOR2X1 U62044 ( .A(n1867), .B(n58121), .Y(n29985) );
  NOR2X1 U62045 ( .A(n1868), .B(n58122), .Y(n29986) );
  NAND2X1 U62046 ( .A(n43381), .B(u_mmu_request_addr_w[15]), .Y(n58103) );
  NAND2X1 U62047 ( .A(n43378), .B(u_mmu_request_addr_w[25]), .Y(n58102) );
  NAND2X1 U62048 ( .A(n58103), .B(n58102), .Y(U1_U7_Z_5) );
  NAND2X1 U62049 ( .A(arb_mmu_addr_w[5]), .B(n44257), .Y(n29984) );
  XNOR2X1 U62050 ( .A(n58104), .B(opcode_opcode_w[26]), .Y(n58105) );
  NOR2X1 U62051 ( .A(n43377), .B(n58105), .Y(n58106) );
  XNOR2X1 U62052 ( .A(n43847), .B(n58106), .Y(u_lsu_mem_addr_r[6]) );
  NOR2X1 U62053 ( .A(n2316), .B(n58121), .Y(n29981) );
  NOR2X1 U62054 ( .A(n2317), .B(n58122), .Y(n29982) );
  NAND2X1 U62055 ( .A(n43381), .B(u_mmu_request_addr_w[16]), .Y(n58108) );
  NAND2X1 U62056 ( .A(n43378), .B(u_mmu_request_addr_w[26]), .Y(n58107) );
  NAND2X1 U62057 ( .A(n58108), .B(n58107), .Y(U1_U7_Z_6) );
  NAND2X1 U62058 ( .A(arb_mmu_addr_w[6]), .B(n44257), .Y(n29980) );
  XNOR2X1 U62059 ( .A(n58109), .B(opcode_opcode_w[27]), .Y(n58110) );
  NOR2X1 U62060 ( .A(n43376), .B(n58110), .Y(n58111) );
  XNOR2X1 U62061 ( .A(n38387), .B(n58111), .Y(u_lsu_mem_addr_r[7]) );
  NOR2X1 U62062 ( .A(n2581), .B(n58121), .Y(n29977) );
  NOR2X1 U62063 ( .A(n2582), .B(n58122), .Y(n29978) );
  NAND2X1 U62064 ( .A(n43381), .B(u_mmu_request_addr_w[17]), .Y(n58113) );
  NAND2X1 U62065 ( .A(n43379), .B(u_mmu_request_addr_w[27]), .Y(n58112) );
  NAND2X1 U62066 ( .A(n58113), .B(n58112), .Y(U1_U7_Z_7) );
  NAND2X1 U62067 ( .A(arb_mmu_addr_w[7]), .B(n44257), .Y(n29976) );
  XNOR2X1 U62068 ( .A(n58114), .B(opcode_opcode_w[28]), .Y(n58115) );
  NOR2X1 U62069 ( .A(n43376), .B(n58115), .Y(n58116) );
  NOR2X1 U62070 ( .A(n2716), .B(n58121), .Y(n29973) );
  NOR2X1 U62071 ( .A(n2717), .B(n58122), .Y(n29974) );
  NAND2X1 U62072 ( .A(n43381), .B(u_mmu_request_addr_w[18]), .Y(n58117) );
  NAND2X1 U62073 ( .A(n42420), .B(n58117), .Y(U1_U7_Z_8) );
  NAND2X1 U62074 ( .A(arb_mmu_addr_w[8]), .B(n44257), .Y(n29972) );
  XNOR2X1 U62075 ( .A(n58118), .B(opcode_opcode_w[29]), .Y(n58119) );
  NOR2X1 U62076 ( .A(n43376), .B(n58119), .Y(n58120) );
  NOR2X1 U62077 ( .A(n2419), .B(n58121), .Y(n29967) );
  NOR2X1 U62078 ( .A(n2420), .B(n58122), .Y(n29968) );
  NAND2X1 U62079 ( .A(n43382), .B(u_mmu_request_addr_w[19]), .Y(n58124) );
  NAND2X1 U62080 ( .A(n42422), .B(n58124), .Y(U1_U7_Z_9) );
  NAND2X1 U62081 ( .A(arb_mmu_addr_w[9]), .B(n44258), .Y(n29966) );
  INVX1 U62082 ( .A(u_lsu_N226), .Y(n58125) );
  NOR2X1 U62083 ( .A(n43734), .B(n58125), .Y(u_lsu_N194) );
  NOR2X1 U62084 ( .A(n43756), .B(n58125), .Y(u_lsu_N195) );
  NOR2X1 U62085 ( .A(n43817), .B(n58125), .Y(u_lsu_N196) );
  NOR2X1 U62086 ( .A(n43807), .B(n58125), .Y(u_lsu_N197) );
  NOR2X1 U62087 ( .A(n43769), .B(n58125), .Y(u_lsu_N198) );
  NOR2X1 U62088 ( .A(n43746), .B(n58125), .Y(u_lsu_N199) );
  NOR2X1 U62089 ( .A(n43793), .B(n58125), .Y(u_lsu_N200) );
  NOR2X1 U62090 ( .A(n43784), .B(n58125), .Y(u_lsu_N201) );
  NAND2X1 U62091 ( .A(n58127), .B(n58126), .Y(n29677) );
  NAND2X1 U62092 ( .A(n44863), .B(n58128), .Y(n29644) );
  NOR2X1 U62093 ( .A(n24422), .B(n58129), .Y(u_decode_N779) );
  NAND2X1 U62094 ( .A(n42757), .B(n40018), .Y(n58131) );
  NOR2X1 U62095 ( .A(n29634), .B(n58131), .Y(n29633) );
  NAND2X1 U62096 ( .A(n44833), .B(opcode_opcode_w[30]), .Y(n25635) );
  INVX1 U62097 ( .A(u_csr_N3162), .Y(n73568) );
  NOR2X1 U62098 ( .A(opcode_opcode_w[29]), .B(n73568), .Y(n58133) );
  NAND2X1 U62099 ( .A(opcode_opcode_w[28]), .B(n73569), .Y(n58132) );
  NOR2X1 U62100 ( .A(n58133), .B(n58132), .Y(n29631) );
  NAND2X1 U62101 ( .A(n73568), .B(opcode_opcode_w[29]), .Y(n29630) );
  INVX1 U62102 ( .A(n27326), .Y(n73543) );
  INVX1 U62103 ( .A(n58213), .Y(n58134) );
  NOR2X1 U62104 ( .A(n27326), .B(n58134), .Y(n29570) );
  NAND2X1 U62105 ( .A(n43607), .B(n58822), .Y(n58135) );
  INVX1 U62106 ( .A(n28813), .Y(n73428) );
  NAND2X1 U62107 ( .A(n58135), .B(n73428), .Y(n58977) );
  INVX1 U62108 ( .A(n58977), .Y(n59114) );
  NAND2X1 U62109 ( .A(n42453), .B(n43608), .Y(n59112) );
  NOR2X1 U62110 ( .A(n42651), .B(n43798), .Y(n58145) );
  NOR2X1 U62111 ( .A(n42632), .B(n40260), .Y(n58144) );
  NOR2X1 U62112 ( .A(n43788), .B(n43724), .Y(n58143) );
  NOR2X1 U62113 ( .A(n40485), .B(n40472), .Y(n58142) );
  NOR2X1 U62114 ( .A(n72820), .B(n40461), .Y(n58141) );
  NOR2X1 U62115 ( .A(n43758), .B(n43821), .Y(n58140) );
  NOR2X1 U62116 ( .A(n43736), .B(n39164), .Y(n58139) );
  NOR2X1 U62117 ( .A(n43791), .B(n43744), .Y(n58138) );
  NOR2X1 U62118 ( .A(n43804), .B(n43766), .Y(n58137) );
  NOR2X1 U62119 ( .A(n43752), .B(n43816), .Y(n58136) );
  NAND2X1 U62120 ( .A(n58136), .B(n43734), .Y(n58988) );
  INVX1 U62121 ( .A(n58988), .Y(n58990) );
  NAND2X1 U62122 ( .A(n58137), .B(n58990), .Y(n58998) );
  INVX1 U62123 ( .A(n58998), .Y(n59000) );
  NAND2X1 U62124 ( .A(n58138), .B(n59000), .Y(n59008) );
  INVX1 U62125 ( .A(n59008), .Y(n59010) );
  NAND2X1 U62126 ( .A(n58139), .B(n59010), .Y(n59018) );
  INVX1 U62127 ( .A(n59018), .Y(n59020) );
  NAND2X1 U62128 ( .A(n58140), .B(n59020), .Y(n59028) );
  INVX1 U62129 ( .A(n59028), .Y(n59030) );
  NAND2X1 U62130 ( .A(n58141), .B(n59030), .Y(n59038) );
  INVX1 U62131 ( .A(n59038), .Y(n59040) );
  NAND2X1 U62132 ( .A(n58142), .B(n59040), .Y(n59048) );
  INVX1 U62133 ( .A(n59048), .Y(n59050) );
  NAND2X1 U62134 ( .A(n58143), .B(n59050), .Y(n59058) );
  INVX1 U62135 ( .A(n59058), .Y(n59060) );
  NAND2X1 U62136 ( .A(n58144), .B(n59060), .Y(n59068) );
  INVX1 U62137 ( .A(n59068), .Y(n59070) );
  NAND2X1 U62138 ( .A(n58145), .B(n59070), .Y(n59075) );
  NOR2X1 U62139 ( .A(n59081), .B(n43776), .Y(n58146) );
  NAND2X1 U62140 ( .A(n43797), .B(n58146), .Y(n59088) );
  INVX1 U62141 ( .A(n59088), .Y(n58147) );
  NAND2X1 U62142 ( .A(n43481), .B(n58147), .Y(n59094) );
  NOR2X1 U62143 ( .A(n43487), .B(n59094), .Y(n58148) );
  NAND2X1 U62144 ( .A(n43485), .B(n58148), .Y(n59101) );
  INVX1 U62145 ( .A(n59101), .Y(n58149) );
  NAND2X1 U62146 ( .A(n58149), .B(n43495), .Y(n59105) );
  INVX1 U62147 ( .A(n59105), .Y(n58150) );
  NAND2X1 U62148 ( .A(n58150), .B(n43498), .Y(n59109) );
  INVX1 U62149 ( .A(n59109), .Y(n58151) );
  NAND2X1 U62150 ( .A(n43504), .B(n58151), .Y(n59115) );
  INVX1 U62151 ( .A(n59115), .Y(n58152) );
  NAND2X1 U62152 ( .A(n58152), .B(n43520), .Y(n58157) );
  NOR2X1 U62153 ( .A(n42980), .B(n58157), .Y(n58153) );
  NOR2X1 U62154 ( .A(n43445), .B(n58153), .Y(n58154) );
  NOR2X1 U62155 ( .A(n43611), .B(n58154), .Y(u_muldiv_N327) );
  NAND2X1 U62156 ( .A(u_csr_writeback_en_q), .B(n37332), .Y(n29321) );
  INVX1 U62157 ( .A(n29321), .Y(n58155) );
  NAND2X1 U62158 ( .A(u_csr_writeback_idx_q[3]), .B(n58155), .Y(n1064) );
  NAND2X1 U62159 ( .A(u_csr_writeback_idx_q[0]), .B(n58155), .Y(n1053) );
  INVX1 U62160 ( .A(n1053), .Y(n29309) );
  NAND2X1 U62161 ( .A(n43383), .B(n58156), .Y(n29256) );
  INVX1 U62162 ( .A(n29256), .Y(n73407) );
  NAND2X1 U62163 ( .A(n43386), .B(n21437), .Y(n29223) );
  INVX1 U62164 ( .A(n29223), .Y(n73406) );
  INVX1 U62165 ( .A(n1064), .Y(n29144) );
  NAND2X1 U62166 ( .A(n58815), .B(n58811), .Y(n28946) );
  NAND2X1 U62167 ( .A(n28934), .B(n73430), .Y(n28932) );
  NAND2X1 U62168 ( .A(opcode_opcode_w[9]), .B(n73374), .Y(n28910) );
  NAND2X1 U62169 ( .A(opcode_opcode_w[8]), .B(n73374), .Y(n28908) );
  NAND2X1 U62170 ( .A(n58158), .B(n58157), .Y(n58160) );
  NAND2X1 U62171 ( .A(n58160), .B(n58159), .Y(n58161) );
  NAND2X1 U62172 ( .A(opcode_instr_w_51), .B(n58161), .Y(n58163) );
  NAND2X1 U62173 ( .A(n8887), .B(n44057), .Y(n58162) );
  NAND2X1 U62174 ( .A(n58163), .B(n58162), .Y(n28848) );
  NAND2X1 U62175 ( .A(n58165), .B(n58164), .Y(n28845) );
  INVX1 U62176 ( .A(n28797), .Y(n73538) );
  NOR2X1 U62177 ( .A(n42975), .B(n58166), .Y(n58167) );
  NAND2X1 U62178 ( .A(u_mmu_store_q[2]), .B(n42464), .Y(n58171) );
  NAND2X1 U62179 ( .A(n58176), .B(n58216), .Y(n58168) );
  NAND2X1 U62180 ( .A(n44073), .B(n58168), .Y(n58169) );
  AND2X1 U62181 ( .A(n58169), .B(n44262), .Y(n58195) );
  NAND2X1 U62182 ( .A(n58195), .B(n37327), .Y(n58170) );
  NAND2X1 U62183 ( .A(n58171), .B(n58170), .Y(mem_d_wr_o[2]) );
  NAND2X1 U62184 ( .A(u_mmu_store_q[1]), .B(n42464), .Y(n58173) );
  NAND2X1 U62185 ( .A(n58195), .B(n37328), .Y(n58172) );
  NAND2X1 U62186 ( .A(n58173), .B(n58172), .Y(mem_d_wr_o[1]) );
  NOR2X1 U62187 ( .A(n29961), .B(n37425), .Y(n58175) );
  NOR2X1 U62188 ( .A(n8574), .B(n44258), .Y(n58174) );
  NOR2X1 U62189 ( .A(n58175), .B(n58174), .Y(n58178) );
  NAND2X1 U62190 ( .A(n58176), .B(n58218), .Y(n58177) );
  NOR2X1 U62191 ( .A(n58178), .B(n58177), .Y(n58182) );
  NAND2X1 U62192 ( .A(n58179), .B(n44261), .Y(n58180) );
  NOR2X1 U62193 ( .A(n8574), .B(n58180), .Y(n58181) );
  NOR2X1 U62194 ( .A(n58182), .B(n58181), .Y(n28744) );
  NAND2X1 U62195 ( .A(n58183), .B(n44258), .Y(n28745) );
  NAND2X1 U62196 ( .A(u_mmu_store_q[3]), .B(n42464), .Y(n58186) );
  NAND2X1 U62197 ( .A(n58195), .B(n58184), .Y(n58185) );
  NAND2X1 U62198 ( .A(n58186), .B(n58185), .Y(mem_d_wr_o[3]) );
  NAND2X1 U62199 ( .A(n58216), .B(n58194), .Y(n58187) );
  NOR2X1 U62200 ( .A(n58188), .B(n58187), .Y(n58193) );
  NOR2X1 U62201 ( .A(n58191), .B(n58190), .Y(n58192) );
  NOR2X1 U62202 ( .A(n58193), .B(n58192), .Y(n28741) );
  NAND2X1 U62203 ( .A(u_mmu_store_q[0]), .B(n42464), .Y(n58197) );
  NAND2X1 U62204 ( .A(n58195), .B(n58194), .Y(n58196) );
  NAND2X1 U62205 ( .A(n58197), .B(n58196), .Y(mem_d_wr_o[0]) );
  NOR2X1 U62206 ( .A(opcode_opcode_w[27]), .B(n58816), .Y(n58198) );
  NAND2X1 U62207 ( .A(n58198), .B(n73367), .Y(n28621) );
  INVX1 U62208 ( .A(n28621), .Y(n73405) );
  NAND2X1 U62209 ( .A(n38501), .B(n73405), .Y(n58199) );
  NAND2X1 U62210 ( .A(n38501), .B(n58233), .Y(n58208) );
  NAND2X1 U62211 ( .A(n58199), .B(n58208), .Y(n26261) );
  NAND2X1 U62212 ( .A(n26261), .B(n27964), .Y(n58209) );
  INVX1 U62213 ( .A(n58209), .Y(n73404) );
  NAND2X1 U62214 ( .A(n58200), .B(n24943), .Y(n58201) );
  NAND2X1 U62215 ( .A(n38824), .B(n58201), .Y(n896) );
  INVX1 U62216 ( .A(n896), .Y(n73403) );
  NAND2X1 U62217 ( .A(n38501), .B(n58243), .Y(n58228) );
  NAND2X1 U62218 ( .A(n58228), .B(n58202), .Y(n28636) );
  NAND2X1 U62219 ( .A(n39198), .B(n73405), .Y(n58255) );
  NOR2X1 U62220 ( .A(n58254), .B(n38501), .Y(n58203) );
  NAND2X1 U62221 ( .A(n58203), .B(n38464), .Y(n58204) );
  NAND2X1 U62222 ( .A(n73506), .B(n58204), .Y(n72829) );
  NAND2X1 U62223 ( .A(n58255), .B(n72829), .Y(n27104) );
  NAND2X1 U62224 ( .A(n39197), .B(n58233), .Y(n58227) );
  NAND2X1 U62225 ( .A(n58205), .B(n58227), .Y(n58206) );
  NOR2X1 U62226 ( .A(n42323), .B(n58206), .Y(n28633) );
  NAND2X1 U62227 ( .A(n28621), .B(n24942), .Y(n58207) );
  NAND2X1 U62228 ( .A(n38825), .B(n58207), .Y(n889) );
  INVX1 U62229 ( .A(n889), .Y(n73402) );
  NAND2X1 U62230 ( .A(n38492), .B(n58243), .Y(n58248) );
  NAND2X1 U62231 ( .A(n73506), .B(n38609), .Y(n58252) );
  NAND2X1 U62232 ( .A(n58248), .B(n58252), .Y(n27401) );
  NOR2X1 U62233 ( .A(n27401), .B(n73539), .Y(n28629) );
  INVX1 U62234 ( .A(n58208), .Y(n58266) );
  INVX1 U62235 ( .A(n26129), .Y(n73577) );
  NAND2X1 U62236 ( .A(n26361), .B(n73230), .Y(n28582) );
  NOR2X1 U62237 ( .A(n58230), .B(n58209), .Y(n58210) );
  NAND2X1 U62238 ( .A(n43911), .B(n58210), .Y(n28579) );
  NAND2X1 U62239 ( .A(n58212), .B(n58211), .Y(n28563) );
  INVX1 U62240 ( .A(n26138), .Y(n73520) );
  NAND2X1 U62241 ( .A(u_csr_csr_medeleg_q[3]), .B(opcode_instr_w_39), .Y(
        n28529) );
  NAND2X1 U62242 ( .A(n28531), .B(opcode_instr_w_38), .Y(n28530) );
  INVX1 U62243 ( .A(n971), .Y(n28524) );
  NAND2X1 U62244 ( .A(n73543), .B(n73418), .Y(n58247) );
  NOR2X1 U62245 ( .A(n58252), .B(n58247), .Y(n28245) );
  NOR2X1 U62246 ( .A(n73539), .B(n58213), .Y(n28241) );
  INVX1 U62247 ( .A(n28234), .Y(n73575) );
  NOR2X1 U62248 ( .A(n58248), .B(n58277), .Y(n28228) );
  NAND2X1 U62249 ( .A(n26138), .B(n73420), .Y(n58214) );
  NAND2X1 U62250 ( .A(n58278), .B(n58214), .Y(n58215) );
  NAND2X1 U62251 ( .A(n42559), .B(n58215), .Y(n28225) );
  NOR2X1 U62252 ( .A(n28034), .B(n58249), .Y(n28224) );
  INVX1 U62253 ( .A(n58252), .Y(n58477) );
  NAND2X1 U62254 ( .A(n58477), .B(n42962), .Y(n25083) );
  NOR2X1 U62255 ( .A(n58248), .B(n58343), .Y(n28205) );
  NAND2X1 U62256 ( .A(n28202), .B(n26138), .Y(n58217) );
  NAND2X1 U62257 ( .A(n58217), .B(n58216), .Y(n58219) );
  NAND2X1 U62258 ( .A(n58219), .B(n58218), .Y(n58220) );
  NAND2X1 U62259 ( .A(n1887), .B(n58220), .Y(n26971) );
  NOR2X1 U62260 ( .A(n58248), .B(n58408), .Y(n28178) );
  NAND2X1 U62261 ( .A(n26957), .B(n73518), .Y(n58221) );
  NAND2X1 U62262 ( .A(n42951), .B(n58221), .Y(n28172) );
  NOR2X1 U62263 ( .A(n58248), .B(n58423), .Y(n28164) );
  NAND2X1 U62264 ( .A(n58278), .B(n26138), .Y(n58223) );
  NAND2X1 U62265 ( .A(n466), .B(opcode_instr_w_38), .Y(n58224) );
  OR2X1 U62266 ( .A(n28034), .B(n58224), .Y(n28163) );
  NOR2X1 U62267 ( .A(opcode_instr_w_39), .B(n28163), .Y(n28155) );
  INVX1 U62268 ( .A(n58248), .Y(n58478) );
  NAND2X1 U62269 ( .A(n58478), .B(n73173), .Y(n58225) );
  NOR2X1 U62270 ( .A(n44060), .B(n58225), .Y(n28151) );
  NOR2X1 U62271 ( .A(n44060), .B(n58230), .Y(n58226) );
  NOR2X1 U62272 ( .A(n73575), .B(n58226), .Y(n28149) );
  INVX1 U62273 ( .A(n58227), .Y(n73172) );
  INVX1 U62274 ( .A(n27401), .Y(n73401) );
  INVX1 U62275 ( .A(n58228), .Y(n73167) );
  NOR2X1 U62276 ( .A(n73167), .B(n73539), .Y(n28098) );
  NAND2X1 U62277 ( .A(n58229), .B(n58451), .Y(n28091) );
  NAND2X1 U62278 ( .A(n43004), .B(n58230), .Y(n27342) );
  NAND2X1 U62279 ( .A(n58229), .B(n73509), .Y(n28070) );
  NAND2X1 U62280 ( .A(n58229), .B(n58452), .Y(n28067) );
  NAND2X1 U62281 ( .A(n58229), .B(n58453), .Y(n28064) );
  NAND2X1 U62282 ( .A(n58229), .B(n58454), .Y(n28059) );
  NAND2X1 U62283 ( .A(n43002), .B(n39945), .Y(n58238) );
  NAND2X1 U62284 ( .A(n28045), .B(n58238), .Y(n28058) );
  NAND2X1 U62285 ( .A(n73173), .B(n39938), .Y(n58267) );
  INVX1 U62286 ( .A(n58267), .Y(n58240) );
  NAND2X1 U62287 ( .A(n58229), .B(n58240), .Y(n28056) );
  NAND2X1 U62288 ( .A(n58229), .B(n73503), .Y(n24958) );
  INVX1 U62289 ( .A(n24958), .Y(n73399) );
  NAND2X1 U62290 ( .A(n44282), .B(n58230), .Y(n26258) );
  NOR2X1 U62291 ( .A(n73172), .B(n73399), .Y(n27465) );
  NAND2X1 U62292 ( .A(n42323), .B(n58451), .Y(n27461) );
  NAND2X1 U62293 ( .A(n42323), .B(n73509), .Y(n27434) );
  NAND2X1 U62294 ( .A(n42323), .B(n58452), .Y(n27431) );
  NAND2X1 U62295 ( .A(n42323), .B(n58453), .Y(n27428) );
  NAND2X1 U62296 ( .A(n42323), .B(n58454), .Y(n27423) );
  NAND2X1 U62297 ( .A(n27407), .B(n58238), .Y(n27422) );
  NAND2X1 U62298 ( .A(n42323), .B(n58240), .Y(n27420) );
  INVX1 U62299 ( .A(n26261), .Y(n887) );
  NAND2X1 U62300 ( .A(n43003), .B(n43967), .Y(n73158) );
  NAND2X1 U62301 ( .A(n27381), .B(n73158), .Y(n27398) );
  NAND2X1 U62302 ( .A(n73173), .B(n38825), .Y(n58237) );
  INVX1 U62303 ( .A(n58237), .Y(n58232) );
  NOR2X1 U62304 ( .A(n24942), .B(n43969), .Y(n58231) );
  NAND2X1 U62305 ( .A(n58232), .B(n58231), .Y(n27395) );
  NAND2X1 U62306 ( .A(n58233), .B(n42306), .Y(n27385) );
  NAND2X1 U62307 ( .A(n27377), .B(n58238), .Y(n27384) );
  NAND2X1 U62308 ( .A(n73402), .B(n58240), .Y(n27382) );
  NAND2X1 U62309 ( .A(n43004), .B(n38387), .Y(n73142) );
  NAND2X1 U62310 ( .A(n27381), .B(n73142), .Y(n27380) );
  NAND2X1 U62311 ( .A(n58233), .B(n42142), .Y(n27379) );
  NAND2X1 U62312 ( .A(n43002), .B(n43855), .Y(n73134) );
  NAND2X1 U62313 ( .A(n27377), .B(n73134), .Y(n27376) );
  NOR2X1 U62314 ( .A(n889), .B(n58234), .Y(n58235) );
  NAND2X1 U62315 ( .A(n43850), .B(n58235), .Y(n27374) );
  NAND2X1 U62316 ( .A(n27353), .B(n73158), .Y(n27364) );
  NAND2X1 U62317 ( .A(n43962), .B(n58243), .Y(n58236) );
  NOR2X1 U62318 ( .A(n58237), .B(n58236), .Y(n27361) );
  NAND2X1 U62319 ( .A(n58243), .B(n42306), .Y(n27349) );
  INVX1 U62320 ( .A(n27342), .Y(n58241) );
  INVX1 U62321 ( .A(n58238), .Y(n58239) );
  NOR2X1 U62322 ( .A(n58241), .B(n58239), .Y(n27346) );
  NAND2X1 U62323 ( .A(n73403), .B(n58240), .Y(n27343) );
  INVX1 U62324 ( .A(n73142), .Y(n58242) );
  NOR2X1 U62325 ( .A(n58242), .B(n58241), .Y(n27339) );
  NAND2X1 U62326 ( .A(n58243), .B(n42142), .Y(n27336) );
  INVX1 U62327 ( .A(n73134), .Y(n58244) );
  NOR2X1 U62328 ( .A(n27332), .B(n58244), .Y(n27331) );
  NAND2X1 U62329 ( .A(n73173), .B(n73403), .Y(n58245) );
  NOR2X1 U62330 ( .A(n43855), .B(n58245), .Y(n27329) );
  NOR2X1 U62331 ( .A(n37663), .B(opcode_opcode_w[29]), .Y(n27322) );
  NOR2X1 U62332 ( .A(n73367), .B(n37688), .Y(n27323) );
  INVX1 U62333 ( .A(n26270), .Y(n58256) );
  INVX1 U62334 ( .A(n58246), .Y(n73514) );
  NAND2X1 U62335 ( .A(n73167), .B(n58451), .Y(n27306) );
  NAND2X1 U62336 ( .A(n73167), .B(n73509), .Y(n27272) );
  NAND2X1 U62337 ( .A(n73167), .B(n58452), .Y(n27239) );
  NAND2X1 U62338 ( .A(n73167), .B(n58453), .Y(n27230) );
  NAND2X1 U62339 ( .A(n73167), .B(n58454), .Y(n27226) );
  NAND2X1 U62340 ( .A(n73172), .B(n58451), .Y(n27205) );
  NAND2X1 U62341 ( .A(n73172), .B(n73509), .Y(n27168) );
  NAND2X1 U62342 ( .A(n73172), .B(n58452), .Y(n27135) );
  NAND2X1 U62343 ( .A(n73172), .B(n58453), .Y(n27126) );
  NAND2X1 U62344 ( .A(n73172), .B(n58454), .Y(n27122) );
  NAND2X1 U62345 ( .A(n73167), .B(n42962), .Y(n26912) );
  NOR2X1 U62346 ( .A(n58248), .B(n58247), .Y(n26995) );
  NOR2X1 U62347 ( .A(n58252), .B(n58277), .Y(n26990) );
  NOR2X1 U62348 ( .A(u_csr_N3161), .B(opcode_instr_w_39), .Y(n26988) );
  INVX1 U62349 ( .A(n28225), .Y(n26986) );
  NOR2X1 U62350 ( .A(n58252), .B(n58343), .Y(n26979) );
  NOR2X1 U62351 ( .A(n26951), .B(n58249), .Y(n26980) );
  NOR2X1 U62352 ( .A(n58252), .B(n58408), .Y(n26961) );
  NAND2X1 U62353 ( .A(n26957), .B(n73508), .Y(n58250) );
  NAND2X1 U62354 ( .A(n42955), .B(n58250), .Y(n26955) );
  NOR2X1 U62355 ( .A(opcode_instr_w_39), .B(n26951), .Y(n26949) );
  NOR2X1 U62356 ( .A(n58252), .B(n58423), .Y(n26941) );
  NAND2X1 U62357 ( .A(n58477), .B(n73173), .Y(n58253) );
  NOR2X1 U62358 ( .A(n44060), .B(n58253), .Y(n26937) );
  NAND2X1 U62359 ( .A(n73506), .B(n58254), .Y(n58425) );
  INVX1 U62360 ( .A(n58425), .Y(n58283) );
  NAND2X1 U62361 ( .A(n58283), .B(n42962), .Y(n58275) );
  INVX1 U62362 ( .A(n58255), .Y(n72834) );
  NAND2X1 U62363 ( .A(n58266), .B(n73173), .Y(n73003) );
  NOR2X1 U62364 ( .A(n43967), .B(n73003), .Y(n58261) );
  INVX1 U62365 ( .A(n58257), .Y(n58258) );
  NOR2X1 U62366 ( .A(n26304), .B(n58258), .Y(n58259) );
  NOR2X1 U62367 ( .A(n58259), .B(n37688), .Y(n58260) );
  NOR2X1 U62368 ( .A(n58261), .B(n58260), .Y(n26306) );
  NOR2X1 U62369 ( .A(n43958), .B(n73003), .Y(n58265) );
  NOR2X1 U62370 ( .A(n43953), .B(n42444), .Y(n58262) );
  NOR2X1 U62371 ( .A(n26304), .B(n58262), .Y(n58263) );
  NOR2X1 U62372 ( .A(n37749), .B(n58263), .Y(n58264) );
  NOR2X1 U62373 ( .A(n58265), .B(n58264), .Y(n26298) );
  NAND2X1 U62374 ( .A(n58266), .B(n58453), .Y(n26290) );
  NOR2X1 U62375 ( .A(n887), .B(n58267), .Y(n26286) );
  NAND2X1 U62376 ( .A(n26270), .B(n58268), .Y(n26281) );
  NAND2X1 U62377 ( .A(n26270), .B(n58269), .Y(n26266) );
  NOR2X1 U62378 ( .A(n38387), .B(n73003), .Y(n58271) );
  NOR2X1 U62379 ( .A(n37748), .B(n73514), .Y(n58270) );
  NOR2X1 U62380 ( .A(n58271), .B(n58270), .Y(n26262) );
  NAND2X1 U62381 ( .A(n26258), .B(n58272), .Y(n26257) );
  NAND2X1 U62382 ( .A(n73173), .B(n44038), .Y(n58273) );
  NOR2X1 U62383 ( .A(n887), .B(n58273), .Y(n26253) );
  NAND2X1 U62384 ( .A(n58275), .B(n58274), .Y(n72833) );
  NAND2X1 U62385 ( .A(n42327), .B(n58451), .Y(n26244) );
  NAND2X1 U62386 ( .A(n42327), .B(n73509), .Y(n26206) );
  NAND2X1 U62387 ( .A(n42327), .B(n58452), .Y(n26173) );
  NAND2X1 U62388 ( .A(n42327), .B(n58453), .Y(n26164) );
  NAND2X1 U62389 ( .A(n42327), .B(n58454), .Y(n26159) );
  NOR2X1 U62390 ( .A(n1858), .B(n43395), .Y(n26139) );
  NOR2X1 U62391 ( .A(n58425), .B(n58277), .Y(n26140) );
  NAND2X1 U62392 ( .A(u_csr_N184), .B(n36766), .Y(n26123) );
  NOR2X1 U62393 ( .A(n1857), .B(n43392), .Y(n26121) );
  NOR2X1 U62394 ( .A(n2350), .B(n43392), .Y(n26117) );
  NOR2X1 U62395 ( .A(n2351), .B(n43395), .Y(n26118) );
  NOR2X1 U62396 ( .A(n58280), .B(n43398), .Y(n26109) );
  NAND2X1 U62397 ( .A(n44075), .B(n43866), .Y(n58281) );
  NAND2X1 U62398 ( .A(n44285), .B(n58281), .Y(n58282) );
  NAND2X1 U62399 ( .A(u_csr_csr_stval_q[10]), .B(n58282), .Y(n58285) );
  NAND2X1 U62400 ( .A(n42138), .B(n43862), .Y(n58284) );
  NAND2X1 U62401 ( .A(n58285), .B(n58284), .Y(n26110) );
  NOR2X1 U62402 ( .A(n2251), .B(n43392), .Y(n26105) );
  NOR2X1 U62403 ( .A(n2252), .B(n43395), .Y(n26106) );
  NOR2X1 U62404 ( .A(n58286), .B(n43398), .Y(n26099) );
  NAND2X1 U62405 ( .A(n44075), .B(n43967), .Y(n58287) );
  NAND2X1 U62406 ( .A(n44285), .B(n58287), .Y(n58288) );
  NAND2X1 U62407 ( .A(u_csr_csr_stval_q[11]), .B(n58288), .Y(n58290) );
  NAND2X1 U62408 ( .A(n42138), .B(n43965), .Y(n58289) );
  NAND2X1 U62409 ( .A(n58290), .B(n58289), .Y(n26100) );
  NOR2X1 U62410 ( .A(n58291), .B(n43398), .Y(n26089) );
  NAND2X1 U62411 ( .A(n44075), .B(n43957), .Y(n58292) );
  NAND2X1 U62412 ( .A(n44285), .B(n58292), .Y(n58293) );
  NAND2X1 U62413 ( .A(u_csr_csr_stval_q[12]), .B(n58293), .Y(n58295) );
  NAND2X1 U62414 ( .A(n42138), .B(n43955), .Y(n58294) );
  NAND2X1 U62415 ( .A(n58295), .B(n58294), .Y(n26090) );
  NOR2X1 U62416 ( .A(n2683), .B(n43395), .Y(n58297) );
  NOR2X1 U62417 ( .A(n8296), .B(n43392), .Y(n58296) );
  NOR2X1 U62418 ( .A(n58297), .B(n58296), .Y(n26087) );
  NOR2X1 U62419 ( .A(n58298), .B(n43398), .Y(n26079) );
  NAND2X1 U62420 ( .A(n44075), .B(n43874), .Y(n58299) );
  NAND2X1 U62421 ( .A(n44284), .B(n58299), .Y(n58300) );
  NAND2X1 U62422 ( .A(u_csr_csr_stval_q[13]), .B(n58300), .Y(n58302) );
  NAND2X1 U62423 ( .A(n43402), .B(n43872), .Y(n58301) );
  NAND2X1 U62424 ( .A(n58302), .B(n58301), .Y(n26080) );
  NOR2X1 U62425 ( .A(n2753), .B(n43395), .Y(n58304) );
  NOR2X1 U62426 ( .A(n8298), .B(n43392), .Y(n58303) );
  NOR2X1 U62427 ( .A(n58304), .B(n58303), .Y(n26077) );
  NOR2X1 U62428 ( .A(n58305), .B(n43398), .Y(n26069) );
  NAND2X1 U62429 ( .A(n44075), .B(n43885), .Y(n58306) );
  NAND2X1 U62430 ( .A(n44284), .B(n58306), .Y(n58307) );
  NAND2X1 U62431 ( .A(u_csr_csr_stval_q[14]), .B(n58307), .Y(n58309) );
  NAND2X1 U62432 ( .A(n43402), .B(n43882), .Y(n58308) );
  NAND2X1 U62433 ( .A(n58309), .B(n58308), .Y(n26070) );
  NOR2X1 U62434 ( .A(n1797), .B(n43395), .Y(n58311) );
  NOR2X1 U62435 ( .A(n8300), .B(n43392), .Y(n58310) );
  NOR2X1 U62436 ( .A(n58311), .B(n58310), .Y(n26067) );
  NOR2X1 U62437 ( .A(n58312), .B(n43398), .Y(n26059) );
  NAND2X1 U62438 ( .A(n44075), .B(n43895), .Y(n58313) );
  NAND2X1 U62439 ( .A(n44284), .B(n58313), .Y(n58314) );
  NAND2X1 U62440 ( .A(u_csr_csr_stval_q[15]), .B(n58314), .Y(n58316) );
  NAND2X1 U62441 ( .A(n43402), .B(n43892), .Y(n58315) );
  NAND2X1 U62442 ( .A(n58316), .B(n58315), .Y(n26060) );
  NOR2X1 U62443 ( .A(n1869), .B(n43395), .Y(n58318) );
  NOR2X1 U62444 ( .A(n8302), .B(n43392), .Y(n58317) );
  NOR2X1 U62445 ( .A(n58318), .B(n58317), .Y(n26057) );
  NOR2X1 U62446 ( .A(n8304), .B(n43392), .Y(n26055) );
  NOR2X1 U62447 ( .A(n2516), .B(n43395), .Y(n26056) );
  NOR2X1 U62448 ( .A(n58319), .B(n43398), .Y(n26049) );
  NAND2X1 U62449 ( .A(n44075), .B(n43901), .Y(n58320) );
  NAND2X1 U62450 ( .A(n44284), .B(n58320), .Y(n58321) );
  NAND2X1 U62451 ( .A(u_csr_csr_stval_q[16]), .B(n58321), .Y(n58323) );
  NAND2X1 U62452 ( .A(n43402), .B(n43898), .Y(n58322) );
  NAND2X1 U62453 ( .A(n58323), .B(n58322), .Y(n26050) );
  NOR2X1 U62454 ( .A(n58324), .B(n43398), .Y(n26039) );
  NAND2X1 U62455 ( .A(n44075), .B(n43908), .Y(n58325) );
  NAND2X1 U62456 ( .A(n44284), .B(n58325), .Y(n58326) );
  NAND2X1 U62457 ( .A(u_csr_csr_stval_q[17]), .B(n58326), .Y(n58328) );
  NAND2X1 U62458 ( .A(n43402), .B(n43906), .Y(n58327) );
  NAND2X1 U62459 ( .A(n58328), .B(n58327), .Y(n26040) );
  NOR2X1 U62460 ( .A(n2882), .B(n43395), .Y(n58330) );
  NOR2X1 U62461 ( .A(n8306), .B(n43392), .Y(n58329) );
  NOR2X1 U62462 ( .A(n58330), .B(n58329), .Y(n26037) );
  NOR2X1 U62463 ( .A(n58331), .B(n43398), .Y(n26029) );
  NAND2X1 U62464 ( .A(n44075), .B(n43915), .Y(n58332) );
  NAND2X1 U62465 ( .A(n44284), .B(n58332), .Y(n58333) );
  NAND2X1 U62466 ( .A(u_csr_csr_stval_q[18]), .B(n58333), .Y(n58335) );
  NAND2X1 U62467 ( .A(n43402), .B(n43911), .Y(n58334) );
  NAND2X1 U62468 ( .A(n58335), .B(n58334), .Y(n26030) );
  NOR2X1 U62469 ( .A(n2650), .B(n43395), .Y(n58337) );
  NOR2X1 U62470 ( .A(n8308), .B(n43392), .Y(n58336) );
  NOR2X1 U62471 ( .A(n58337), .B(n58336), .Y(n26027) );
  NOR2X1 U62472 ( .A(n8310), .B(n43392), .Y(n26025) );
  NOR2X1 U62473 ( .A(n2283), .B(n43395), .Y(n26026) );
  NOR2X1 U62474 ( .A(n58338), .B(n43398), .Y(n26019) );
  NAND2X1 U62475 ( .A(n44075), .B(n43923), .Y(n58339) );
  NAND2X1 U62476 ( .A(n44284), .B(n58339), .Y(n58340) );
  NAND2X1 U62477 ( .A(u_csr_csr_stval_q[19]), .B(n58340), .Y(n58342) );
  NAND2X1 U62478 ( .A(n43402), .B(n43920), .Y(n58341) );
  NAND2X1 U62479 ( .A(n58342), .B(n58341), .Y(n26020) );
  NOR2X1 U62480 ( .A(n1860), .B(n43395), .Y(n26015) );
  NOR2X1 U62481 ( .A(n58425), .B(n58343), .Y(n26016) );
  NAND2X1 U62482 ( .A(opcode_pc_w[1]), .B(n36766), .Y(n26010) );
  NOR2X1 U62483 ( .A(n1859), .B(n43392), .Y(n26008) );
  NOR2X1 U62484 ( .A(n8314), .B(n43393), .Y(n26004) );
  NOR2X1 U62485 ( .A(n2383), .B(n43396), .Y(n26005) );
  NOR2X1 U62486 ( .A(n58344), .B(n43398), .Y(n25998) );
  NAND2X1 U62487 ( .A(n44075), .B(n43931), .Y(n58345) );
  NAND2X1 U62488 ( .A(n44284), .B(n58345), .Y(n58346) );
  NAND2X1 U62489 ( .A(u_csr_csr_stval_q[20]), .B(n58346), .Y(n58348) );
  NAND2X1 U62490 ( .A(n43402), .B(n43929), .Y(n58347) );
  NAND2X1 U62491 ( .A(n58348), .B(n58347), .Y(n25999) );
  NOR2X1 U62492 ( .A(n58349), .B(n43398), .Y(n25988) );
  NAND2X1 U62493 ( .A(n44075), .B(n43939), .Y(n58350) );
  NAND2X1 U62494 ( .A(n44284), .B(n58350), .Y(n58351) );
  NAND2X1 U62495 ( .A(u_csr_csr_stval_q[21]), .B(n58351), .Y(n58353) );
  NAND2X1 U62496 ( .A(n43402), .B(n43936), .Y(n58352) );
  NAND2X1 U62497 ( .A(n58353), .B(n58352), .Y(n25989) );
  NOR2X1 U62498 ( .A(n2549), .B(n43396), .Y(n58355) );
  NOR2X1 U62499 ( .A(n8316), .B(n43393), .Y(n58354) );
  NOR2X1 U62500 ( .A(n58355), .B(n58354), .Y(n25986) );
  NOR2X1 U62501 ( .A(n58356), .B(n43399), .Y(n25978) );
  NAND2X1 U62502 ( .A(n44076), .B(n43948), .Y(n58357) );
  NAND2X1 U62503 ( .A(n44284), .B(n58357), .Y(n58358) );
  NAND2X1 U62504 ( .A(u_csr_csr_stval_q[22]), .B(n58358), .Y(n58360) );
  NAND2X1 U62505 ( .A(n43402), .B(n43945), .Y(n58359) );
  NAND2X1 U62506 ( .A(n58360), .B(n58359), .Y(n25979) );
  NOR2X1 U62507 ( .A(n2483), .B(n43396), .Y(n58362) );
  NOR2X1 U62508 ( .A(n8318), .B(n43393), .Y(n58361) );
  NOR2X1 U62509 ( .A(n58362), .B(n58361), .Y(n25976) );
  NOR2X1 U62510 ( .A(n58363), .B(n43399), .Y(n25968) );
  NAND2X1 U62511 ( .A(n44076), .B(n43978), .Y(n58364) );
  NAND2X1 U62512 ( .A(n44284), .B(n58364), .Y(n58365) );
  NAND2X1 U62513 ( .A(u_csr_csr_stval_q[23]), .B(n58365), .Y(n58367) );
  NAND2X1 U62514 ( .A(n43402), .B(n43975), .Y(n58366) );
  NAND2X1 U62515 ( .A(n58367), .B(n58366), .Y(n25969) );
  NOR2X1 U62516 ( .A(n2451), .B(n43396), .Y(n58369) );
  NOR2X1 U62517 ( .A(n8320), .B(n43393), .Y(n58368) );
  NOR2X1 U62518 ( .A(n58369), .B(n58368), .Y(n25966) );
  NOR2X1 U62519 ( .A(n58370), .B(n43399), .Y(n25958) );
  NAND2X1 U62520 ( .A(n44076), .B(n43988), .Y(n58371) );
  NAND2X1 U62521 ( .A(n44284), .B(n58371), .Y(n58372) );
  NAND2X1 U62522 ( .A(u_csr_csr_stval_q[24]), .B(n58372), .Y(n58374) );
  NAND2X1 U62523 ( .A(n43402), .B(n43985), .Y(n58373) );
  NAND2X1 U62524 ( .A(n58374), .B(n58373), .Y(n25959) );
  NOR2X1 U62525 ( .A(n2850), .B(n43396), .Y(n58376) );
  NOR2X1 U62526 ( .A(n8322), .B(n43393), .Y(n58375) );
  NOR2X1 U62527 ( .A(n58376), .B(n58375), .Y(n25956) );
  NOR2X1 U62528 ( .A(n8324), .B(n43393), .Y(n25954) );
  NOR2X1 U62529 ( .A(n2817), .B(n43396), .Y(n25955) );
  NOR2X1 U62530 ( .A(n58377), .B(n43399), .Y(n25948) );
  NAND2X1 U62531 ( .A(n44076), .B(n43996), .Y(n58378) );
  NAND2X1 U62532 ( .A(n44283), .B(n58378), .Y(n58379) );
  NAND2X1 U62533 ( .A(u_csr_csr_stval_q[25]), .B(n58379), .Y(n58381) );
  NAND2X1 U62534 ( .A(n43401), .B(n43994), .Y(n58380) );
  NAND2X1 U62535 ( .A(n58381), .B(n58380), .Y(n25949) );
  NOR2X1 U62536 ( .A(n58382), .B(n43399), .Y(n25938) );
  NAND2X1 U62537 ( .A(n44076), .B(n44006), .Y(n58383) );
  NAND2X1 U62538 ( .A(n44283), .B(n58383), .Y(n58384) );
  NAND2X1 U62539 ( .A(u_csr_csr_stval_q[26]), .B(n58384), .Y(n58386) );
  NAND2X1 U62540 ( .A(n43401), .B(n44002), .Y(n58385) );
  NAND2X1 U62541 ( .A(n58386), .B(n58385), .Y(n25939) );
  NOR2X1 U62542 ( .A(n2617), .B(n43396), .Y(n58388) );
  NOR2X1 U62543 ( .A(n8326), .B(n43393), .Y(n58387) );
  NOR2X1 U62544 ( .A(n58388), .B(n58387), .Y(n25936) );
  NOR2X1 U62545 ( .A(n58389), .B(n43399), .Y(n25928) );
  NAND2X1 U62546 ( .A(n44076), .B(n44012), .Y(n58390) );
  NAND2X1 U62547 ( .A(n44283), .B(n58390), .Y(n58391) );
  NAND2X1 U62548 ( .A(u_csr_csr_stval_q[27]), .B(n58391), .Y(n58393) );
  NAND2X1 U62549 ( .A(n43401), .B(n44010), .Y(n58392) );
  NAND2X1 U62550 ( .A(n58393), .B(n58392), .Y(n25929) );
  NOR2X1 U62551 ( .A(n2785), .B(n43396), .Y(n58395) );
  NOR2X1 U62552 ( .A(n8328), .B(n43393), .Y(n58394) );
  NOR2X1 U62553 ( .A(n58395), .B(n58394), .Y(n25926) );
  NOR2X1 U62554 ( .A(n58396), .B(n43399), .Y(n25918) );
  NAND2X1 U62555 ( .A(n44076), .B(n44021), .Y(n58397) );
  NAND2X1 U62556 ( .A(n44283), .B(n58397), .Y(n58398) );
  NAND2X1 U62557 ( .A(u_csr_csr_stval_q[28]), .B(n58398), .Y(n58400) );
  NAND2X1 U62558 ( .A(n43401), .B(n44019), .Y(n58399) );
  NAND2X1 U62559 ( .A(n58400), .B(n58399), .Y(n25919) );
  NOR2X1 U62560 ( .A(n1870), .B(n43396), .Y(n58402) );
  NOR2X1 U62561 ( .A(n8330), .B(n43393), .Y(n58401) );
  NOR2X1 U62562 ( .A(n58402), .B(n58401), .Y(n25916) );
  NOR2X1 U62563 ( .A(n8332), .B(n43393), .Y(n25914) );
  NOR2X1 U62564 ( .A(n1801), .B(n43396), .Y(n25915) );
  NOR2X1 U62565 ( .A(n58403), .B(n43399), .Y(n25908) );
  NAND2X1 U62566 ( .A(n44076), .B(n44028), .Y(n58404) );
  NAND2X1 U62567 ( .A(n44283), .B(n58404), .Y(n58405) );
  NAND2X1 U62568 ( .A(u_csr_csr_stval_q[29]), .B(n58405), .Y(n58407) );
  NAND2X1 U62569 ( .A(n43401), .B(n44027), .Y(n58406) );
  NAND2X1 U62570 ( .A(n58407), .B(n58406), .Y(n25909) );
  NOR2X1 U62571 ( .A(n1862), .B(n43396), .Y(n25904) );
  NOR2X1 U62572 ( .A(n58425), .B(n58408), .Y(n25905) );
  NAND2X1 U62573 ( .A(opcode_pc_w[2]), .B(n36766), .Y(n25899) );
  NOR2X1 U62574 ( .A(n1861), .B(n43393), .Y(n25897) );
  NOR2X1 U62575 ( .A(n58409), .B(n43399), .Y(n25887) );
  NAND2X1 U62576 ( .A(n44076), .B(n44053), .Y(n58410) );
  NAND2X1 U62577 ( .A(n44283), .B(n58410), .Y(n58411) );
  NAND2X1 U62578 ( .A(u_csr_csr_stval_q[30]), .B(n58411), .Y(n58413) );
  NAND2X1 U62579 ( .A(n43401), .B(n44050), .Y(n58412) );
  NAND2X1 U62580 ( .A(n58413), .B(n58412), .Y(n25888) );
  NOR2X1 U62581 ( .A(n1871), .B(n43396), .Y(n58415) );
  NOR2X1 U62582 ( .A(n8336), .B(n43393), .Y(n58414) );
  NOR2X1 U62583 ( .A(n58415), .B(n58414), .Y(n25885) );
  NOR2X1 U62584 ( .A(n58416), .B(n43399), .Y(n25877) );
  NAND2X1 U62585 ( .A(n44076), .B(n44060), .Y(n58417) );
  NAND2X1 U62586 ( .A(n44283), .B(n58417), .Y(n58418) );
  NAND2X1 U62587 ( .A(u_csr_csr_stval_q[31]), .B(n58418), .Y(n58420) );
  NAND2X1 U62588 ( .A(n43401), .B(n44057), .Y(n58419) );
  NAND2X1 U62589 ( .A(n58420), .B(n58419), .Y(n25878) );
  NOR2X1 U62590 ( .A(n1872), .B(n43397), .Y(n58422) );
  NOR2X1 U62591 ( .A(n8338), .B(n43394), .Y(n58421) );
  NOR2X1 U62592 ( .A(n58422), .B(n58421), .Y(n25875) );
  NOR2X1 U62593 ( .A(n1864), .B(n43397), .Y(n25873) );
  NOR2X1 U62594 ( .A(n58425), .B(n58423), .Y(n25874) );
  NAND2X1 U62595 ( .A(opcode_pc_w[3]), .B(n36766), .Y(n25868) );
  NOR2X1 U62596 ( .A(n1863), .B(n43394), .Y(n25866) );
  NOR2X1 U62597 ( .A(n1866), .B(n43397), .Y(n25861) );
  NOR2X1 U62598 ( .A(n58425), .B(n58424), .Y(n25862) );
  NAND2X1 U62599 ( .A(opcode_pc_w[4]), .B(n36766), .Y(n25855) );
  NOR2X1 U62600 ( .A(n1865), .B(n43394), .Y(n25853) );
  NOR2X1 U62601 ( .A(n1867), .B(n43394), .Y(n25849) );
  NOR2X1 U62602 ( .A(n1868), .B(n43397), .Y(n25850) );
  NOR2X1 U62603 ( .A(n58426), .B(n43399), .Y(n25843) );
  NAND2X1 U62604 ( .A(n44076), .B(n39944), .Y(n58427) );
  NAND2X1 U62605 ( .A(n44283), .B(n58427), .Y(n58428) );
  NAND2X1 U62606 ( .A(u_csr_csr_stval_q[5]), .B(n58428), .Y(n58430) );
  NAND2X1 U62607 ( .A(n43401), .B(n39939), .Y(n58429) );
  NAND2X1 U62608 ( .A(n58430), .B(n58429), .Y(n25844) );
  NOR2X1 U62609 ( .A(n2316), .B(n43394), .Y(n25839) );
  NOR2X1 U62610 ( .A(n2317), .B(n43397), .Y(n25840) );
  NOR2X1 U62611 ( .A(n58431), .B(n43399), .Y(n25833) );
  NAND2X1 U62612 ( .A(n44076), .B(n43847), .Y(n58432) );
  NAND2X1 U62613 ( .A(n44283), .B(n58432), .Y(n58433) );
  NAND2X1 U62614 ( .A(u_csr_csr_stval_q[6]), .B(n58433), .Y(n58435) );
  NAND2X1 U62615 ( .A(n43401), .B(n43843), .Y(n58434) );
  NAND2X1 U62616 ( .A(n58435), .B(n58434), .Y(n25834) );
  NOR2X1 U62617 ( .A(n2581), .B(n43394), .Y(n25829) );
  NOR2X1 U62618 ( .A(n2582), .B(n43397), .Y(n25830) );
  NOR2X1 U62619 ( .A(n58436), .B(n43400), .Y(n25823) );
  NAND2X1 U62620 ( .A(n42210), .B(n38386), .Y(n58437) );
  NAND2X1 U62621 ( .A(n44283), .B(n58437), .Y(n58438) );
  NAND2X1 U62622 ( .A(u_csr_csr_stval_q[7]), .B(n58438), .Y(n58440) );
  NAND2X1 U62623 ( .A(n43401), .B(n38382), .Y(n58439) );
  NAND2X1 U62624 ( .A(n58440), .B(n58439), .Y(n25824) );
  NOR2X1 U62625 ( .A(n2716), .B(n43394), .Y(n25819) );
  NOR2X1 U62626 ( .A(n2717), .B(n43397), .Y(n25820) );
  NOR2X1 U62627 ( .A(n58441), .B(n43400), .Y(n25813) );
  NAND2X1 U62628 ( .A(n42210), .B(n44040), .Y(n58442) );
  NAND2X1 U62629 ( .A(n44283), .B(n58442), .Y(n58443) );
  NAND2X1 U62630 ( .A(u_csr_csr_stval_q[8]), .B(n58443), .Y(n58445) );
  NAND2X1 U62631 ( .A(n43401), .B(n44038), .Y(n58444) );
  NAND2X1 U62632 ( .A(n58445), .B(n58444), .Y(n25814) );
  NOR2X1 U62633 ( .A(n2419), .B(n43394), .Y(n25807) );
  NOR2X1 U62634 ( .A(n2420), .B(n43397), .Y(n25808) );
  NOR2X1 U62635 ( .A(n58446), .B(n43400), .Y(n25797) );
  NAND2X1 U62636 ( .A(n42210), .B(n43855), .Y(n58447) );
  NAND2X1 U62637 ( .A(n44283), .B(n58447), .Y(n58448) );
  NAND2X1 U62638 ( .A(u_csr_csr_stval_q[9]), .B(n58448), .Y(n58450) );
  NAND2X1 U62639 ( .A(n43401), .B(n43853), .Y(n58449) );
  NAND2X1 U62640 ( .A(n58450), .B(n58449), .Y(n25798) );
  NAND2X1 U62641 ( .A(n72834), .B(n58451), .Y(n25788) );
  NAND2X1 U62642 ( .A(n72834), .B(n73509), .Y(n25741) );
  NAND2X1 U62643 ( .A(n72834), .B(n58452), .Y(n25696) );
  NAND2X1 U62644 ( .A(n72834), .B(n58453), .Y(n25683) );
  NAND2X1 U62645 ( .A(n72834), .B(n58454), .Y(n25677) );
  NOR2X1 U62646 ( .A(n42966), .B(n58455), .Y(n25652) );
  NOR2X1 U62647 ( .A(n42963), .B(n58456), .Y(n25647) );
  NAND2X1 U62648 ( .A(n73367), .B(n58457), .Y(n25639) );
  NAND2X1 U62649 ( .A(n58818), .B(n73364), .Y(n25640) );
  OR2X1 U62650 ( .A(n42747), .B(n25635), .Y(n58460) );
  NAND2X1 U62651 ( .A(n38501), .B(n73503), .Y(n58459) );
  NOR2X1 U62652 ( .A(n58460), .B(n58459), .Y(n25637) );
  NAND2X1 U62653 ( .A(n38824), .B(n42962), .Y(n58501) );
  NOR2X1 U62654 ( .A(n25635), .B(n58501), .Y(n25631) );
  NAND2X1 U62655 ( .A(n42748), .B(opcode_opcode_w[29]), .Y(n58461) );
  NOR2X1 U62656 ( .A(n58462), .B(n58461), .Y(n25632) );
  NOR2X1 U62657 ( .A(n42967), .B(n58463), .Y(n25613) );
  NOR2X1 U62658 ( .A(n42964), .B(n58464), .Y(n25609) );
  NOR2X1 U62659 ( .A(n42965), .B(n58465), .Y(n25588) );
  NOR2X1 U62660 ( .A(n42963), .B(n58466), .Y(n25583) );
  NOR2X1 U62661 ( .A(n25574), .B(n58501), .Y(n25572) );
  INVX1 U62662 ( .A(n58467), .Y(n73500) );
  INVX1 U62663 ( .A(n58468), .Y(n73502) );
  OR2X1 U62664 ( .A(n24877), .B(n38464), .Y(n58470) );
  NOR2X1 U62665 ( .A(n24942), .B(n58470), .Y(n24910) );
  INVX1 U62666 ( .A(n58471), .Y(n73498) );
  INVX1 U62667 ( .A(n58472), .Y(n73499) );
  INVX1 U62668 ( .A(n58473), .Y(n73496) );
  INVX1 U62669 ( .A(n58474), .Y(n73497) );
  NOR2X1 U62670 ( .A(n42966), .B(n58475), .Y(n25378) );
  NOR2X1 U62671 ( .A(n42963), .B(n58476), .Y(n25373) );
  NAND2X1 U62672 ( .A(u_csr_csr_scause_q[1]), .B(n58477), .Y(n25364) );
  NAND2X1 U62673 ( .A(u_csr_csr_mcause_q[1]), .B(n58478), .Y(n25361) );
  NOR2X1 U62674 ( .A(n42967), .B(n58479), .Y(n25304) );
  NAND2X1 U62675 ( .A(u_csr_csr_mepc_q[22]), .B(n42131), .Y(n25300) );
  NOR2X1 U62676 ( .A(n42965), .B(n58480), .Y(n25284) );
  NAND2X1 U62677 ( .A(u_csr_csr_mepc_q[23]), .B(n42131), .Y(n25280) );
  NOR2X1 U62678 ( .A(n42966), .B(n58481), .Y(n25264) );
  NAND2X1 U62679 ( .A(u_csr_csr_mepc_q[24]), .B(n42131), .Y(n25260) );
  NOR2X1 U62680 ( .A(n42967), .B(n58482), .Y(n25244) );
  NAND2X1 U62681 ( .A(u_csr_csr_mepc_q[25]), .B(n42131), .Y(n25240) );
  NOR2X1 U62682 ( .A(n42965), .B(n58483), .Y(n25224) );
  NAND2X1 U62683 ( .A(u_csr_csr_mepc_q[26]), .B(n42131), .Y(n25220) );
  NOR2X1 U62684 ( .A(n42966), .B(n58484), .Y(n25204) );
  NAND2X1 U62685 ( .A(u_csr_csr_mepc_q[27]), .B(n42131), .Y(n25200) );
  NOR2X1 U62686 ( .A(n42967), .B(n58485), .Y(n25184) );
  NAND2X1 U62687 ( .A(u_csr_csr_mepc_q[28]), .B(n42131), .Y(n25180) );
  NOR2X1 U62688 ( .A(n42965), .B(n58486), .Y(n25164) );
  NAND2X1 U62689 ( .A(u_csr_csr_mepc_q[29]), .B(n42131), .Y(n25160) );
  NOR2X1 U62690 ( .A(n42966), .B(n58487), .Y(n25142) );
  NOR2X1 U62691 ( .A(n42964), .B(n58488), .Y(n25137) );
  NAND2X1 U62692 ( .A(u_csr_csr_sepc_q[30]), .B(n73501), .Y(n25114) );
  NOR2X1 U62693 ( .A(n42963), .B(n58489), .Y(n25112) );
  NAND2X1 U62694 ( .A(u_csr_csr_sepc_q[31]), .B(n73501), .Y(n25093) );
  NOR2X1 U62695 ( .A(n42963), .B(n58490), .Y(n25091) );
  INVX1 U62696 ( .A(n25083), .Y(n73400) );
  NOR2X1 U62697 ( .A(n42967), .B(n58491), .Y(n25069) );
  NOR2X1 U62698 ( .A(n42964), .B(n58492), .Y(n25062) );
  NOR2X1 U62699 ( .A(n25051), .B(n58501), .Y(n25049) );
  NOR2X1 U62700 ( .A(n42965), .B(n58493), .Y(n25035) );
  NOR2X1 U62701 ( .A(n42963), .B(n58494), .Y(n25031) );
  NOR2X1 U62702 ( .A(n42966), .B(n58495), .Y(n25010) );
  NOR2X1 U62703 ( .A(n42963), .B(n58496), .Y(n25005) );
  NOR2X1 U62704 ( .A(n42967), .B(n58497), .Y(n24982) );
  NOR2X1 U62705 ( .A(n42964), .B(n58498), .Y(n24978) );
  NOR2X1 U62706 ( .A(n42965), .B(n58499), .Y(n24955) );
  NOR2X1 U62707 ( .A(n42963), .B(n58500), .Y(n24950) );
  NOR2X1 U62708 ( .A(n24938), .B(n58501), .Y(n24936) );
  NOR2X1 U62709 ( .A(n42966), .B(n58502), .Y(n24923) );
  NOR2X1 U62710 ( .A(n42963), .B(n58503), .Y(n24918) );
  NOR2X1 U62711 ( .A(n42967), .B(n58504), .Y(n24895) );
  NOR2X1 U62712 ( .A(n42964), .B(n58505), .Y(n24889) );
  NAND2X1 U62713 ( .A(mem_i_inst_i[0]), .B(n43319), .Y(n58507) );
  NAND2X1 U62714 ( .A(n58510), .B(n58507), .Y(net2336) );
  NAND2X1 U62715 ( .A(u_fetch_skid_buffer_q[0]), .B(n43406), .Y(n24855) );
  INVX1 U62716 ( .A(mem_i_inst_i[2]), .Y(n58508) );
  NOR2X1 U62717 ( .A(n43404), .B(n58508), .Y(net2339) );
  NAND2X1 U62718 ( .A(u_fetch_skid_buffer_q[2]), .B(n43406), .Y(n24852) );
  NAND2X1 U62719 ( .A(mem_i_inst_i[1]), .B(n43319), .Y(n58509) );
  NAND2X1 U62720 ( .A(n58510), .B(n58509), .Y(net2337) );
  NAND2X1 U62721 ( .A(u_fetch_skid_buffer_q[1]), .B(n43407), .Y(n24850) );
  NAND2X1 U62722 ( .A(n58512), .B(n8801), .Y(n24504) );
  NOR2X1 U62723 ( .A(n24464), .B(n58513), .Y(n24462) );
  INVX1 U62724 ( .A(n58514), .Y(n73541) );
  INVX1 U62725 ( .A(n24436), .Y(n602) );
  INVX1 U62726 ( .A(n24422), .Y(n73530) );
  INVX1 U62727 ( .A(n58515), .Y(n73515) );
  NOR2X1 U62728 ( .A(n24539), .B(n24535), .Y(n58516) );
  NAND2X1 U62729 ( .A(n37568), .B(n58516), .Y(n73389) );
  INVX1 U62730 ( .A(n73389), .Y(n73398) );
  INVX1 U62731 ( .A(n58517), .Y(n73531) );
  INVX1 U62732 ( .A(n58518), .Y(n24237) );
  INVX1 U62733 ( .A(n58519), .Y(n73423) );
  NOR2X1 U62734 ( .A(u_csr_writeback_idx_q[1]), .B(n37537), .Y(n24337) );
  INVX1 U62735 ( .A(n58520), .Y(n73426) );
  NOR2X1 U62736 ( .A(opcode_opcode_w[8]), .B(opcode_opcode_w[9]), .Y(n58522)
         );
  NAND2X1 U62737 ( .A(n58522), .B(n58521), .Y(n58536) );
  NOR2X1 U62738 ( .A(n58523), .B(n58536), .Y(n58524) );
  NOR2X1 U62739 ( .A(n24306), .B(n58524), .Y(n24299) );
  NOR2X1 U62740 ( .A(n24237), .B(n37537), .Y(n24295) );
  NOR2X1 U62741 ( .A(n58525), .B(n58536), .Y(n58526) );
  NOR2X1 U62742 ( .A(n24298), .B(n58526), .Y(n24291) );
  INVX1 U62743 ( .A(n58536), .Y(n58532) );
  NAND2X1 U62744 ( .A(n58532), .B(n58527), .Y(n58528) );
  NAND2X1 U62745 ( .A(n24275), .B(n58528), .Y(n24273) );
  INVX1 U62746 ( .A(n24180), .Y(n73424) );
  NOR2X1 U62747 ( .A(n58529), .B(n58536), .Y(n58530) );
  NOR2X1 U62748 ( .A(n24239), .B(n58530), .Y(n24232) );
  NAND2X1 U62749 ( .A(n58532), .B(n58531), .Y(n58533) );
  NAND2X1 U62750 ( .A(n24229), .B(n58533), .Y(n24227) );
  INVX1 U62751 ( .A(n24135), .Y(n73422) );
  NOR2X1 U62752 ( .A(n58534), .B(n58536), .Y(n58535) );
  NOR2X1 U62753 ( .A(n24125), .B(n58535), .Y(n24119) );
  NOR2X1 U62754 ( .A(n58537), .B(n58536), .Y(n58538) );
  NOR2X1 U62755 ( .A(n24117), .B(n58538), .Y(n24112) );
  INVX1 U62756 ( .A(n24217), .Y(n552) );
  INVX1 U62757 ( .A(n24203), .Y(n549) );
  INVX1 U62758 ( .A(n24188), .Y(n73425) );
  INVX1 U62759 ( .A(n24170), .Y(n567) );
  INVX1 U62760 ( .A(n24336), .Y(n497) );
  INVX1 U62761 ( .A(n24328), .Y(n503) );
  INVX1 U62762 ( .A(n24316), .Y(n495) );
  INVX1 U62763 ( .A(n24283), .Y(n559) );
  INVX1 U62764 ( .A(n24263), .Y(n555) );
  INVX1 U62765 ( .A(n24247), .Y(n563) );
  NAND2X1 U62766 ( .A(n42949), .B(n15977), .Y(n16922) );
  INVX1 U62767 ( .A(n16922), .Y(n17949) );
  NAND2X1 U62768 ( .A(n43420), .B(n15805), .Y(n17944) );
  NAND2X1 U62769 ( .A(n43424), .B(n16042), .Y(n16566) );
  INVX1 U62770 ( .A(n15594), .Y(n73524) );
  INVX1 U62771 ( .A(n15410), .Y(n73572) );
  INVX1 U62772 ( .A(n15498), .Y(n58542) );
  NAND2X1 U62773 ( .A(n43420), .B(n58542), .Y(n358) );
  NOR2X1 U62774 ( .A(n1890), .B(n58539), .Y(n17900) );
  NAND2X1 U62775 ( .A(n58541), .B(n58540), .Y(n17899) );
  NAND2X1 U62776 ( .A(n42947), .B(n58542), .Y(n360) );
  NOR2X1 U62777 ( .A(n73448), .B(n43414), .Y(n17868) );
  NOR2X1 U62778 ( .A(n73450), .B(n40690), .Y(n17869) );
  NOR2X1 U62779 ( .A(n73452), .B(n43422), .Y(n17858) );
  NOR2X1 U62780 ( .A(n73446), .B(n43417), .Y(n17859) );
  NAND2X1 U62781 ( .A(n42948), .B(n16563), .Y(n16708) );
  INVX1 U62782 ( .A(n16708), .Y(n17845) );
  NOR2X1 U62783 ( .A(n73468), .B(n43422), .Y(n17835) );
  NOR2X1 U62784 ( .A(n73462), .B(n43417), .Y(n17836) );
  NOR2X1 U62785 ( .A(n73456), .B(n43414), .Y(n17824) );
  NOR2X1 U62786 ( .A(n73460), .B(n43422), .Y(n17814) );
  NOR2X1 U62787 ( .A(n73454), .B(n43417), .Y(n17815) );
  INVX1 U62788 ( .A(n15737), .Y(n73432) );
  NAND2X1 U62789 ( .A(n58542), .B(n43425), .Y(n17796) );
  NOR2X1 U62790 ( .A(n58544), .B(n58543), .Y(n58545) );
  NAND2X1 U62791 ( .A(n58545), .B(n73513), .Y(n16080) );
  NOR2X1 U62792 ( .A(n73439), .B(n43414), .Y(n17781) );
  NOR2X1 U62793 ( .A(n73438), .B(n43417), .Y(n17782) );
  NOR2X1 U62794 ( .A(n73444), .B(n43421), .Y(n17770) );
  NOR2X1 U62795 ( .A(n73442), .B(n40690), .Y(n17771) );
  NAND2X1 U62796 ( .A(n43736), .B(n39164), .Y(n58546) );
  NOR2X1 U62797 ( .A(n43412), .B(n58546), .Y(n58550) );
  NAND2X1 U62798 ( .A(opcode_opcode_w[27]), .B(opcode_opcode_w[28]), .Y(n58547) );
  NOR2X1 U62799 ( .A(n58548), .B(n58547), .Y(n58549) );
  NOR2X1 U62800 ( .A(n58550), .B(n58549), .Y(n17578) );
  NAND2X1 U62801 ( .A(n58659), .B(n73523), .Y(n58551) );
  NAND2X1 U62802 ( .A(n58551), .B(n73492), .Y(n58553) );
  NAND2X1 U62803 ( .A(n42435), .B(n58577), .Y(n58552) );
  NAND2X1 U62804 ( .A(n58553), .B(n58552), .Y(n17572) );
  NOR2X1 U62805 ( .A(n73364), .B(n58817), .Y(n58555) );
  NAND2X1 U62806 ( .A(n58555), .B(n58554), .Y(n58559) );
  NOR2X1 U62807 ( .A(n43746), .B(n43793), .Y(n58557) );
  NAND2X1 U62808 ( .A(n58557), .B(n43410), .Y(n58558) );
  NAND2X1 U62809 ( .A(n58559), .B(n58558), .Y(n17551) );
  INVX1 U62810 ( .A(n58561), .Y(n58562) );
  NAND2X1 U62811 ( .A(n58562), .B(n43759), .Y(n58564) );
  NAND2X1 U62812 ( .A(n17203), .B(n73482), .Y(n58563) );
  NAND2X1 U62813 ( .A(n58564), .B(n58563), .Y(n17531) );
  NAND2X1 U62814 ( .A(n43419), .B(n15728), .Y(n17427) );
  NAND2X1 U62815 ( .A(n43424), .B(n15447), .Y(n16817) );
  NOR2X1 U62816 ( .A(n73460), .B(n43414), .Y(n17416) );
  NOR2X1 U62817 ( .A(n73458), .B(n43417), .Y(n17417) );
  NOR2X1 U62818 ( .A(n73464), .B(n43421), .Y(n17415) );
  NOR2X1 U62819 ( .A(n58577), .B(n43414), .Y(n58566) );
  NOR2X1 U62820 ( .A(n73491), .B(n43421), .Y(n58565) );
  NOR2X1 U62821 ( .A(n58566), .B(n58565), .Y(n58568) );
  NAND2X1 U62822 ( .A(n42949), .B(n16596), .Y(n58567) );
  NAND2X1 U62823 ( .A(n58568), .B(n58567), .Y(n16182) );
  INVX1 U62824 ( .A(n16182), .Y(n73397) );
  NOR2X1 U62825 ( .A(n73448), .B(n43422), .Y(n17404) );
  NOR2X1 U62826 ( .A(n73446), .B(n40690), .Y(n17405) );
  NOR2X1 U62827 ( .A(n73444), .B(n43414), .Y(n17402) );
  NOR2X1 U62828 ( .A(n73442), .B(n43417), .Y(n17403) );
  NOR2X1 U62829 ( .A(n73488), .B(n40690), .Y(n17399) );
  NOR2X1 U62830 ( .A(n73495), .B(n43417), .Y(n17397) );
  NOR2X1 U62831 ( .A(n73490), .B(n43414), .Y(n17398) );
  NOR2X1 U62832 ( .A(n73452), .B(n43414), .Y(n17388) );
  NOR2X1 U62833 ( .A(n73456), .B(n43422), .Y(n17386) );
  NOR2X1 U62834 ( .A(n73450), .B(n43417), .Y(n17387) );
  NAND2X1 U62835 ( .A(n73492), .B(n58658), .Y(n17376) );
  INVX1 U62836 ( .A(n58658), .Y(n58654) );
  NAND2X1 U62837 ( .A(n58654), .B(n16596), .Y(n58569) );
  NAND2X1 U62838 ( .A(n17375), .B(n58569), .Y(n15932) );
  NAND2X1 U62839 ( .A(n17156), .B(n43429), .Y(n58571) );
  OR2X1 U62840 ( .A(n43437), .B(n58573), .Y(n58570) );
  NAND2X1 U62841 ( .A(n58571), .B(n58570), .Y(n17340) );
  INVX1 U62842 ( .A(n58759), .Y(n58807) );
  NOR2X1 U62843 ( .A(n17156), .B(n43431), .Y(n58572) );
  NOR2X1 U62844 ( .A(n43441), .B(n58572), .Y(n58575) );
  NAND2X1 U62845 ( .A(n43432), .B(n58573), .Y(n58574) );
  NAND2X1 U62846 ( .A(n42451), .B(n16775), .Y(n17331) );
  NAND2X1 U62847 ( .A(n42948), .B(n15805), .Y(n16815) );
  NAND2X1 U62848 ( .A(n43420), .B(n16563), .Y(n16562) );
  NAND2X1 U62849 ( .A(n42949), .B(n58580), .Y(n17326) );
  NAND2X1 U62850 ( .A(n42316), .B(n15862), .Y(n17327) );
  NAND2X1 U62851 ( .A(n43420), .B(n58576), .Y(n363) );
  NOR2X1 U62852 ( .A(n73439), .B(n43417), .Y(n17192) );
  NOR2X1 U62853 ( .A(n73446), .B(n43421), .Y(n17193) );
  NOR2X1 U62854 ( .A(n73444), .B(n40691), .Y(n17190) );
  NOR2X1 U62855 ( .A(n73442), .B(n43414), .Y(n17191) );
  NOR2X1 U62856 ( .A(n73491), .B(n40689), .Y(n17182) );
  NOR2X1 U62857 ( .A(n73495), .B(n43422), .Y(n17183) );
  NOR2X1 U62858 ( .A(n58577), .B(n43417), .Y(n58579) );
  NOR2X1 U62859 ( .A(n73492), .B(n43414), .Y(n58578) );
  NOR2X1 U62860 ( .A(n58579), .B(n58578), .Y(n17180) );
  NOR2X1 U62861 ( .A(n73486), .B(n40691), .Y(n17178) );
  NOR2X1 U62862 ( .A(n73484), .B(n43421), .Y(n17179) );
  NOR2X1 U62863 ( .A(n73490), .B(n43417), .Y(n17176) );
  NOR2X1 U62864 ( .A(n73488), .B(n43414), .Y(n17177) );
  NAND2X1 U62865 ( .A(n43424), .B(n58580), .Y(n15530) );
  NAND2X1 U62866 ( .A(n42947), .B(n16775), .Y(n16774) );
  NAND2X1 U62867 ( .A(n42451), .B(n16563), .Y(n16668) );
  NAND2X1 U62868 ( .A(n43425), .B(n15805), .Y(n17159) );
  NAND2X1 U62869 ( .A(n17083), .B(n43429), .Y(n58583) );
  INVX1 U62870 ( .A(n58581), .Y(n58584) );
  NAND2X1 U62871 ( .A(n58584), .B(n43433), .Y(n58582) );
  NOR2X1 U62872 ( .A(n58584), .B(n43436), .Y(n58585) );
  NOR2X1 U62873 ( .A(n58807), .B(n58585), .Y(n58588) );
  INVX1 U62874 ( .A(n17083), .Y(n58586) );
  NAND2X1 U62875 ( .A(n43427), .B(n58586), .Y(n58587) );
  NAND2X1 U62876 ( .A(n58588), .B(n58587), .Y(n17143) );
  NAND2X1 U62877 ( .A(n42948), .B(n16042), .Y(n17028) );
  INVX1 U62878 ( .A(n17028), .Y(n17131) );
  NAND2X1 U62879 ( .A(n43420), .B(n15846), .Y(n17130) );
  NOR2X1 U62880 ( .A(n73448), .B(n43418), .Y(n17127) );
  NOR2X1 U62881 ( .A(n73450), .B(n43414), .Y(n17128) );
  NOR2X1 U62882 ( .A(n73454), .B(n43423), .Y(n17125) );
  NOR2X1 U62883 ( .A(n73452), .B(n40689), .Y(n17126) );
  NOR2X1 U62884 ( .A(n73456), .B(n43418), .Y(n17119) );
  NOR2X1 U62885 ( .A(n73458), .B(n43414), .Y(n17120) );
  NOR2X1 U62886 ( .A(n73462), .B(n43423), .Y(n17118) );
  NOR2X1 U62887 ( .A(n73486), .B(n43413), .Y(n17095) );
  NAND2X1 U62888 ( .A(n17094), .B(n43420), .Y(n17093) );
  NOR2X1 U62889 ( .A(n73490), .B(n43423), .Y(n17090) );
  NOR2X1 U62890 ( .A(n73492), .B(n43416), .Y(n17091) );
  NOR2X1 U62891 ( .A(n73491), .B(n43413), .Y(n17088) );
  NOR2X1 U62892 ( .A(n73495), .B(n40689), .Y(n17089) );
  NAND2X1 U62893 ( .A(n17018), .B(n43428), .Y(n58591) );
  INVX1 U62894 ( .A(n58589), .Y(n58592) );
  NAND2X1 U62895 ( .A(n58592), .B(n43433), .Y(n58590) );
  NOR2X1 U62896 ( .A(n58592), .B(n43435), .Y(n58593) );
  NOR2X1 U62897 ( .A(n58807), .B(n58593), .Y(n58596) );
  INVX1 U62898 ( .A(n17018), .Y(n58594) );
  NAND2X1 U62899 ( .A(n43427), .B(n58594), .Y(n58595) );
  NAND2X1 U62900 ( .A(n58596), .B(n58595), .Y(n17070) );
  NOR2X1 U62901 ( .A(n73482), .B(n43418), .Y(n17058) );
  NAND2X1 U62902 ( .A(n42948), .B(n15728), .Y(n17057) );
  NAND2X1 U62903 ( .A(n43425), .B(n73511), .Y(n15672) );
  NAND2X1 U62904 ( .A(n43425), .B(n16596), .Y(n58599) );
  NAND2X1 U62905 ( .A(n42949), .B(n58597), .Y(n58598) );
  NOR2X1 U62906 ( .A(n73466), .B(n43423), .Y(n17043) );
  NOR2X1 U62907 ( .A(n73460), .B(n43416), .Y(n17044) );
  NOR2X1 U62908 ( .A(n73462), .B(n43413), .Y(n17042) );
  NOR2X1 U62909 ( .A(n73494), .B(n40691), .Y(n17036) );
  NOR2X1 U62910 ( .A(n73482), .B(n43423), .Y(n17037) );
  NOR2X1 U62911 ( .A(n73486), .B(n43416), .Y(n17034) );
  NOR2X1 U62912 ( .A(n73484), .B(n43413), .Y(n17035) );
  NOR2X1 U62913 ( .A(n73480), .B(n43418), .Y(n17029) );
  NAND2X1 U62914 ( .A(n43419), .B(n16775), .Y(n17025) );
  NAND2X1 U62915 ( .A(n16953), .B(n43428), .Y(n58602) );
  INVX1 U62916 ( .A(n58600), .Y(n58603) );
  NAND2X1 U62917 ( .A(n58603), .B(n43433), .Y(n58601) );
  NOR2X1 U62918 ( .A(n58603), .B(n43436), .Y(n58604) );
  NOR2X1 U62919 ( .A(n58807), .B(n58604), .Y(n58607) );
  INVX1 U62920 ( .A(n16953), .Y(n58605) );
  NAND2X1 U62921 ( .A(n43427), .B(n58605), .Y(n58606) );
  NAND2X1 U62922 ( .A(n58607), .B(n58606), .Y(n17004) );
  NOR2X1 U62923 ( .A(n73446), .B(n43413), .Y(n16994) );
  NOR2X1 U62924 ( .A(n73448), .B(n40691), .Y(n16995) );
  NOR2X1 U62925 ( .A(n73444), .B(n43418), .Y(n16992) );
  NOR2X1 U62926 ( .A(n73450), .B(n43423), .Y(n16993) );
  NOR2X1 U62927 ( .A(n73458), .B(n43423), .Y(n16986) );
  NOR2X1 U62928 ( .A(n73452), .B(n43416), .Y(n16987) );
  NOR2X1 U62929 ( .A(n73439), .B(n40690), .Y(n16982) );
  NOR2X1 U62930 ( .A(n73438), .B(n43413), .Y(n16983) );
  NAND2X1 U62931 ( .A(n17322), .B(n42455), .Y(n15887) );
  NOR2X1 U62932 ( .A(n15887), .B(n43416), .Y(n16980) );
  NOR2X1 U62933 ( .A(n73442), .B(n43423), .Y(n16981) );
  NOR2X1 U62934 ( .A(n73490), .B(n40689), .Y(n16974) );
  NOR2X1 U62935 ( .A(n73488), .B(n43423), .Y(n16975) );
  NOR2X1 U62936 ( .A(n73491), .B(n43418), .Y(n16972) );
  NOR2X1 U62937 ( .A(n73495), .B(n43413), .Y(n16973) );
  OR2X1 U62938 ( .A(n43439), .B(n58611), .Y(n58609) );
  NAND2X1 U62939 ( .A(n16892), .B(n43428), .Y(n58608) );
  NAND2X1 U62940 ( .A(n58609), .B(n58608), .Y(n16937) );
  NOR2X1 U62941 ( .A(n16892), .B(n43431), .Y(n58610) );
  NOR2X1 U62942 ( .A(n58807), .B(n58610), .Y(n58613) );
  NAND2X1 U62943 ( .A(n43432), .B(n58611), .Y(n58612) );
  INVX1 U62944 ( .A(n361), .Y(n15416) );
  NOR2X1 U62945 ( .A(n73484), .B(n43416), .Y(n16926) );
  NOR2X1 U62946 ( .A(n73494), .B(n43413), .Y(n16927) );
  INVX1 U62947 ( .A(n17427), .Y(n16923) );
  NAND2X1 U62948 ( .A(n43424), .B(n15728), .Y(n15727) );
  INVX1 U62949 ( .A(n15727), .Y(n16899) );
  NOR2X1 U62950 ( .A(n73494), .B(n43418), .Y(n16897) );
  NOR2X1 U62951 ( .A(n73482), .B(n43413), .Y(n16898) );
  INVX1 U62952 ( .A(n15530), .Y(n73396) );
  NAND2X1 U62953 ( .A(n16845), .B(n43428), .Y(n58616) );
  INVX1 U62954 ( .A(n58614), .Y(n58617) );
  NAND2X1 U62955 ( .A(n58617), .B(n43433), .Y(n58615) );
  NOR2X1 U62956 ( .A(n58617), .B(n43437), .Y(n58618) );
  NOR2X1 U62957 ( .A(n58807), .B(n58618), .Y(n58621) );
  INVX1 U62958 ( .A(n16845), .Y(n58619) );
  NAND2X1 U62959 ( .A(n43427), .B(n58619), .Y(n58620) );
  NAND2X1 U62960 ( .A(n58621), .B(n58620), .Y(n16878) );
  INVX1 U62961 ( .A(n58622), .Y(n58627) );
  NOR2X1 U62962 ( .A(n58627), .B(n43436), .Y(n58623) );
  NOR2X1 U62963 ( .A(n43441), .B(n58623), .Y(n58626) );
  INVX1 U62964 ( .A(n16793), .Y(n58624) );
  NAND2X1 U62965 ( .A(n43427), .B(n58624), .Y(n58625) );
  NAND2X1 U62966 ( .A(n58626), .B(n58625), .Y(n16826) );
  NAND2X1 U62967 ( .A(n16793), .B(n43427), .Y(n58629) );
  NAND2X1 U62968 ( .A(n58627), .B(n43433), .Y(n58628) );
  NAND2X1 U62969 ( .A(n16342), .B(n42310), .Y(n15965) );
  NOR2X1 U62970 ( .A(n15965), .B(n58734), .Y(n16829) );
  INVX1 U62971 ( .A(n58630), .Y(n58635) );
  NOR2X1 U62972 ( .A(n58635), .B(n43436), .Y(n58631) );
  NOR2X1 U62973 ( .A(n58807), .B(n58631), .Y(n58634) );
  INVX1 U62974 ( .A(n16740), .Y(n58632) );
  NAND2X1 U62975 ( .A(n43427), .B(n58632), .Y(n58633) );
  NAND2X1 U62976 ( .A(n58634), .B(n58633), .Y(n16769) );
  NAND2X1 U62977 ( .A(n16740), .B(n43428), .Y(n58637) );
  NAND2X1 U62978 ( .A(n58635), .B(n43433), .Y(n58636) );
  INVX1 U62979 ( .A(n17130), .Y(n16776) );
  INVX1 U62980 ( .A(n58638), .Y(n58643) );
  NOR2X1 U62981 ( .A(n58643), .B(n43437), .Y(n58639) );
  NOR2X1 U62982 ( .A(n43442), .B(n58639), .Y(n58642) );
  INVX1 U62983 ( .A(n16686), .Y(n58640) );
  NAND2X1 U62984 ( .A(n43427), .B(n58640), .Y(n58641) );
  NAND2X1 U62985 ( .A(n58642), .B(n58641), .Y(n16719) );
  NAND2X1 U62986 ( .A(n16686), .B(n43428), .Y(n58645) );
  NAND2X1 U62987 ( .A(n58643), .B(n43434), .Y(n58644) );
  INVX1 U62988 ( .A(n17944), .Y(n16709) );
  INVX1 U62989 ( .A(n17331), .Y(n16710) );
  INVX1 U62990 ( .A(n58646), .Y(n58651) );
  NOR2X1 U62991 ( .A(n58651), .B(n43435), .Y(n58647) );
  NOR2X1 U62992 ( .A(n43442), .B(n58647), .Y(n58650) );
  INVX1 U62993 ( .A(n16558), .Y(n58648) );
  NAND2X1 U62994 ( .A(n43426), .B(n58648), .Y(n58649) );
  NAND2X1 U62995 ( .A(n58650), .B(n58649), .Y(n16663) );
  NAND2X1 U62996 ( .A(n16558), .B(n43427), .Y(n58653) );
  NAND2X1 U62997 ( .A(n58651), .B(n43434), .Y(n58652) );
  INVX1 U62998 ( .A(n17025), .Y(n16669) );
  INVX1 U62999 ( .A(n17159), .Y(n16656) );
  NAND2X1 U63000 ( .A(n43419), .B(n16042), .Y(n16637) );
  INVX1 U63001 ( .A(n16637), .Y(n16653) );
  NAND2X1 U63002 ( .A(n43424), .B(n15977), .Y(n16507) );
  NOR2X1 U63003 ( .A(n58654), .B(n43431), .Y(n58655) );
  NOR2X1 U63004 ( .A(n43442), .B(n58655), .Y(n58657) );
  NAND2X1 U63005 ( .A(n43432), .B(n58659), .Y(n58656) );
  NAND2X1 U63006 ( .A(n58657), .B(n58656), .Y(n16597) );
  NOR2X1 U63007 ( .A(n58805), .B(n58658), .Y(n58661) );
  NOR2X1 U63008 ( .A(n43436), .B(n58659), .Y(n58660) );
  NOR2X1 U63009 ( .A(n58661), .B(n58660), .Y(n16598) );
  NOR2X1 U63010 ( .A(n16599), .B(n43423), .Y(n16590) );
  NAND2X1 U63011 ( .A(n16505), .B(n43427), .Y(n58664) );
  INVX1 U63012 ( .A(n58662), .Y(n58665) );
  NAND2X1 U63013 ( .A(n58665), .B(n43434), .Y(n58663) );
  NOR2X1 U63014 ( .A(n58665), .B(n43438), .Y(n58666) );
  NOR2X1 U63015 ( .A(n43442), .B(n58666), .Y(n58669) );
  INVX1 U63016 ( .A(n16505), .Y(n58667) );
  NAND2X1 U63017 ( .A(n43426), .B(n58667), .Y(n58668) );
  NAND2X1 U63018 ( .A(n58669), .B(n58668), .Y(n16544) );
  NAND2X1 U63019 ( .A(n42310), .B(n73432), .Y(n15966) );
  NOR2X1 U63020 ( .A(n15966), .B(n58734), .Y(n16529) );
  INVX1 U63021 ( .A(n58670), .Y(n58673) );
  NAND2X1 U63022 ( .A(n58673), .B(n43434), .Y(n58672) );
  NAND2X1 U63023 ( .A(n16451), .B(n43427), .Y(n58671) );
  NAND2X1 U63024 ( .A(n58672), .B(n58671), .Y(n16488) );
  NOR2X1 U63025 ( .A(n58673), .B(n43439), .Y(n58674) );
  NOR2X1 U63026 ( .A(n43442), .B(n58674), .Y(n58677) );
  INVX1 U63027 ( .A(n16451), .Y(n58675) );
  NAND2X1 U63028 ( .A(n43426), .B(n58675), .Y(n58676) );
  NAND2X1 U63029 ( .A(n58677), .B(n58676), .Y(n16489) );
  INVX1 U63030 ( .A(n364), .Y(n73510) );
  INVX1 U63031 ( .A(n15672), .Y(n73395) );
  NAND2X1 U63032 ( .A(n43424), .B(n73512), .Y(n16148) );
  INVX1 U63033 ( .A(n58678), .Y(n58681) );
  NAND2X1 U63034 ( .A(n58681), .B(n43434), .Y(n58680) );
  NAND2X1 U63035 ( .A(n16397), .B(n43428), .Y(n58679) );
  NAND2X1 U63036 ( .A(n58680), .B(n58679), .Y(n16433) );
  NOR2X1 U63037 ( .A(n58681), .B(n43439), .Y(n58682) );
  NOR2X1 U63038 ( .A(n43442), .B(n58682), .Y(n58685) );
  INVX1 U63039 ( .A(n16397), .Y(n58683) );
  NAND2X1 U63040 ( .A(n43426), .B(n58683), .Y(n58684) );
  NAND2X1 U63041 ( .A(n58685), .B(n58684), .Y(n16434) );
  INVX1 U63042 ( .A(n58686), .Y(n58689) );
  NAND2X1 U63043 ( .A(n58689), .B(n43433), .Y(n58688) );
  NAND2X1 U63044 ( .A(n16339), .B(n43428), .Y(n58687) );
  NAND2X1 U63045 ( .A(n58688), .B(n58687), .Y(n16380) );
  NOR2X1 U63046 ( .A(n58689), .B(n43438), .Y(n58690) );
  NOR2X1 U63047 ( .A(n43442), .B(n58690), .Y(n58693) );
  INVX1 U63048 ( .A(n16339), .Y(n58691) );
  NAND2X1 U63049 ( .A(n43426), .B(n58691), .Y(n58692) );
  NAND2X1 U63050 ( .A(n58693), .B(n58692), .Y(n16381) );
  NAND2X1 U63051 ( .A(n16342), .B(n42315), .Y(n15829) );
  NOR2X1 U63052 ( .A(n15829), .B(n58734), .Y(n16341) );
  INVX1 U63053 ( .A(n58694), .Y(n58697) );
  NAND2X1 U63054 ( .A(n58697), .B(n43433), .Y(n58696) );
  NAND2X1 U63055 ( .A(n16279), .B(n43428), .Y(n58695) );
  NAND2X1 U63056 ( .A(n58696), .B(n58695), .Y(n16322) );
  NOR2X1 U63057 ( .A(n58697), .B(n43437), .Y(n58698) );
  NOR2X1 U63058 ( .A(n43442), .B(n58698), .Y(n58701) );
  INVX1 U63059 ( .A(n16279), .Y(n58699) );
  NAND2X1 U63060 ( .A(n43426), .B(n58699), .Y(n58700) );
  NAND2X1 U63061 ( .A(n58701), .B(n58700), .Y(n16323) );
  INVX1 U63062 ( .A(n363), .Y(n15442) );
  NAND2X1 U63063 ( .A(n73511), .B(n43420), .Y(n15880) );
  NAND2X1 U63064 ( .A(n73511), .B(n42451), .Y(n16084) );
  INVX1 U63065 ( .A(n58702), .Y(n58707) );
  NOR2X1 U63066 ( .A(n58707), .B(n43438), .Y(n58703) );
  NOR2X1 U63067 ( .A(n43442), .B(n58703), .Y(n58706) );
  INVX1 U63068 ( .A(n16215), .Y(n58704) );
  NAND2X1 U63069 ( .A(n43426), .B(n58704), .Y(n58705) );
  NAND2X1 U63070 ( .A(n58706), .B(n58705), .Y(n16263) );
  NAND2X1 U63071 ( .A(n58707), .B(n43433), .Y(n58709) );
  NAND2X1 U63072 ( .A(n16215), .B(n43429), .Y(n58708) );
  NAND2X1 U63073 ( .A(n58709), .B(n58708), .Y(n16262) );
  INVX1 U63074 ( .A(n58710), .Y(n58715) );
  NOR2X1 U63075 ( .A(n58715), .B(n43439), .Y(n58711) );
  NOR2X1 U63076 ( .A(n43442), .B(n58711), .Y(n58714) );
  INVX1 U63077 ( .A(n16145), .Y(n58712) );
  NAND2X1 U63078 ( .A(n43426), .B(n58712), .Y(n58713) );
  NAND2X1 U63079 ( .A(n58714), .B(n58713), .Y(n16198) );
  NAND2X1 U63080 ( .A(n58715), .B(n43433), .Y(n58717) );
  NAND2X1 U63081 ( .A(n16145), .B(n43428), .Y(n58716) );
  NAND2X1 U63082 ( .A(n58717), .B(n58716), .Y(n16197) );
  NAND2X1 U63083 ( .A(n16009), .B(n43424), .Y(n16178) );
  INVX1 U63084 ( .A(n58718), .Y(n58721) );
  NAND2X1 U63085 ( .A(n58721), .B(n43433), .Y(n58720) );
  NAND2X1 U63086 ( .A(n16079), .B(n43428), .Y(n58719) );
  NAND2X1 U63087 ( .A(n58720), .B(n58719), .Y(n16127) );
  NOR2X1 U63088 ( .A(n58721), .B(n43438), .Y(n58722) );
  NOR2X1 U63089 ( .A(n43442), .B(n58722), .Y(n58725) );
  INVX1 U63090 ( .A(n16079), .Y(n58723) );
  NAND2X1 U63091 ( .A(n43426), .B(n58723), .Y(n58724) );
  NAND2X1 U63092 ( .A(n58725), .B(n58724), .Y(n16128) );
  INVX1 U63093 ( .A(n58726), .Y(n58729) );
  NAND2X1 U63094 ( .A(n58729), .B(n43433), .Y(n58728) );
  NAND2X1 U63095 ( .A(n16005), .B(n43428), .Y(n58727) );
  NAND2X1 U63096 ( .A(n58728), .B(n58727), .Y(n16061) );
  INVX1 U63097 ( .A(n16080), .Y(n981) );
  NOR2X1 U63098 ( .A(n58729), .B(n43436), .Y(n58730) );
  NOR2X1 U63099 ( .A(n43441), .B(n58730), .Y(n58733) );
  INVX1 U63100 ( .A(n16005), .Y(n58731) );
  NAND2X1 U63101 ( .A(n43426), .B(n58731), .Y(n58732) );
  NAND2X1 U63102 ( .A(n58733), .B(n58732), .Y(n16062) );
  NOR2X1 U63103 ( .A(n229), .B(n43423), .Y(n16032) );
  NAND2X1 U63104 ( .A(n42315), .B(n73432), .Y(n15824) );
  NOR2X1 U63105 ( .A(n15824), .B(n58734), .Y(n16033) );
  NOR2X1 U63106 ( .A(n16008), .B(n43418), .Y(n16006) );
  NAND2X1 U63107 ( .A(n15876), .B(n43429), .Y(n58737) );
  INVX1 U63108 ( .A(n58735), .Y(n58738) );
  NAND2X1 U63109 ( .A(n58738), .B(n43433), .Y(n58736) );
  NOR2X1 U63110 ( .A(n58738), .B(n43435), .Y(n58739) );
  NOR2X1 U63111 ( .A(n43441), .B(n58739), .Y(n58742) );
  INVX1 U63112 ( .A(n15876), .Y(n58740) );
  NAND2X1 U63113 ( .A(n43426), .B(n58740), .Y(n58741) );
  NAND2X1 U63114 ( .A(n58742), .B(n58741), .Y(n15990) );
  NOR2X1 U63115 ( .A(n37340), .B(n43423), .Y(n15969) );
  NOR2X1 U63116 ( .A(n229), .B(n40690), .Y(n15970) );
  NOR2X1 U63117 ( .A(n15879), .B(n43413), .Y(n15957) );
  NOR2X1 U63118 ( .A(n15932), .B(n58805), .Y(n58743) );
  NOR2X1 U63119 ( .A(n43441), .B(n58743), .Y(n58745) );
  NAND2X1 U63120 ( .A(n43432), .B(n58746), .Y(n58744) );
  NAND2X1 U63121 ( .A(n58745), .B(n58744), .Y(n15920) );
  NOR2X1 U63122 ( .A(n43437), .B(n58746), .Y(n58749) );
  INVX1 U63123 ( .A(n15932), .Y(n58747) );
  NOR2X1 U63124 ( .A(n58747), .B(n58805), .Y(n58748) );
  NOR2X1 U63125 ( .A(n58749), .B(n58748), .Y(n15921) );
  NAND2X1 U63126 ( .A(n43425), .B(n15846), .Y(n15593) );
  INVX1 U63127 ( .A(n17057), .Y(n15909) );
  NOR2X1 U63128 ( .A(n15879), .B(n43418), .Y(n15878) );
  NAND2X1 U63129 ( .A(n15811), .B(n43429), .Y(n58752) );
  INVX1 U63130 ( .A(n58750), .Y(n58753) );
  NAND2X1 U63131 ( .A(n58753), .B(n43432), .Y(n58751) );
  NOR2X1 U63132 ( .A(n58753), .B(n43439), .Y(n58754) );
  NOR2X1 U63133 ( .A(n43441), .B(n58754), .Y(n58757) );
  INVX1 U63134 ( .A(n15811), .Y(n58755) );
  NAND2X1 U63135 ( .A(n43426), .B(n58755), .Y(n58756) );
  NAND2X1 U63136 ( .A(n58757), .B(n58756), .Y(n15860) );
  NOR2X1 U63137 ( .A(n15784), .B(n43422), .Y(n15837) );
  NOR2X1 U63138 ( .A(n37340), .B(n40691), .Y(n15838) );
  NOR2X1 U63139 ( .A(n229), .B(n43418), .Y(n15822) );
  XNOR2X1 U63140 ( .A(n58760), .B(n15807), .Y(n58758) );
  NOR2X1 U63141 ( .A(n43431), .B(n58758), .Y(n15793) );
  NOR2X1 U63142 ( .A(n15795), .B(n43422), .Y(n15794) );
  NOR2X1 U63143 ( .A(n58760), .B(n58759), .Y(n15782) );
  NOR2X1 U63144 ( .A(n15784), .B(n40689), .Y(n15783) );
  NOR2X1 U63145 ( .A(n15756), .B(n58805), .Y(n58762) );
  NOR2X1 U63146 ( .A(n43441), .B(n58762), .Y(n58764) );
  NAND2X1 U63147 ( .A(n43432), .B(n58765), .Y(n58763) );
  NAND2X1 U63148 ( .A(n58764), .B(n58763), .Y(n15743) );
  NOR2X1 U63149 ( .A(n43435), .B(n58765), .Y(n58768) );
  INVX1 U63150 ( .A(n15756), .Y(n58766) );
  NOR2X1 U63151 ( .A(n58805), .B(n58766), .Y(n58767) );
  NOR2X1 U63152 ( .A(n58768), .B(n58767), .Y(n15744) );
  NOR2X1 U63153 ( .A(n15695), .B(n43431), .Y(n58769) );
  NOR2X1 U63154 ( .A(n43441), .B(n58769), .Y(n58771) );
  NAND2X1 U63155 ( .A(n43432), .B(n58772), .Y(n58770) );
  NAND2X1 U63156 ( .A(n58771), .B(n58770), .Y(n15683) );
  NOR2X1 U63157 ( .A(n43435), .B(n58772), .Y(n58775) );
  INVX1 U63158 ( .A(n15695), .Y(n58773) );
  NOR2X1 U63159 ( .A(n58805), .B(n58773), .Y(n58774) );
  NOR2X1 U63160 ( .A(n58775), .B(n58774), .Y(n15684) );
  NOR2X1 U63161 ( .A(n15641), .B(n58805), .Y(n58776) );
  NOR2X1 U63162 ( .A(n43441), .B(n58776), .Y(n58778) );
  NAND2X1 U63163 ( .A(n43432), .B(n58779), .Y(n58777) );
  NAND2X1 U63164 ( .A(n58778), .B(n58777), .Y(n15632) );
  NAND2X1 U63165 ( .A(n15641), .B(n43429), .Y(n58781) );
  OR2X1 U63166 ( .A(n43435), .B(n58779), .Y(n58780) );
  NAND2X1 U63167 ( .A(n58781), .B(n58780), .Y(n15631) );
  INVX1 U63168 ( .A(n358), .Y(n15600) );
  NAND2X1 U63169 ( .A(n15580), .B(n43429), .Y(n58783) );
  OR2X1 U63170 ( .A(n43438), .B(n58785), .Y(n58782) );
  NAND2X1 U63171 ( .A(n58783), .B(n58782), .Y(n15575) );
  NOR2X1 U63172 ( .A(n15580), .B(n43431), .Y(n58784) );
  NOR2X1 U63173 ( .A(n43441), .B(n58784), .Y(n58787) );
  NAND2X1 U63174 ( .A(n43432), .B(n58785), .Y(n58786) );
  NAND2X1 U63175 ( .A(n58787), .B(n58786), .Y(n15568) );
  INVX1 U63176 ( .A(n15568), .Y(n343) );
  NOR2X1 U63177 ( .A(n15539), .B(n43431), .Y(n58788) );
  NOR2X1 U63178 ( .A(n43441), .B(n58788), .Y(n58790) );
  NAND2X1 U63179 ( .A(n43432), .B(n58791), .Y(n58789) );
  NAND2X1 U63180 ( .A(n58790), .B(n58789), .Y(n15525) );
  NOR2X1 U63181 ( .A(n43435), .B(n58791), .Y(n58794) );
  INVX1 U63182 ( .A(n15539), .Y(n58792) );
  NOR2X1 U63183 ( .A(n58805), .B(n58792), .Y(n58793) );
  NOR2X1 U63184 ( .A(n58794), .B(n58793), .Y(n15526) );
  NAND2X1 U63185 ( .A(n15481), .B(n43429), .Y(n58796) );
  OR2X1 U63186 ( .A(n43436), .B(n58798), .Y(n58795) );
  NAND2X1 U63187 ( .A(n58796), .B(n58795), .Y(n15473) );
  NOR2X1 U63188 ( .A(n15481), .B(n43431), .Y(n58797) );
  NOR2X1 U63189 ( .A(n43441), .B(n58797), .Y(n58800) );
  NAND2X1 U63190 ( .A(n43432), .B(n58798), .Y(n58799) );
  NAND2X1 U63191 ( .A(n15433), .B(n43428), .Y(n58804) );
  OR2X1 U63192 ( .A(n43435), .B(n58808), .Y(n58803) );
  NAND2X1 U63193 ( .A(n58804), .B(n58803), .Y(n15422) );
  NOR2X1 U63194 ( .A(n15433), .B(n43431), .Y(n58806) );
  NOR2X1 U63195 ( .A(n43442), .B(n58806), .Y(n58810) );
  NAND2X1 U63196 ( .A(n43432), .B(n58808), .Y(n58809) );
  NAND2X1 U63197 ( .A(n58812), .B(n58811), .Y(n15319) );
  OR2X1 U63198 ( .A(opcode_instr_w_36), .B(n28943), .Y(n58813) );
  NAND2X1 U63199 ( .A(n73431), .B(n58813), .Y(n58814) );
  NAND2X1 U63200 ( .A(n58815), .B(n58814), .Y(n15320) );
  INVX1 U63201 ( .A(n58816), .Y(n73542) );
  NOR2X1 U63202 ( .A(n58818), .B(n58817), .Y(n58819) );
  NAND2X1 U63203 ( .A(n58819), .B(n43377), .Y(n73366) );
  INVX1 U63204 ( .A(n73366), .Y(n73394) );
  NOR2X1 U63205 ( .A(n73367), .B(n38802), .Y(n58821) );
  NAND2X1 U63206 ( .A(n42760), .B(n58821), .Y(n15220) );
  NAND2X1 U63207 ( .A(n44054), .B(n58822), .Y(n58823) );
  NAND2X1 U63208 ( .A(n58823), .B(n73428), .Y(n73383) );
  INVX1 U63209 ( .A(n73383), .Y(n58970) );
  NAND2X1 U63210 ( .A(n42453), .B(n44057), .Y(n73382) );
  NOR2X1 U63211 ( .A(n73384), .B(n44064), .Y(n58824) );
  NOR2X1 U63212 ( .A(n43443), .B(n58824), .Y(n58826) );
  NAND2X1 U63213 ( .A(n44061), .B(n44070), .Y(n58825) );
  MX2X1 U63214 ( .A(n58826), .B(n58825), .S0(n43461), .Y(n14878) );
  NAND2X1 U63215 ( .A(n36719), .B(n43463), .Y(n58830) );
  NOR2X1 U63216 ( .A(n58830), .B(n44067), .Y(n58827) );
  NOR2X1 U63217 ( .A(n43443), .B(n58827), .Y(n58829) );
  NAND2X1 U63218 ( .A(n44061), .B(n58830), .Y(n58828) );
  MX2X1 U63219 ( .A(n58829), .B(n58828), .S0(n40627), .Y(n14864) );
  INVX1 U63220 ( .A(n58830), .Y(n58831) );
  NAND2X1 U63221 ( .A(n58831), .B(n40627), .Y(n58835) );
  NOR2X1 U63222 ( .A(n58835), .B(n44067), .Y(n58832) );
  NOR2X1 U63223 ( .A(n43443), .B(n58832), .Y(n58834) );
  NAND2X1 U63224 ( .A(n44061), .B(n58835), .Y(n58833) );
  MX2X1 U63225 ( .A(n58834), .B(n58833), .S0(n43475), .Y(n14845) );
  INVX1 U63226 ( .A(n58835), .Y(n58836) );
  NAND2X1 U63227 ( .A(n58836), .B(n43474), .Y(n58840) );
  NOR2X1 U63228 ( .A(n58840), .B(n44067), .Y(n58837) );
  NOR2X1 U63229 ( .A(n43443), .B(n58837), .Y(n58839) );
  NAND2X1 U63230 ( .A(n44061), .B(n58840), .Y(n58838) );
  MX2X1 U63231 ( .A(n58839), .B(n58838), .S0(n43470), .Y(n14831) );
  INVX1 U63232 ( .A(n58840), .Y(n58841) );
  NAND2X1 U63233 ( .A(n58841), .B(n43470), .Y(n58845) );
  NOR2X1 U63234 ( .A(n58845), .B(n44067), .Y(n58842) );
  NOR2X1 U63235 ( .A(n43443), .B(n58842), .Y(n58844) );
  NAND2X1 U63236 ( .A(n44061), .B(n58845), .Y(n58843) );
  MX2X1 U63237 ( .A(n58844), .B(n58843), .S0(n39946), .Y(n14817) );
  INVX1 U63238 ( .A(n58845), .Y(n58846) );
  NAND2X1 U63239 ( .A(n58846), .B(n39944), .Y(n58850) );
  NOR2X1 U63240 ( .A(n58850), .B(n44067), .Y(n58847) );
  NOR2X1 U63241 ( .A(n43443), .B(n58847), .Y(n58849) );
  NAND2X1 U63242 ( .A(n44061), .B(n58850), .Y(n58848) );
  MX2X1 U63243 ( .A(n58849), .B(n58848), .S0(n43846), .Y(n14803) );
  INVX1 U63244 ( .A(n58850), .Y(n58851) );
  NAND2X1 U63245 ( .A(n58851), .B(n43846), .Y(n58855) );
  NOR2X1 U63246 ( .A(n58855), .B(n44066), .Y(n58852) );
  NOR2X1 U63247 ( .A(n43443), .B(n58852), .Y(n58854) );
  NAND2X1 U63248 ( .A(n44061), .B(n58855), .Y(n58853) );
  MX2X1 U63249 ( .A(n58854), .B(n58853), .S0(n38387), .Y(n14789) );
  INVX1 U63250 ( .A(n58855), .Y(n58856) );
  NAND2X1 U63251 ( .A(n58856), .B(n38387), .Y(n58865) );
  NOR2X1 U63252 ( .A(n58865), .B(n44067), .Y(n58857) );
  NOR2X1 U63253 ( .A(n43443), .B(n58857), .Y(n58859) );
  NAND2X1 U63254 ( .A(n44061), .B(n58865), .Y(n58858) );
  MX2X1 U63255 ( .A(n58859), .B(n58858), .S0(n44041), .Y(n14775) );
  INVX1 U63256 ( .A(n58865), .Y(n58860) );
  NAND2X1 U63257 ( .A(n58860), .B(n44040), .Y(n58862) );
  NOR2X1 U63258 ( .A(n44064), .B(n58862), .Y(n58861) );
  NOR2X1 U63259 ( .A(n43443), .B(n58861), .Y(n58864) );
  NAND2X1 U63260 ( .A(n44061), .B(n58862), .Y(n58863) );
  MX2X1 U63261 ( .A(n58864), .B(n58863), .S0(n43856), .Y(n14761) );
  NOR2X1 U63262 ( .A(n43851), .B(n58865), .Y(n58866) );
  NAND2X1 U63263 ( .A(n58866), .B(n44040), .Y(n58870) );
  NOR2X1 U63264 ( .A(n58870), .B(n44066), .Y(n58867) );
  NOR2X1 U63265 ( .A(n43443), .B(n58867), .Y(n58869) );
  NAND2X1 U63266 ( .A(n44061), .B(n58870), .Y(n58868) );
  MX2X1 U63267 ( .A(n58869), .B(n58868), .S0(n43865), .Y(n14747) );
  INVX1 U63268 ( .A(n58870), .Y(n58871) );
  NAND2X1 U63269 ( .A(n58871), .B(n43865), .Y(n58880) );
  NOR2X1 U63270 ( .A(n58880), .B(n44066), .Y(n58872) );
  NOR2X1 U63271 ( .A(n43443), .B(n58872), .Y(n58874) );
  NAND2X1 U63272 ( .A(n44061), .B(n58880), .Y(n58873) );
  MX2X1 U63273 ( .A(n58874), .B(n58873), .S0(n43968), .Y(n14733) );
  INVX1 U63274 ( .A(n58880), .Y(n58875) );
  NAND2X1 U63275 ( .A(n58875), .B(n43968), .Y(n58877) );
  NOR2X1 U63276 ( .A(n44065), .B(n58877), .Y(n58876) );
  NOR2X1 U63277 ( .A(n43443), .B(n58876), .Y(n58879) );
  NAND2X1 U63278 ( .A(n44061), .B(n58877), .Y(n58878) );
  MX2X1 U63279 ( .A(n58879), .B(n58878), .S0(n43958), .Y(n14719) );
  NOR2X1 U63280 ( .A(n43953), .B(n58880), .Y(n58881) );
  NAND2X1 U63281 ( .A(n58881), .B(n43967), .Y(n58885) );
  NOR2X1 U63282 ( .A(n58885), .B(n44066), .Y(n58882) );
  NOR2X1 U63283 ( .A(n43444), .B(n58882), .Y(n58884) );
  NAND2X1 U63284 ( .A(n44062), .B(n58885), .Y(n58883) );
  MX2X1 U63285 ( .A(n58884), .B(n58883), .S0(n43876), .Y(n14705) );
  INVX1 U63286 ( .A(n58885), .Y(n58886) );
  NAND2X1 U63287 ( .A(n58886), .B(n43875), .Y(n58890) );
  NOR2X1 U63288 ( .A(n58890), .B(n44066), .Y(n58887) );
  NOR2X1 U63289 ( .A(n43444), .B(n58887), .Y(n58889) );
  NAND2X1 U63290 ( .A(n44062), .B(n58890), .Y(n58888) );
  MX2X1 U63291 ( .A(n58889), .B(n58888), .S0(n43885), .Y(n14691) );
  INVX1 U63292 ( .A(n58890), .Y(n58891) );
  NAND2X1 U63293 ( .A(n58891), .B(n43885), .Y(n58895) );
  NOR2X1 U63294 ( .A(n58895), .B(n44067), .Y(n58892) );
  NOR2X1 U63295 ( .A(n43444), .B(n58892), .Y(n58894) );
  NAND2X1 U63296 ( .A(n44062), .B(n58895), .Y(n58893) );
  MX2X1 U63297 ( .A(n58894), .B(n58893), .S0(n43895), .Y(n14677) );
  INVX1 U63298 ( .A(n58895), .Y(n58896) );
  NAND2X1 U63299 ( .A(n58896), .B(n43895), .Y(n58911) );
  INVX1 U63300 ( .A(n58911), .Y(n58907) );
  NAND2X1 U63301 ( .A(n44062), .B(n58907), .Y(n58904) );
  INVX1 U63302 ( .A(n58904), .Y(n58897) );
  NOR2X1 U63303 ( .A(n43444), .B(n58897), .Y(n58899) );
  NAND2X1 U63304 ( .A(n44062), .B(n58911), .Y(n58898) );
  MX2X1 U63305 ( .A(n58899), .B(n58898), .S0(n43902), .Y(n14663) );
  NOR2X1 U63306 ( .A(n43898), .B(n58904), .Y(n58900) );
  NOR2X1 U63307 ( .A(n43444), .B(n58900), .Y(n58903) );
  NAND2X1 U63308 ( .A(n58907), .B(n43901), .Y(n58901) );
  NAND2X1 U63309 ( .A(n44062), .B(n58901), .Y(n58902) );
  MX2X1 U63310 ( .A(n58903), .B(n58902), .S0(n43908), .Y(n14649) );
  NOR2X1 U63311 ( .A(n58905), .B(n58904), .Y(n58906) );
  NOR2X1 U63312 ( .A(n43444), .B(n58906), .Y(n58910) );
  NAND2X1 U63313 ( .A(n58912), .B(n58907), .Y(n58908) );
  NAND2X1 U63314 ( .A(n44062), .B(n58908), .Y(n58909) );
  MX2X1 U63315 ( .A(n58910), .B(n58909), .S0(n43915), .Y(n14635) );
  NOR2X1 U63316 ( .A(n43911), .B(n58911), .Y(n58913) );
  NAND2X1 U63317 ( .A(n58913), .B(n58912), .Y(n58917) );
  NOR2X1 U63318 ( .A(n58917), .B(n44064), .Y(n58914) );
  NOR2X1 U63319 ( .A(n43444), .B(n58914), .Y(n58916) );
  NAND2X1 U63320 ( .A(n44062), .B(n58917), .Y(n58915) );
  MX2X1 U63321 ( .A(n58916), .B(n58915), .S0(n43924), .Y(n14621) );
  INVX1 U63322 ( .A(n58917), .Y(n58918) );
  NAND2X1 U63323 ( .A(n58918), .B(n43924), .Y(n58922) );
  NOR2X1 U63324 ( .A(n58922), .B(n44067), .Y(n58919) );
  NOR2X1 U63325 ( .A(n43444), .B(n58919), .Y(n58921) );
  NAND2X1 U63326 ( .A(n44062), .B(n58922), .Y(n58920) );
  MX2X1 U63327 ( .A(n58921), .B(n58920), .S0(n43932), .Y(n14607) );
  INVX1 U63328 ( .A(n58922), .Y(n58927) );
  NAND2X1 U63329 ( .A(n58927), .B(n43931), .Y(n58924) );
  NOR2X1 U63330 ( .A(n44065), .B(n58924), .Y(n58923) );
  NOR2X1 U63331 ( .A(n43444), .B(n58923), .Y(n58926) );
  NAND2X1 U63332 ( .A(n44062), .B(n58924), .Y(n58925) );
  MX2X1 U63333 ( .A(n58926), .B(n58925), .S0(n43939), .Y(n14593) );
  NAND2X1 U63334 ( .A(n58928), .B(n58927), .Y(n58932) );
  NOR2X1 U63335 ( .A(n58932), .B(n44065), .Y(n58929) );
  NOR2X1 U63336 ( .A(n43444), .B(n58929), .Y(n58931) );
  NAND2X1 U63337 ( .A(n44062), .B(n58932), .Y(n58930) );
  MX2X1 U63338 ( .A(n58931), .B(n58930), .S0(n43949), .Y(n14579) );
  INVX1 U63339 ( .A(n58932), .Y(n58933) );
  NAND2X1 U63340 ( .A(n58933), .B(n43949), .Y(n58942) );
  NOR2X1 U63341 ( .A(n58942), .B(n44065), .Y(n58934) );
  NOR2X1 U63342 ( .A(n43444), .B(n58934), .Y(n58936) );
  NAND2X1 U63343 ( .A(n44062), .B(n58942), .Y(n58935) );
  MX2X1 U63344 ( .A(n58936), .B(n58935), .S0(n43978), .Y(n14565) );
  INVX1 U63345 ( .A(n58942), .Y(n58937) );
  NAND2X1 U63346 ( .A(n58937), .B(n43979), .Y(n58939) );
  NOR2X1 U63347 ( .A(n44066), .B(n58939), .Y(n58938) );
  NOR2X1 U63348 ( .A(n43444), .B(n58938), .Y(n58941) );
  NAND2X1 U63349 ( .A(n44063), .B(n58939), .Y(n58940) );
  MX2X1 U63350 ( .A(n58941), .B(n58940), .S0(n43989), .Y(n14551) );
  NOR2X1 U63351 ( .A(n43982), .B(n58942), .Y(n58943) );
  NAND2X1 U63352 ( .A(n58943), .B(n43978), .Y(n58947) );
  NOR2X1 U63353 ( .A(n58947), .B(n44066), .Y(n58944) );
  NOR2X1 U63354 ( .A(n58970), .B(n58944), .Y(n58946) );
  NAND2X1 U63355 ( .A(n44063), .B(n58947), .Y(n58945) );
  MX2X1 U63356 ( .A(n58946), .B(n58945), .S0(n43996), .Y(n14537) );
  INVX1 U63357 ( .A(n58947), .Y(n58948) );
  NAND2X1 U63358 ( .A(n58948), .B(n43996), .Y(n58957) );
  NOR2X1 U63359 ( .A(n58957), .B(n44064), .Y(n58949) );
  NOR2X1 U63360 ( .A(n58970), .B(n58949), .Y(n58951) );
  NAND2X1 U63361 ( .A(n44063), .B(n58957), .Y(n58950) );
  MX2X1 U63362 ( .A(n58951), .B(n58950), .S0(n44006), .Y(n14523) );
  INVX1 U63363 ( .A(n58957), .Y(n58952) );
  NAND2X1 U63364 ( .A(n58952), .B(n44006), .Y(n58954) );
  NOR2X1 U63365 ( .A(n44065), .B(n58954), .Y(n58953) );
  NOR2X1 U63366 ( .A(n43443), .B(n58953), .Y(n58956) );
  NAND2X1 U63367 ( .A(n44063), .B(n58954), .Y(n58955) );
  MX2X1 U63368 ( .A(n58956), .B(n58955), .S0(n44013), .Y(n14509) );
  NOR2X1 U63369 ( .A(n58957), .B(n44010), .Y(n58958) );
  NAND2X1 U63370 ( .A(n58958), .B(n44006), .Y(n58962) );
  NOR2X1 U63371 ( .A(n58962), .B(n44064), .Y(n58959) );
  NOR2X1 U63372 ( .A(n58970), .B(n58959), .Y(n58961) );
  NAND2X1 U63373 ( .A(n44063), .B(n58962), .Y(n58960) );
  MX2X1 U63374 ( .A(n58961), .B(n58960), .S0(n44021), .Y(n14495) );
  INVX1 U63375 ( .A(n58962), .Y(n58963) );
  NAND2X1 U63376 ( .A(n58963), .B(n44021), .Y(n58967) );
  NOR2X1 U63377 ( .A(n58967), .B(n44065), .Y(n58964) );
  NOR2X1 U63378 ( .A(n58970), .B(n58964), .Y(n58966) );
  NAND2X1 U63379 ( .A(n44063), .B(n58967), .Y(n58965) );
  MX2X1 U63380 ( .A(n58966), .B(n58965), .S0(n44029), .Y(n14481) );
  INVX1 U63381 ( .A(n58967), .Y(n58968) );
  NAND2X1 U63382 ( .A(n58968), .B(n44028), .Y(n73376) );
  NOR2X1 U63383 ( .A(n73376), .B(n44064), .Y(n58969) );
  NOR2X1 U63384 ( .A(n58970), .B(n58969), .Y(n58972) );
  NAND2X1 U63385 ( .A(n44063), .B(n73376), .Y(n58971) );
  MX2X1 U63386 ( .A(n58972), .B(n58971), .S0(n44053), .Y(n14462) );
  INVX1 U63387 ( .A(n59112), .Y(n59116) );
  NAND2X1 U63388 ( .A(n43447), .B(n43731), .Y(n58975) );
  INVX1 U63389 ( .A(n58975), .Y(n58981) );
  NOR2X1 U63390 ( .A(n43734), .B(n58977), .Y(n58973) );
  NOR2X1 U63391 ( .A(n58981), .B(n58973), .Y(n14443) );
  NAND2X1 U63392 ( .A(n43447), .B(n43734), .Y(n58974) );
  NAND2X1 U63393 ( .A(n58974), .B(n58977), .Y(n58978) );
  INVX1 U63394 ( .A(n58978), .Y(n58976) );
  MX2X1 U63395 ( .A(n58976), .B(n58975), .S0(n43756), .Y(n14436) );
  NAND2X1 U63396 ( .A(n58977), .B(n43753), .Y(n58979) );
  NAND2X1 U63397 ( .A(n58979), .B(n58978), .Y(n58983) );
  NOR2X1 U63398 ( .A(n43756), .B(n42980), .Y(n58980) );
  NOR2X1 U63399 ( .A(n58981), .B(n58980), .Y(n58982) );
  MX2X1 U63400 ( .A(n58983), .B(n58982), .S0(n43817), .Y(n14426) );
  NOR2X1 U63401 ( .A(n58988), .B(n42981), .Y(n58984) );
  NOR2X1 U63402 ( .A(n43445), .B(n58984), .Y(n58986) );
  NAND2X1 U63403 ( .A(n43447), .B(n58988), .Y(n58985) );
  MX2X1 U63404 ( .A(n58986), .B(n58985), .S0(n43808), .Y(n14419) );
  NAND2X1 U63405 ( .A(n43447), .B(n43807), .Y(n58987) );
  NOR2X1 U63406 ( .A(n58988), .B(n58987), .Y(n58989) );
  NOR2X1 U63407 ( .A(n43445), .B(n58989), .Y(n58993) );
  NAND2X1 U63408 ( .A(n58990), .B(n43807), .Y(n58991) );
  NAND2X1 U63409 ( .A(n43447), .B(n58991), .Y(n58992) );
  NOR2X1 U63410 ( .A(n58998), .B(n42980), .Y(n58994) );
  NOR2X1 U63411 ( .A(n43445), .B(n58994), .Y(n58996) );
  NAND2X1 U63412 ( .A(n43447), .B(n58998), .Y(n58995) );
  MX2X1 U63413 ( .A(n58996), .B(n58995), .S0(n43747), .Y(n14403) );
  NAND2X1 U63414 ( .A(n43447), .B(n43746), .Y(n58997) );
  NOR2X1 U63415 ( .A(n58998), .B(n58997), .Y(n58999) );
  NOR2X1 U63416 ( .A(n43445), .B(n58999), .Y(n59003) );
  NAND2X1 U63417 ( .A(n59000), .B(n43747), .Y(n59001) );
  NAND2X1 U63418 ( .A(n43447), .B(n59001), .Y(n59002) );
  MX2X1 U63419 ( .A(n59003), .B(n59002), .S0(n43793), .Y(n14394) );
  NOR2X1 U63420 ( .A(n59008), .B(n42981), .Y(n59004) );
  NOR2X1 U63421 ( .A(n43445), .B(n59004), .Y(n59006) );
  NAND2X1 U63422 ( .A(n43447), .B(n59008), .Y(n59005) );
  NAND2X1 U63423 ( .A(n43447), .B(n43785), .Y(n59007) );
  NOR2X1 U63424 ( .A(n59008), .B(n59007), .Y(n59009) );
  NOR2X1 U63425 ( .A(n43445), .B(n59009), .Y(n59013) );
  NAND2X1 U63426 ( .A(n59010), .B(n43783), .Y(n59011) );
  NAND2X1 U63427 ( .A(n43447), .B(n59011), .Y(n59012) );
  MX2X1 U63428 ( .A(n59013), .B(n59012), .S0(n43740), .Y(n14378) );
  NOR2X1 U63429 ( .A(n59018), .B(n59112), .Y(n59014) );
  NOR2X1 U63430 ( .A(n43445), .B(n59014), .Y(n59016) );
  NAND2X1 U63431 ( .A(n43447), .B(n59018), .Y(n59015) );
  MX2X1 U63432 ( .A(n59016), .B(n59015), .S0(n43760), .Y(n14371) );
  NAND2X1 U63433 ( .A(n43448), .B(n43760), .Y(n59017) );
  NOR2X1 U63434 ( .A(n59018), .B(n59017), .Y(n59019) );
  NOR2X1 U63435 ( .A(n43445), .B(n59019), .Y(n59023) );
  NAND2X1 U63436 ( .A(n59020), .B(n43760), .Y(n59021) );
  NAND2X1 U63437 ( .A(n43448), .B(n59021), .Y(n59022) );
  MX2X1 U63438 ( .A(n59023), .B(n59022), .S0(n43822), .Y(n14362) );
  NOR2X1 U63439 ( .A(n59028), .B(n42980), .Y(n59024) );
  NOR2X1 U63440 ( .A(n43445), .B(n59024), .Y(n59026) );
  NAND2X1 U63441 ( .A(n43448), .B(n59028), .Y(n59025) );
  NAND2X1 U63442 ( .A(n43448), .B(n43813), .Y(n59027) );
  NOR2X1 U63443 ( .A(n59028), .B(n59027), .Y(n59029) );
  NOR2X1 U63444 ( .A(n43445), .B(n59029), .Y(n59033) );
  NAND2X1 U63445 ( .A(n59030), .B(n43813), .Y(n59031) );
  NAND2X1 U63446 ( .A(n43448), .B(n59031), .Y(n59032) );
  MX2X1 U63447 ( .A(n59033), .B(n59032), .S0(n40460), .Y(n14346) );
  NOR2X1 U63448 ( .A(n59038), .B(n42981), .Y(n59034) );
  NOR2X1 U63449 ( .A(n43445), .B(n59034), .Y(n59036) );
  NAND2X1 U63450 ( .A(n43448), .B(n59038), .Y(n59035) );
  MX2X1 U63451 ( .A(n59036), .B(n59035), .S0(n40477), .Y(n14339) );
  NAND2X1 U63452 ( .A(n43448), .B(n40477), .Y(n59037) );
  NOR2X1 U63453 ( .A(n59038), .B(n59037), .Y(n59039) );
  NOR2X1 U63454 ( .A(n43446), .B(n59039), .Y(n59043) );
  NAND2X1 U63455 ( .A(n59040), .B(n40477), .Y(n59041) );
  NAND2X1 U63456 ( .A(n43448), .B(n59041), .Y(n59042) );
  MX2X1 U63457 ( .A(n59043), .B(n59042), .S0(n43722), .Y(n14330) );
  NOR2X1 U63458 ( .A(n59048), .B(n59112), .Y(n59044) );
  NOR2X1 U63459 ( .A(n43446), .B(n59044), .Y(n59046) );
  NAND2X1 U63460 ( .A(n43448), .B(n59048), .Y(n59045) );
  NAND2X1 U63461 ( .A(n43448), .B(n43789), .Y(n59047) );
  NOR2X1 U63462 ( .A(n59048), .B(n59047), .Y(n59049) );
  NOR2X1 U63463 ( .A(n43446), .B(n59049), .Y(n59053) );
  NAND2X1 U63464 ( .A(n59050), .B(n43789), .Y(n59051) );
  NAND2X1 U63465 ( .A(n43448), .B(n59051), .Y(n59052) );
  MX2X1 U63466 ( .A(n59053), .B(n59052), .S0(n43728), .Y(n14314) );
  NOR2X1 U63467 ( .A(n59058), .B(n42980), .Y(n59054) );
  NOR2X1 U63468 ( .A(n43446), .B(n59054), .Y(n59056) );
  NAND2X1 U63469 ( .A(n43448), .B(n59058), .Y(n59055) );
  MX2X1 U63470 ( .A(n59056), .B(n59055), .S0(n42634), .Y(n14307) );
  NAND2X1 U63471 ( .A(n43449), .B(n42635), .Y(n59057) );
  NOR2X1 U63472 ( .A(n59058), .B(n59057), .Y(n59059) );
  NOR2X1 U63473 ( .A(n43446), .B(n59059), .Y(n59063) );
  NAND2X1 U63474 ( .A(n59060), .B(n42642), .Y(n59061) );
  NAND2X1 U63475 ( .A(n43449), .B(n59061), .Y(n59062) );
  MX2X1 U63476 ( .A(n59063), .B(n59062), .S0(n40538), .Y(n14298) );
  NOR2X1 U63477 ( .A(n59068), .B(n42981), .Y(n59064) );
  NOR2X1 U63478 ( .A(n43446), .B(n59064), .Y(n59066) );
  NAND2X1 U63479 ( .A(n43449), .B(n59068), .Y(n59065) );
  NAND2X1 U63480 ( .A(n43449), .B(n42701), .Y(n59067) );
  NOR2X1 U63481 ( .A(n59068), .B(n59067), .Y(n59069) );
  NOR2X1 U63482 ( .A(n43446), .B(n59069), .Y(n59073) );
  NAND2X1 U63483 ( .A(n59070), .B(n42701), .Y(n59071) );
  NAND2X1 U63484 ( .A(n43449), .B(n59071), .Y(n59072) );
  NOR2X1 U63485 ( .A(n59075), .B(n59112), .Y(n59074) );
  NOR2X1 U63486 ( .A(n43446), .B(n59074), .Y(n59077) );
  NAND2X1 U63487 ( .A(n43449), .B(n59075), .Y(n59076) );
  NOR2X1 U63488 ( .A(n59081), .B(n42980), .Y(n59078) );
  NOR2X1 U63489 ( .A(n43446), .B(n59078), .Y(n59080) );
  NAND2X1 U63490 ( .A(n43449), .B(n59081), .Y(n59079) );
  MX2X1 U63491 ( .A(n59080), .B(n59079), .S0(n43797), .Y(n14266) );
  INVX1 U63492 ( .A(n59081), .Y(n59082) );
  NAND2X1 U63493 ( .A(n43797), .B(n59082), .Y(n59084) );
  NOR2X1 U63494 ( .A(n42981), .B(n59084), .Y(n59083) );
  NOR2X1 U63495 ( .A(n43446), .B(n59083), .Y(n59086) );
  NAND2X1 U63496 ( .A(n43449), .B(n59084), .Y(n59085) );
  NOR2X1 U63497 ( .A(n59088), .B(n42981), .Y(n59087) );
  NOR2X1 U63498 ( .A(n43446), .B(n59087), .Y(n59090) );
  NAND2X1 U63499 ( .A(n43449), .B(n59088), .Y(n59089) );
  MX2X1 U63500 ( .A(n59090), .B(n59089), .S0(n43480), .Y(n14250) );
  NOR2X1 U63501 ( .A(n59094), .B(n59112), .Y(n59091) );
  NOR2X1 U63502 ( .A(n43446), .B(n59091), .Y(n59093) );
  NAND2X1 U63503 ( .A(n43449), .B(n59094), .Y(n59092) );
  INVX1 U63504 ( .A(n59094), .Y(n59095) );
  NAND2X1 U63505 ( .A(n43485), .B(n59095), .Y(n59097) );
  NOR2X1 U63506 ( .A(n59112), .B(n59097), .Y(n59096) );
  NOR2X1 U63507 ( .A(n59114), .B(n59096), .Y(n59099) );
  NAND2X1 U63508 ( .A(n43449), .B(n59097), .Y(n59098) );
  MX2X1 U63509 ( .A(n59099), .B(n59098), .S0(n43489), .Y(n14234) );
  NOR2X1 U63510 ( .A(n59101), .B(n42980), .Y(n59100) );
  NOR2X1 U63511 ( .A(n59114), .B(n59100), .Y(n59103) );
  NAND2X1 U63512 ( .A(n43449), .B(n59101), .Y(n59102) );
  MX2X1 U63513 ( .A(n59103), .B(n59102), .S0(n43495), .Y(n14227) );
  NOR2X1 U63514 ( .A(n59105), .B(n42981), .Y(n59104) );
  NOR2X1 U63515 ( .A(n59114), .B(n59104), .Y(n59107) );
  NAND2X1 U63516 ( .A(n59116), .B(n59105), .Y(n59106) );
  MX2X1 U63517 ( .A(n59107), .B(n59106), .S0(n43498), .Y(n14218) );
  NOR2X1 U63518 ( .A(n59109), .B(n59112), .Y(n59108) );
  NOR2X1 U63519 ( .A(n59114), .B(n59108), .Y(n59111) );
  NAND2X1 U63520 ( .A(n59116), .B(n59109), .Y(n59110) );
  MX2X1 U63521 ( .A(n59111), .B(n59110), .S0(n43504), .Y(n14210) );
  NOR2X1 U63522 ( .A(n42980), .B(n59115), .Y(n59113) );
  NOR2X1 U63523 ( .A(n59114), .B(n59113), .Y(n59118) );
  NAND2X1 U63524 ( .A(n59116), .B(n59115), .Y(n59117) );
  MX2X1 U63525 ( .A(n59118), .B(n59117), .S0(n36706), .Y(n14202) );
  NAND2X1 U63526 ( .A(n43612), .B(n43731), .Y(n72708) );
  NAND2X1 U63527 ( .A(n43926), .B(n43758), .Y(n60566) );
  NAND2X1 U63528 ( .A(n43809), .B(n43905), .Y(n60187) );
  NAND2X1 U63529 ( .A(n40473), .B(n43882), .Y(n59968) );
  NAND2X1 U63530 ( .A(n43952), .B(n40484), .Y(n59764) );
  NAND2X1 U63531 ( .A(n43962), .B(n43788), .Y(n59754) );
  NAND2X1 U63532 ( .A(n43724), .B(n43862), .Y(n59744) );
  NAND2X1 U63533 ( .A(n43850), .B(n42631), .Y(n59669) );
  NAND2X1 U63534 ( .A(n40260), .B(n44038), .Y(n59736) );
  NAND2X1 U63535 ( .A(n43799), .B(n38384), .Y(n59728) );
  NAND2X1 U63536 ( .A(n42652), .B(n39941), .Y(n59270) );
  NAND2X1 U63537 ( .A(n59226), .B(n63194), .Y(n59122) );
  NAND2X1 U63538 ( .A(n59124), .B(n40229), .Y(n59121) );
  NAND2X1 U63539 ( .A(n59122), .B(n59121), .Y(n59123) );
  NAND2X1 U63540 ( .A(n59231), .B(n59123), .Y(n59135) );
  NAND2X1 U63541 ( .A(n42838), .B(n42350), .Y(n59166) );
  NAND2X1 U63542 ( .A(n42825), .B(n39794), .Y(n59134) );
  XNOR2X1 U63543 ( .A(n59245), .B(n40446), .Y(n59125) );
  INVX1 U63544 ( .A(n59189), .Y(n59165) );
  NAND2X1 U63545 ( .A(n59168), .B(n40228), .Y(n59173) );
  NAND2X1 U63546 ( .A(n59166), .B(n40390), .Y(n59174) );
  INVX1 U63547 ( .A(n59175), .Y(n59129) );
  NAND2X1 U63548 ( .A(n59128), .B(n59134), .Y(n59130) );
  NAND2X1 U63549 ( .A(n59129), .B(n36722), .Y(n59160) );
  NAND2X1 U63550 ( .A(n59160), .B(n59161), .Y(n59131) );
  INVX1 U63551 ( .A(n59131), .Y(n59132) );
  NAND2X1 U63552 ( .A(n59132), .B(n59189), .Y(n59133) );
  INVX1 U63553 ( .A(n59252), .Y(n59254) );
  XNOR2X1 U63554 ( .A(n39761), .B(n40619), .Y(n59140) );
  INVX1 U63555 ( .A(n59140), .Y(n59137) );
  NOR2X1 U63556 ( .A(n59137), .B(n40379), .Y(n59139) );
  INVX1 U63557 ( .A(n59245), .Y(n59136) );
  NAND2X1 U63558 ( .A(n59136), .B(n40278), .Y(n59242) );
  NOR2X1 U63559 ( .A(n59137), .B(n40429), .Y(n59138) );
  NOR2X1 U63560 ( .A(n59139), .B(n59138), .Y(n59143) );
  NOR2X1 U63561 ( .A(n59140), .B(n42812), .Y(n59141) );
  NAND2X1 U63562 ( .A(n59141), .B(n40429), .Y(n59142) );
  NAND2X1 U63563 ( .A(n59143), .B(n59142), .Y(n59154) );
  NAND2X1 U63564 ( .A(n59224), .B(n42347), .Y(n59676) );
  NAND2X1 U63565 ( .A(n38493), .B(n38827), .Y(n61185) );
  NAND2X1 U63566 ( .A(n40371), .B(n42822), .Y(n59678) );
  NAND2X1 U63567 ( .A(n38527), .B(n59147), .Y(n59152) );
  NAND2X1 U63568 ( .A(n59150), .B(n38527), .Y(n59151) );
  NAND2X1 U63569 ( .A(n59152), .B(n59151), .Y(n59153) );
  INVX1 U63570 ( .A(n59231), .Y(n59232) );
  XNOR2X1 U63571 ( .A(n42817), .B(n59154), .Y(n59155) );
  XNOR2X1 U63572 ( .A(n59254), .B(n59155), .Y(n59264) );
  INVX1 U63573 ( .A(n59264), .Y(n59266) );
  NAND2X1 U63574 ( .A(n39022), .B(n41751), .Y(n59156) );
  NOR2X1 U63575 ( .A(n36636), .B(n59156), .Y(n59159) );
  NOR2X1 U63576 ( .A(n59157), .B(n59160), .Y(n59158) );
  NOR2X1 U63577 ( .A(n59159), .B(n59158), .Y(n59164) );
  NOR2X1 U63578 ( .A(n39022), .B(n38485), .Y(n59162) );
  NAND2X1 U63579 ( .A(n59162), .B(n59161), .Y(n59163) );
  NAND2X1 U63580 ( .A(n59164), .B(n59163), .Y(n59192) );
  NAND2X1 U63581 ( .A(n59167), .B(n59168), .Y(n59171) );
  INVX1 U63582 ( .A(n59168), .Y(n59169) );
  NOR2X1 U63583 ( .A(n43459), .B(n59169), .Y(n59170) );
  XNOR2X1 U63584 ( .A(n59171), .B(n59170), .Y(n59172) );
  XNOR2X1 U63585 ( .A(n36722), .B(n59172), .Y(n59181) );
  INVX1 U63586 ( .A(n59181), .Y(n59208) );
  NAND2X1 U63587 ( .A(n59201), .B(n63824), .Y(n59198) );
  INVX1 U63588 ( .A(n59200), .Y(n59196) );
  NAND2X1 U63589 ( .A(n59174), .B(n59173), .Y(n59176) );
  NAND2X1 U63590 ( .A(n59176), .B(n59175), .Y(n59177) );
  NAND2X1 U63591 ( .A(n72783), .B(n43457), .Y(n59194) );
  INVX1 U63592 ( .A(n59194), .Y(n59179) );
  NAND2X1 U63593 ( .A(n59177), .B(n59200), .Y(n59178) );
  NAND2X1 U63594 ( .A(n59208), .B(n59180), .Y(n59182) );
  NAND2X1 U63595 ( .A(n42648), .B(n40392), .Y(n59209) );
  NAND2X1 U63596 ( .A(n59182), .B(n59183), .Y(n59193) );
  NAND2X1 U63597 ( .A(n42815), .B(n59193), .Y(n59188) );
  NAND2X1 U63598 ( .A(n42651), .B(n43466), .Y(n59190) );
  INVX1 U63599 ( .A(n59190), .Y(n59186) );
  NAND2X1 U63600 ( .A(n59183), .B(n59182), .Y(n59184) );
  OR2X1 U63601 ( .A(n42815), .B(n59184), .Y(n59185) );
  NAND2X1 U63602 ( .A(n59186), .B(n59185), .Y(n59187) );
  NAND2X1 U63603 ( .A(n59188), .B(n59187), .Y(n59265) );
  XNOR2X1 U63604 ( .A(n59190), .B(n59189), .Y(n59191) );
  XNOR2X1 U63605 ( .A(n59194), .B(n38859), .Y(n59195) );
  XNOR2X1 U63606 ( .A(n59196), .B(n59195), .Y(n59307) );
  INVX1 U63607 ( .A(n59307), .Y(n59204) );
  NAND2X1 U63608 ( .A(n39698), .B(n43458), .Y(n59299) );
  INVX1 U63609 ( .A(n59299), .Y(n59282) );
  NAND2X1 U63610 ( .A(n59199), .B(n59198), .Y(n59197) );
  NAND2X1 U63611 ( .A(n59282), .B(n59197), .Y(n59203) );
  NAND2X1 U63612 ( .A(n39698), .B(n38813), .Y(n59284) );
  NAND2X1 U63613 ( .A(n59201), .B(n44071), .Y(n59285) );
  INVX1 U63614 ( .A(n59294), .Y(n59202) );
  NAND2X1 U63615 ( .A(n40596), .B(n59202), .Y(n59297) );
  NAND2X1 U63616 ( .A(n59203), .B(n59297), .Y(n59205) );
  NAND2X1 U63617 ( .A(n43800), .B(n40393), .Y(n59298) );
  INVX1 U63618 ( .A(n59298), .Y(n59207) );
  XNOR2X1 U63619 ( .A(n59209), .B(n59208), .Y(n59210) );
  XNOR2X1 U63620 ( .A(n59210), .B(n39051), .Y(n59212) );
  NAND2X1 U63621 ( .A(n43800), .B(n43465), .Y(n59280) );
  INVX1 U63622 ( .A(n59280), .Y(n59214) );
  INVX1 U63623 ( .A(n59212), .Y(n59279) );
  NAND2X1 U63624 ( .A(n42840), .B(n59279), .Y(n59213) );
  NAND2X1 U63625 ( .A(n43800), .B(n39942), .Y(n59313) );
  INVX1 U63626 ( .A(n59313), .Y(n59217) );
  INVX1 U63627 ( .A(n59215), .Y(n59312) );
  NAND2X1 U63628 ( .A(n40628), .B(n59312), .Y(n59216) );
  NAND2X1 U63629 ( .A(n43800), .B(n43843), .Y(n59278) );
  INVX1 U63630 ( .A(n59278), .Y(n59327) );
  NAND2X1 U63631 ( .A(n39754), .B(n59330), .Y(n59218) );
  NOR2X1 U63632 ( .A(n42828), .B(n59244), .Y(n59220) );
  NOR2X1 U63633 ( .A(n42817), .B(n42828), .Y(n59219) );
  NOR2X1 U63634 ( .A(n59220), .B(n59219), .Y(n59223) );
  NAND2X1 U63635 ( .A(n40619), .B(n59221), .Y(n59222) );
  NAND2X1 U63636 ( .A(n42221), .B(n40253), .Y(n59890) );
  NAND2X1 U63637 ( .A(n40391), .B(n59890), .Y(n59883) );
  NAND2X1 U63638 ( .A(n36715), .B(n42347), .Y(n60243) );
  NAND2X1 U63639 ( .A(n60243), .B(n63824), .Y(n59882) );
  NAND2X1 U63640 ( .A(n59883), .B(n59882), .Y(n59225) );
  NAND2X1 U63641 ( .A(n59225), .B(n42816), .Y(n59679) );
  NAND2X1 U63642 ( .A(n59226), .B(n43458), .Y(n59230) );
  NOR2X1 U63643 ( .A(n59228), .B(n59227), .Y(n59229) );
  NOR2X1 U63644 ( .A(n59684), .B(n39909), .Y(n59234) );
  NAND2X1 U63645 ( .A(n59686), .B(n59689), .Y(n59233) );
  NOR2X1 U63646 ( .A(n59234), .B(n59233), .Y(n59239) );
  OR2X1 U63647 ( .A(n59689), .B(n59686), .Y(n59237) );
  NOR2X1 U63648 ( .A(n59684), .B(n59689), .Y(n59235) );
  NAND2X1 U63649 ( .A(n59235), .B(n59685), .Y(n59236) );
  NAND2X1 U63650 ( .A(n59237), .B(n59236), .Y(n59238) );
  NOR2X1 U63651 ( .A(n59239), .B(n59238), .Y(n59240) );
  XOR2X1 U63652 ( .A(n59691), .B(n59240), .Y(n59696) );
  XNOR2X1 U63653 ( .A(n59696), .B(n41779), .Y(n59241) );
  XNOR2X1 U63654 ( .A(n40662), .B(n59241), .Y(n59705) );
  NAND2X1 U63655 ( .A(n40379), .B(n59244), .Y(n59243) );
  NOR2X1 U63656 ( .A(n38994), .B(n59243), .Y(n59250) );
  NAND2X1 U63657 ( .A(n40619), .B(n42812), .Y(n59248) );
  NOR2X1 U63658 ( .A(n59245), .B(n59244), .Y(n59246) );
  NAND2X1 U63659 ( .A(n59246), .B(n40278), .Y(n59247) );
  NAND2X1 U63660 ( .A(n59248), .B(n59247), .Y(n59249) );
  NOR2X1 U63661 ( .A(n59250), .B(n59249), .Y(n59251) );
  XNOR2X1 U63662 ( .A(n42817), .B(n59251), .Y(n59253) );
  NAND2X1 U63663 ( .A(n59253), .B(n59252), .Y(n59701) );
  NAND2X1 U63664 ( .A(n39942), .B(n42709), .Y(n59702) );
  NAND2X1 U63665 ( .A(n59701), .B(n59702), .Y(n59256) );
  NAND2X1 U63666 ( .A(n39761), .B(n59258), .Y(n59700) );
  INVX1 U63667 ( .A(n59700), .Y(n59255) );
  NOR2X1 U63668 ( .A(n59256), .B(n59255), .Y(n59263) );
  OR2X1 U63669 ( .A(n59702), .B(n59701), .Y(n59261) );
  NOR2X1 U63670 ( .A(n59257), .B(n59702), .Y(n59259) );
  NAND2X1 U63671 ( .A(n59259), .B(n59258), .Y(n59260) );
  NAND2X1 U63672 ( .A(n59261), .B(n59260), .Y(n59262) );
  NAND2X1 U63673 ( .A(n59265), .B(n59264), .Y(n59712) );
  NAND2X1 U63674 ( .A(n42653), .B(n43843), .Y(n59717) );
  NAND2X1 U63675 ( .A(n59712), .B(n59717), .Y(n59269) );
  INVX1 U63676 ( .A(n59270), .Y(n59267) );
  NAND2X1 U63677 ( .A(n59267), .B(n59271), .Y(n59711) );
  INVX1 U63678 ( .A(n59711), .Y(n59268) );
  NOR2X1 U63679 ( .A(n59269), .B(n59268), .Y(n59276) );
  OR2X1 U63680 ( .A(n59717), .B(n59712), .Y(n59274) );
  NOR2X1 U63681 ( .A(n59270), .B(n59717), .Y(n59272) );
  NAND2X1 U63682 ( .A(n59272), .B(n59271), .Y(n59273) );
  NAND2X1 U63683 ( .A(n59274), .B(n59273), .Y(n59275) );
  XNOR2X1 U63684 ( .A(n59736), .B(n38765), .Y(n59325) );
  NAND2X1 U63685 ( .A(n40260), .B(n38381), .Y(n59321) );
  NOR2X1 U63686 ( .A(n59318), .B(n59321), .Y(n59320) );
  XNOR2X1 U63687 ( .A(n59280), .B(n59279), .Y(n59281) );
  XNOR2X1 U63688 ( .A(n59281), .B(n42840), .Y(n59378) );
  INVX1 U63689 ( .A(n59378), .Y(n59308) );
  XNOR2X1 U63690 ( .A(n59294), .B(n59282), .Y(n59283) );
  XNOR2X1 U63691 ( .A(n40596), .B(n59283), .Y(n59363) );
  INVX1 U63692 ( .A(n59363), .Y(n59289) );
  NAND2X1 U63693 ( .A(n72815), .B(n44070), .Y(n59341) );
  INVX1 U63694 ( .A(n59342), .Y(n59338) );
  NAND2X1 U63695 ( .A(n59285), .B(n59284), .Y(n59287) );
  NAND2X1 U63696 ( .A(n39699), .B(n38471), .Y(n59286) );
  NAND2X1 U63697 ( .A(n59287), .B(n59286), .Y(n59288) );
  INVX1 U63698 ( .A(n59288), .Y(n59339) );
  NAND2X1 U63699 ( .A(n59338), .B(n59339), .Y(n59353) );
  NAND2X1 U63700 ( .A(n59288), .B(n59342), .Y(n59356) );
  NAND2X1 U63701 ( .A(n43772), .B(n40393), .Y(n59354) );
  INVX1 U63702 ( .A(n59354), .Y(n59292) );
  NAND2X1 U63703 ( .A(n40597), .B(n59363), .Y(n59291) );
  NAND2X1 U63704 ( .A(n59294), .B(n59293), .Y(n59300) );
  NAND2X1 U63705 ( .A(n59297), .B(n59298), .Y(n59295) );
  NOR2X1 U63706 ( .A(n59296), .B(n59295), .Y(n59305) );
  OR2X1 U63707 ( .A(n59298), .B(n59297), .Y(n59303) );
  NOR2X1 U63708 ( .A(n59299), .B(n59298), .Y(n59301) );
  NAND2X1 U63709 ( .A(n59301), .B(n59300), .Y(n59302) );
  NAND2X1 U63710 ( .A(n59303), .B(n59302), .Y(n59304) );
  NOR2X1 U63711 ( .A(n59305), .B(n59304), .Y(n59306) );
  NAND2X1 U63712 ( .A(n59336), .B(n36771), .Y(n59368) );
  NAND2X1 U63713 ( .A(n40260), .B(n43465), .Y(n59370) );
  INVX1 U63714 ( .A(n59370), .Y(n59335) );
  NAND2X1 U63715 ( .A(n40259), .B(n39937), .Y(n59369) );
  INVX1 U63716 ( .A(n59369), .Y(n59311) );
  XNOR2X1 U63717 ( .A(n59313), .B(n59312), .Y(n59314) );
  XNOR2X1 U63718 ( .A(n59314), .B(n40628), .Y(n59315) );
  INVX1 U63719 ( .A(n59315), .Y(n59332) );
  NAND2X1 U63720 ( .A(n40259), .B(n43843), .Y(n59333) );
  INVX1 U63721 ( .A(n59333), .Y(n59317) );
  NAND2X1 U63722 ( .A(n40638), .B(n59315), .Y(n59316) );
  NOR2X1 U63723 ( .A(n42829), .B(n59318), .Y(n59319) );
  NOR2X1 U63724 ( .A(n59320), .B(n59319), .Y(n59324) );
  INVX1 U63725 ( .A(n59321), .Y(n59326) );
  NAND2X1 U63726 ( .A(n59326), .B(n59322), .Y(n59323) );
  NAND2X1 U63727 ( .A(n59324), .B(n59323), .Y(n59735) );
  INVX1 U63728 ( .A(n59735), .Y(n59738) );
  XNOR2X1 U63729 ( .A(n59669), .B(n38294), .Y(n59385) );
  XNOR2X1 U63730 ( .A(n59327), .B(n59326), .Y(n59328) );
  XNOR2X1 U63731 ( .A(n59328), .B(n39754), .Y(n59329) );
  XNOR2X1 U63732 ( .A(n59330), .B(n59329), .Y(n59331) );
  XNOR2X1 U63733 ( .A(n42829), .B(n59331), .Y(n59452) );
  INVX1 U63734 ( .A(n59452), .Y(n59381) );
  XNOR2X1 U63735 ( .A(n59333), .B(n59332), .Y(n59334) );
  XNOR2X1 U63736 ( .A(n59334), .B(n40638), .Y(n59443) );
  XNOR2X1 U63737 ( .A(n59336), .B(n59335), .Y(n59337) );
  XNOR2X1 U63738 ( .A(n36771), .B(n59337), .Y(n59436) );
  INVX1 U63739 ( .A(n59419), .Y(n59346) );
  INVX1 U63740 ( .A(n59396), .Y(n59392) );
  NAND2X1 U63741 ( .A(n59341), .B(n59340), .Y(n59343) );
  NAND2X1 U63742 ( .A(n59343), .B(n59342), .Y(n59344) );
  NAND2X1 U63743 ( .A(n59392), .B(n39898), .Y(n59410) );
  NAND2X1 U63744 ( .A(n43456), .B(n36499), .Y(n59412) );
  INVX1 U63745 ( .A(n59412), .Y(n59345) );
  NAND2X1 U63746 ( .A(n59344), .B(n59396), .Y(n59413) );
  NAND2X1 U63747 ( .A(n59345), .B(n59413), .Y(n59407) );
  NAND2X1 U63748 ( .A(n43472), .B(n42636), .Y(n59411) );
  INVX1 U63749 ( .A(n59411), .Y(n59349) );
  NAND2X1 U63750 ( .A(n59353), .B(n59354), .Y(n59352) );
  INVX1 U63751 ( .A(n59350), .Y(n59351) );
  NOR2X1 U63752 ( .A(n59352), .B(n59351), .Y(n59361) );
  OR2X1 U63753 ( .A(n59354), .B(n59353), .Y(n59359) );
  NOR2X1 U63754 ( .A(n59355), .B(n59354), .Y(n59357) );
  NAND2X1 U63755 ( .A(n59357), .B(n59356), .Y(n59358) );
  NAND2X1 U63756 ( .A(n59359), .B(n59358), .Y(n59360) );
  NOR2X1 U63757 ( .A(n59361), .B(n59360), .Y(n59362) );
  NAND2X1 U63758 ( .A(n59390), .B(n37378), .Y(n59426) );
  NAND2X1 U63759 ( .A(n43465), .B(n42638), .Y(n59428) );
  INVX1 U63760 ( .A(n59428), .Y(n59389) );
  NAND2X1 U63761 ( .A(n59389), .B(n59429), .Y(n59423) );
  NAND2X1 U63762 ( .A(n59426), .B(n59423), .Y(n59364) );
  NAND2X1 U63763 ( .A(n39940), .B(n42639), .Y(n59427) );
  INVX1 U63764 ( .A(n59427), .Y(n59366) );
  NAND2X1 U63765 ( .A(n59368), .B(n59369), .Y(n59367) );
  NOR2X1 U63766 ( .A(n59367), .B(n39046), .Y(n59376) );
  OR2X1 U63767 ( .A(n59369), .B(n59368), .Y(n59374) );
  NOR2X1 U63768 ( .A(n59370), .B(n59369), .Y(n59372) );
  NAND2X1 U63769 ( .A(n59372), .B(n59371), .Y(n59373) );
  NAND2X1 U63770 ( .A(n59374), .B(n59373), .Y(n59375) );
  NOR2X1 U63771 ( .A(n59376), .B(n59375), .Y(n59377) );
  XOR2X1 U63772 ( .A(n59378), .B(n59377), .Y(n59379) );
  INVX1 U63773 ( .A(n59379), .Y(n59388) );
  NAND2X1 U63774 ( .A(n59379), .B(n40583), .Y(n59380) );
  NAND2X1 U63775 ( .A(n59443), .B(n39090), .Y(n59382) );
  NAND2X1 U63776 ( .A(n38379), .B(n42641), .Y(n59444) );
  NAND2X1 U63777 ( .A(n59382), .B(n59383), .Y(n59451) );
  XNOR2X1 U63778 ( .A(n59386), .B(n41483), .Y(n59387) );
  XNOR2X1 U63779 ( .A(n59388), .B(n59387), .Y(n59510) );
  XNOR2X1 U63780 ( .A(n59390), .B(n59389), .Y(n59391) );
  XNOR2X1 U63781 ( .A(n37378), .B(n59391), .Y(n59421) );
  XNOR2X1 U63782 ( .A(n59412), .B(n59392), .Y(n59393) );
  XNOR2X1 U63783 ( .A(n39898), .B(n59393), .Y(n59403) );
  INVX1 U63784 ( .A(n59403), .Y(n59485) );
  NAND2X1 U63785 ( .A(n38110), .B(n42718), .Y(n59473) );
  INVX1 U63786 ( .A(n59475), .Y(n59470) );
  NAND2X1 U63787 ( .A(n59397), .B(n59396), .Y(n59398) );
  NAND2X1 U63788 ( .A(n59470), .B(n39421), .Y(n59402) );
  NAND2X1 U63789 ( .A(n38111), .B(n43458), .Y(n59471) );
  INVX1 U63790 ( .A(n59471), .Y(n59400) );
  NAND2X1 U63791 ( .A(n59398), .B(n59475), .Y(n59399) );
  NAND2X1 U63792 ( .A(n59400), .B(n59399), .Y(n59401) );
  NAND2X1 U63793 ( .A(n59402), .B(n59401), .Y(n59483) );
  NAND2X1 U63794 ( .A(n59485), .B(n59483), .Y(n59406) );
  NAND2X1 U63795 ( .A(n40343), .B(n59403), .Y(n59404) );
  NAND2X1 U63796 ( .A(n42150), .B(n59404), .Y(n59405) );
  NAND2X1 U63797 ( .A(n59410), .B(n59411), .Y(n59409) );
  INVX1 U63798 ( .A(n59407), .Y(n59408) );
  NOR2X1 U63799 ( .A(n59409), .B(n59408), .Y(n59418) );
  OR2X1 U63800 ( .A(n59411), .B(n59410), .Y(n59416) );
  NOR2X1 U63801 ( .A(n59412), .B(n59411), .Y(n59414) );
  NAND2X1 U63802 ( .A(n59414), .B(n59413), .Y(n59415) );
  NAND2X1 U63803 ( .A(n59416), .B(n59415), .Y(n59417) );
  INVX1 U63804 ( .A(n59420), .Y(n59469) );
  INVX1 U63805 ( .A(n59421), .Y(n59494) );
  NAND2X1 U63806 ( .A(n38529), .B(n59494), .Y(n59422) );
  NAND2X1 U63807 ( .A(n59426), .B(n59427), .Y(n59425) );
  INVX1 U63808 ( .A(n59423), .Y(n59424) );
  NOR2X1 U63809 ( .A(n59425), .B(n59424), .Y(n59434) );
  OR2X1 U63810 ( .A(n59427), .B(n59426), .Y(n59432) );
  NOR2X1 U63811 ( .A(n59428), .B(n59427), .Y(n59430) );
  NAND2X1 U63812 ( .A(n59430), .B(n59429), .Y(n59431) );
  NAND2X1 U63813 ( .A(n59432), .B(n59431), .Y(n59433) );
  NOR2X1 U63814 ( .A(n59434), .B(n59433), .Y(n59435) );
  XOR2X1 U63815 ( .A(n59436), .B(n59435), .Y(n59437) );
  NAND2X1 U63816 ( .A(n43725), .B(n43842), .Y(n59502) );
  INVX1 U63817 ( .A(n59502), .Y(n59463) );
  INVX1 U63818 ( .A(n59437), .Y(n59466) );
  NAND2X1 U63819 ( .A(n59463), .B(n59503), .Y(n59499) );
  NAND2X1 U63820 ( .A(n38803), .B(n59499), .Y(n59438) );
  NAND2X1 U63821 ( .A(n59510), .B(n59438), .Y(n59442) );
  NAND2X1 U63822 ( .A(n43724), .B(n38381), .Y(n59501) );
  INVX1 U63823 ( .A(n59501), .Y(n59440) );
  NAND2X1 U63824 ( .A(n59440), .B(n59439), .Y(n59441) );
  NAND2X1 U63825 ( .A(n59442), .B(n59441), .Y(n59447) );
  XNOR2X1 U63826 ( .A(n59445), .B(n59444), .Y(n59446) );
  INVX1 U63827 ( .A(n59448), .Y(n59460) );
  NAND2X1 U63828 ( .A(n43724), .B(n44038), .Y(n59461) );
  INVX1 U63829 ( .A(n59461), .Y(n59450) );
  INVX1 U63830 ( .A(n59447), .Y(n59462) );
  NAND2X1 U63831 ( .A(n59462), .B(n59448), .Y(n59449) );
  XNOR2X1 U63832 ( .A(n59452), .B(n41495), .Y(n59453) );
  NAND2X1 U63833 ( .A(n59454), .B(n59455), .Y(n59459) );
  NAND2X1 U63834 ( .A(n43724), .B(n43853), .Y(n59521) );
  INVX1 U63835 ( .A(n59521), .Y(n59457) );
  INVX1 U63836 ( .A(n59455), .Y(n59520) );
  NAND2X1 U63837 ( .A(n59457), .B(n59456), .Y(n59458) );
  NAND2X1 U63838 ( .A(n59459), .B(n59458), .Y(n59743) );
  INVX1 U63839 ( .A(n59749), .Y(n59750) );
  XNOR2X1 U63840 ( .A(n59754), .B(n59750), .Y(n59527) );
  XNOR2X1 U63841 ( .A(n59464), .B(n59463), .Y(n59465) );
  XNOR2X1 U63842 ( .A(n59467), .B(n42155), .Y(n59468) );
  XNOR2X1 U63843 ( .A(n59469), .B(n59468), .Y(n59491) );
  XNOR2X1 U63844 ( .A(n59471), .B(n59470), .Y(n59472) );
  XNOR2X1 U63845 ( .A(n39421), .B(n59472), .Y(n59480) );
  INVX1 U63846 ( .A(n59480), .Y(n59555) );
  NAND2X1 U63847 ( .A(n42718), .B(n72807), .Y(n59543) );
  NAND2X1 U63848 ( .A(n38110), .B(n73384), .Y(n59544) );
  INVX1 U63849 ( .A(n59545), .Y(n59540) );
  NAND2X1 U63850 ( .A(n59474), .B(n59473), .Y(n59476) );
  NAND2X1 U63851 ( .A(n59476), .B(n59475), .Y(n59477) );
  NAND2X1 U63852 ( .A(n43456), .B(n43786), .Y(n59541) );
  INVX1 U63853 ( .A(n59541), .Y(n59479) );
  NAND2X1 U63854 ( .A(n59477), .B(n59545), .Y(n59478) );
  INVX1 U63855 ( .A(n59553), .Y(n59481) );
  NAND2X1 U63856 ( .A(n59481), .B(n59480), .Y(n59482) );
  XNOR2X1 U63857 ( .A(n59483), .B(n42150), .Y(n59484) );
  NAND2X1 U63858 ( .A(n59538), .B(n59486), .Y(n59490) );
  INVX1 U63859 ( .A(n59538), .Y(n59487) );
  NAND2X1 U63860 ( .A(n59487), .B(n38216), .Y(n59488) );
  NAND2X1 U63861 ( .A(n41795), .B(n59488), .Y(n59489) );
  NAND2X1 U63862 ( .A(n59490), .B(n59489), .Y(n59561) );
  INVX1 U63863 ( .A(n59491), .Y(n59563) );
  XNOR2X1 U63864 ( .A(n36524), .B(n42160), .Y(n59493) );
  XNOR2X1 U63865 ( .A(n59494), .B(n59493), .Y(n59495) );
  INVX1 U63866 ( .A(n59495), .Y(n59537) );
  NAND2X1 U63867 ( .A(n43840), .B(n43787), .Y(n59571) );
  INVX1 U63868 ( .A(n59571), .Y(n59534) );
  NAND2X1 U63869 ( .A(n38378), .B(n43788), .Y(n59570) );
  INVX1 U63870 ( .A(n59570), .Y(n59498) );
  NAND2X1 U63871 ( .A(n38803), .B(n59501), .Y(n59500) );
  NOR2X1 U63872 ( .A(n59500), .B(n39780), .Y(n59508) );
  OR2X1 U63873 ( .A(n59501), .B(n38803), .Y(n59506) );
  NOR2X1 U63874 ( .A(n59502), .B(n59501), .Y(n59504) );
  NAND2X1 U63875 ( .A(n59504), .B(n59503), .Y(n59505) );
  NAND2X1 U63876 ( .A(n59506), .B(n59505), .Y(n59507) );
  NOR2X1 U63877 ( .A(n59508), .B(n59507), .Y(n59509) );
  XOR2X1 U63878 ( .A(n59510), .B(n59509), .Y(n59512) );
  NAND2X1 U63879 ( .A(n44035), .B(n43788), .Y(n59532) );
  INVX1 U63880 ( .A(n59532), .Y(n59514) );
  INVX1 U63881 ( .A(n59512), .Y(n59531) );
  NAND2X1 U63882 ( .A(n40580), .B(n59531), .Y(n59513) );
  NAND2X1 U63883 ( .A(n59515), .B(n36602), .Y(n59519) );
  NAND2X1 U63884 ( .A(n43850), .B(n43788), .Y(n59585) );
  INVX1 U63885 ( .A(n59585), .Y(n59517) );
  NAND2X1 U63886 ( .A(n40622), .B(n38705), .Y(n59516) );
  NAND2X1 U63887 ( .A(n59517), .B(n59516), .Y(n59518) );
  NAND2X1 U63888 ( .A(n59519), .B(n59518), .Y(n59530) );
  INVX1 U63889 ( .A(n59530), .Y(n59522) );
  NOR2X1 U63890 ( .A(n59522), .B(n59528), .Y(n59524) );
  NAND2X1 U63891 ( .A(n43859), .B(n43788), .Y(n59529) );
  NOR2X1 U63892 ( .A(n59522), .B(n59529), .Y(n59523) );
  NOR2X1 U63893 ( .A(n59524), .B(n59523), .Y(n59526) );
  OR2X1 U63894 ( .A(n59528), .B(n59529), .Y(n59525) );
  NAND2X1 U63895 ( .A(n59526), .B(n59525), .Y(n59748) );
  INVX1 U63896 ( .A(n59748), .Y(n59751) );
  XNOR2X1 U63897 ( .A(n59527), .B(n59751), .Y(n59765) );
  INVX1 U63898 ( .A(n59765), .Y(n59762) );
  XNOR2X1 U63899 ( .A(n59532), .B(n59531), .Y(n59533) );
  XNOR2X1 U63900 ( .A(n59535), .B(n59534), .Y(n59536) );
  XNOR2X1 U63901 ( .A(n59538), .B(n41795), .Y(n59539) );
  XNOR2X1 U63902 ( .A(n38216), .B(n59539), .Y(n59558) );
  INVX1 U63903 ( .A(n59558), .Y(n59628) );
  XNOR2X1 U63904 ( .A(n59541), .B(n59540), .Y(n59542) );
  XNOR2X1 U63905 ( .A(n39795), .B(n59542), .Y(n59551) );
  INVX1 U63906 ( .A(n59551), .Y(n59618) );
  NAND2X1 U63907 ( .A(n42716), .B(n72741), .Y(n59606) );
  NAND2X1 U63908 ( .A(n40390), .B(n72807), .Y(n59607) );
  NAND2X1 U63909 ( .A(n59544), .B(n59543), .Y(n59546) );
  NAND2X1 U63910 ( .A(n59546), .B(n59545), .Y(n59604) );
  INVX1 U63911 ( .A(n59604), .Y(n59547) );
  NAND2X1 U63912 ( .A(n39361), .B(n59547), .Y(n59550) );
  NAND2X1 U63913 ( .A(n59608), .B(n59604), .Y(n59548) );
  NAND2X1 U63914 ( .A(n41760), .B(n59548), .Y(n59549) );
  NAND2X1 U63915 ( .A(n59550), .B(n59549), .Y(n59616) );
  NAND2X1 U63916 ( .A(n39774), .B(n59551), .Y(n59552) );
  XNOR2X1 U63917 ( .A(n59553), .B(n41773), .Y(n59554) );
  XNOR2X1 U63918 ( .A(n59555), .B(n59554), .Y(n59556) );
  INVX1 U63919 ( .A(n59556), .Y(n59603) );
  NAND2X1 U63920 ( .A(n40653), .B(n59603), .Y(n59557) );
  INVX1 U63921 ( .A(n59626), .Y(n59559) );
  NAND2X1 U63922 ( .A(n59558), .B(n59559), .Y(n59560) );
  XNOR2X1 U63923 ( .A(n59561), .B(n41808), .Y(n59562) );
  XNOR2X1 U63924 ( .A(n59563), .B(n59562), .Y(n59564) );
  INVX1 U63925 ( .A(n59564), .Y(n59600) );
  NAND2X1 U63926 ( .A(n59564), .B(n40362), .Y(n59565) );
  NAND2X1 U63927 ( .A(n40047), .B(n40578), .Y(n59567) );
  NAND2X1 U63928 ( .A(n59569), .B(n59570), .Y(n59568) );
  NOR2X1 U63929 ( .A(n59568), .B(n38505), .Y(n59577) );
  OR2X1 U63930 ( .A(n59570), .B(n59569), .Y(n59575) );
  NOR2X1 U63931 ( .A(n59571), .B(n59570), .Y(n59573) );
  NAND2X1 U63932 ( .A(n59573), .B(n59572), .Y(n59574) );
  NAND2X1 U63933 ( .A(n59575), .B(n59574), .Y(n59576) );
  NAND2X1 U63934 ( .A(n59597), .B(n40598), .Y(n59580) );
  NAND2X1 U63935 ( .A(n41854), .B(n59578), .Y(n59579) );
  NAND2X1 U63936 ( .A(n59580), .B(n59579), .Y(n59581) );
  NAND2X1 U63937 ( .A(n43850), .B(n40483), .Y(n59645) );
  INVX1 U63938 ( .A(n59645), .Y(n59584) );
  INVX1 U63939 ( .A(n59581), .Y(n59646) );
  NAND2X1 U63940 ( .A(n59646), .B(n59582), .Y(n59583) );
  XNOR2X1 U63941 ( .A(n59585), .B(n38705), .Y(n59586) );
  XNOR2X1 U63942 ( .A(n59586), .B(n40622), .Y(n59587) );
  INVX1 U63943 ( .A(n59587), .Y(n59594) );
  NAND2X1 U63944 ( .A(n43859), .B(n40482), .Y(n59595) );
  INVX1 U63945 ( .A(n59595), .Y(n59589) );
  NAND2X1 U63946 ( .A(n39762), .B(n59587), .Y(n59588) );
  NAND2X1 U63947 ( .A(n59590), .B(n36527), .Y(n59766) );
  NAND2X1 U63948 ( .A(n43962), .B(n40483), .Y(n59591) );
  INVX1 U63949 ( .A(n59590), .Y(n59592) );
  NAND2X1 U63950 ( .A(n59766), .B(n59767), .Y(n59763) );
  XNOR2X1 U63951 ( .A(n59591), .B(n39592), .Y(n59593) );
  XNOR2X1 U63952 ( .A(n59593), .B(n59592), .Y(n59661) );
  INVX1 U63953 ( .A(n59661), .Y(n59844) );
  XNOR2X1 U63954 ( .A(n59595), .B(n59594), .Y(n59596) );
  XNOR2X1 U63955 ( .A(n39762), .B(n59596), .Y(n59655) );
  XNOR2X1 U63956 ( .A(n59597), .B(n41854), .Y(n59598) );
  XNOR2X1 U63957 ( .A(n40598), .B(n59598), .Y(n59642) );
  XNOR2X1 U63958 ( .A(n38796), .B(n41827), .Y(n59599) );
  XNOR2X1 U63959 ( .A(n59600), .B(n59599), .Y(n59632) );
  XNOR2X1 U63960 ( .A(n59601), .B(n41797), .Y(n59602) );
  XNOR2X1 U63961 ( .A(n59603), .B(n59602), .Y(n59623) );
  INVX1 U63962 ( .A(n59623), .Y(n59812) );
  XNOR2X1 U63963 ( .A(n59604), .B(n39361), .Y(n59605) );
  XNOR2X1 U63964 ( .A(n59605), .B(n41760), .Y(n59612) );
  INVX1 U63965 ( .A(n59612), .Y(n59803) );
  NAND2X1 U63966 ( .A(n73384), .B(n72741), .Y(n59792) );
  INVX1 U63967 ( .A(n59793), .Y(n59788) );
  NAND2X1 U63968 ( .A(n59607), .B(n59606), .Y(n59609) );
  NAND2X1 U63969 ( .A(n59609), .B(n59608), .Y(n59789) );
  INVX1 U63970 ( .A(n59789), .Y(n59610) );
  NAND2X1 U63971 ( .A(n59793), .B(n59789), .Y(n59611) );
  NAND2X1 U63972 ( .A(n59803), .B(n39607), .Y(n59615) );
  NAND2X1 U63973 ( .A(n40264), .B(n59612), .Y(n59613) );
  NAND2X1 U63974 ( .A(n41778), .B(n59613), .Y(n59614) );
  NAND2X1 U63975 ( .A(n59615), .B(n59614), .Y(n59785) );
  XNOR2X1 U63976 ( .A(n59616), .B(n41774), .Y(n59617) );
  XNOR2X1 U63977 ( .A(n59618), .B(n59617), .Y(n59619) );
  NAND2X1 U63978 ( .A(n59785), .B(n59619), .Y(n59622) );
  INVX1 U63979 ( .A(n59619), .Y(n59787) );
  NAND2X1 U63980 ( .A(n41794), .B(n59620), .Y(n59621) );
  NAND2X1 U63981 ( .A(n59622), .B(n59621), .Y(n59810) );
  INVX1 U63982 ( .A(n59810), .Y(n59624) );
  NAND2X1 U63983 ( .A(n59624), .B(n59623), .Y(n59625) );
  XNOR2X1 U63984 ( .A(n59626), .B(n41812), .Y(n59627) );
  XNOR2X1 U63985 ( .A(n59628), .B(n59627), .Y(n59629) );
  INVX1 U63986 ( .A(n59782), .Y(n59630) );
  INVX1 U63987 ( .A(n59629), .Y(n59784) );
  NAND2X1 U63988 ( .A(n59630), .B(n59784), .Y(n59631) );
  INVX1 U63989 ( .A(n59819), .Y(n59633) );
  INVX1 U63990 ( .A(n59632), .Y(n59821) );
  NAND2X1 U63991 ( .A(n59633), .B(n59821), .Y(n59634) );
  XNOR2X1 U63992 ( .A(n59635), .B(n41842), .Y(n59636) );
  XNOR2X1 U63993 ( .A(n40578), .B(n59636), .Y(n59637) );
  INVX1 U63994 ( .A(n59637), .Y(n59781) );
  NAND2X1 U63995 ( .A(n36419), .B(n59781), .Y(n59640) );
  NAND2X1 U63996 ( .A(n40666), .B(n59637), .Y(n59638) );
  NAND2X1 U63997 ( .A(n41849), .B(n59638), .Y(n59639) );
  NAND2X1 U63998 ( .A(n59640), .B(n59639), .Y(n59641) );
  NAND2X1 U63999 ( .A(n40470), .B(n43853), .Y(n59831) );
  INVX1 U64000 ( .A(n59831), .Y(n59644) );
  INVX1 U64001 ( .A(n59641), .Y(n59832) );
  INVX1 U64002 ( .A(n59642), .Y(n59830) );
  NAND2X1 U64003 ( .A(n59832), .B(n59830), .Y(n59643) );
  XNOR2X1 U64004 ( .A(n59645), .B(n38232), .Y(n59647) );
  XNOR2X1 U64005 ( .A(n59647), .B(n59646), .Y(n59649) );
  NAND2X1 U64006 ( .A(n59648), .B(n59649), .Y(n59653) );
  NAND2X1 U64007 ( .A(n40470), .B(n43862), .Y(n59777) );
  INVX1 U64008 ( .A(n59777), .Y(n59651) );
  INVX1 U64009 ( .A(n59648), .Y(n59778) );
  INVX1 U64010 ( .A(n59649), .Y(n59776) );
  NAND2X1 U64011 ( .A(n59651), .B(n59650), .Y(n59652) );
  NAND2X1 U64012 ( .A(n59653), .B(n59652), .Y(n59654) );
  NAND2X1 U64013 ( .A(n59655), .B(n59654), .Y(n59659) );
  NAND2X1 U64014 ( .A(n40471), .B(n43965), .Y(n59773) );
  INVX1 U64015 ( .A(n59773), .Y(n59657) );
  INVX1 U64016 ( .A(n59654), .Y(n59774) );
  INVX1 U64017 ( .A(n59655), .Y(n59772) );
  NAND2X1 U64018 ( .A(n59657), .B(n59656), .Y(n59658) );
  NAND2X1 U64019 ( .A(n59659), .B(n59658), .Y(n59660) );
  NAND2X1 U64020 ( .A(n40472), .B(n43955), .Y(n59845) );
  INVX1 U64021 ( .A(n59845), .Y(n59663) );
  INVX1 U64022 ( .A(n59660), .Y(n59846) );
  NAND2X1 U64023 ( .A(n59846), .B(n59661), .Y(n59662) );
  INVX1 U64024 ( .A(n59664), .Y(n59852) );
  INVX1 U64025 ( .A(n59665), .Y(n59854) );
  XNOR2X1 U64026 ( .A(n59968), .B(n39313), .Y(n59771) );
  NAND2X1 U64027 ( .A(n43869), .B(n40485), .Y(n59962) );
  NAND2X1 U64028 ( .A(n43724), .B(n43964), .Y(n59951) );
  NAND2X1 U64029 ( .A(n43859), .B(n42643), .Y(n59941) );
  NAND2X1 U64030 ( .A(n59668), .B(n59667), .Y(n59673) );
  INVX1 U64031 ( .A(n59669), .Y(n59671) );
  NAND2X1 U64032 ( .A(n36437), .B(n38294), .Y(n59670) );
  NAND2X1 U64033 ( .A(n59671), .B(n59670), .Y(n59672) );
  NAND2X1 U64034 ( .A(n59673), .B(n59672), .Y(n59936) );
  XNOR2X1 U64035 ( .A(n59941), .B(n36723), .Y(n59742) );
  NAND2X1 U64036 ( .A(n40259), .B(n43853), .Y(n59931) );
  NAND2X1 U64037 ( .A(n43840), .B(n42709), .Y(n59900) );
  NAND2X1 U64038 ( .A(n39938), .B(n43795), .Y(n59864) );
  NAND2X1 U64039 ( .A(n43465), .B(n43776), .Y(n59868) );
  NAND2X1 U64040 ( .A(n43471), .B(n43479), .Y(n59874) );
  NAND2X1 U64041 ( .A(n38614), .B(n40574), .Y(n60240) );
  NAND2X1 U64042 ( .A(n40391), .B(n71033), .Y(n59675) );
  NAND2X1 U64043 ( .A(n40524), .B(n40394), .Y(n59674) );
  NAND2X1 U64044 ( .A(n40121), .B(n60227), .Y(n59881) );
  NAND2X1 U64045 ( .A(n60243), .B(n38527), .Y(n59879) );
  INVX1 U64046 ( .A(n59875), .Y(n59873) );
  XNOR2X1 U64047 ( .A(n59874), .B(n59873), .Y(n59683) );
  OR2X1 U64048 ( .A(n59679), .B(n59678), .Y(n59682) );
  NOR2X1 U64049 ( .A(n43481), .B(n43460), .Y(n59680) );
  NAND2X1 U64050 ( .A(n59682), .B(n59681), .Y(n59872) );
  XNOR2X1 U64051 ( .A(n59683), .B(n38444), .Y(n59867) );
  INVX1 U64052 ( .A(n59867), .Y(n59869) );
  INVX1 U64053 ( .A(n59691), .Y(n59688) );
  NAND2X1 U64054 ( .A(n40626), .B(n59685), .Y(n59687) );
  NAND2X1 U64055 ( .A(n59687), .B(n59686), .Y(n59690) );
  INVX1 U64056 ( .A(n59689), .Y(n59693) );
  NAND2X1 U64057 ( .A(n38107), .B(n59691), .Y(n59692) );
  XNOR2X1 U64058 ( .A(n59864), .B(n38280), .Y(n59699) );
  INVX1 U64059 ( .A(n59696), .Y(n59695) );
  NAND2X1 U64060 ( .A(n59695), .B(n59694), .Y(n59698) );
  NAND2X1 U64061 ( .A(n59698), .B(n59697), .Y(n59863) );
  INVX1 U64062 ( .A(n59863), .Y(n59866) );
  XNOR2X1 U64063 ( .A(n59699), .B(n59866), .Y(n59898) );
  INVX1 U64064 ( .A(n59898), .Y(n59901) );
  XNOR2X1 U64065 ( .A(n59900), .B(n59901), .Y(n59710) );
  NAND2X1 U64066 ( .A(n59701), .B(n59700), .Y(n59704) );
  NOR2X1 U64067 ( .A(n59705), .B(n59704), .Y(n59703) );
  NOR2X1 U64068 ( .A(n59703), .B(n59702), .Y(n59709) );
  INVX1 U64069 ( .A(n59704), .Y(n59707) );
  INVX1 U64070 ( .A(n59705), .Y(n59706) );
  NOR2X1 U64071 ( .A(n59707), .B(n59706), .Y(n59708) );
  OR2X1 U64072 ( .A(n59709), .B(n59708), .Y(n59899) );
  INVX1 U64073 ( .A(n59899), .Y(n59902) );
  XNOR2X1 U64074 ( .A(n59710), .B(n59902), .Y(n60213) );
  NAND2X1 U64075 ( .A(n59712), .B(n59711), .Y(n59713) );
  NAND2X1 U64076 ( .A(n59713), .B(n59714), .Y(n59909) );
  NAND2X1 U64077 ( .A(n42654), .B(n38383), .Y(n59913) );
  NAND2X1 U64078 ( .A(n59909), .B(n59913), .Y(n59716) );
  INVX1 U64079 ( .A(n59717), .Y(n59715) );
  NAND2X1 U64080 ( .A(n59715), .B(n59718), .Y(n59908) );
  NOR2X1 U64081 ( .A(n59716), .B(n36618), .Y(n59723) );
  OR2X1 U64082 ( .A(n59913), .B(n59909), .Y(n59721) );
  NOR2X1 U64083 ( .A(n59717), .B(n59913), .Y(n59719) );
  NAND2X1 U64084 ( .A(n59719), .B(n59718), .Y(n59720) );
  NAND2X1 U64085 ( .A(n59721), .B(n59720), .Y(n59722) );
  NAND2X1 U64086 ( .A(n59725), .B(n59724), .Y(n59922) );
  NAND2X1 U64087 ( .A(n43798), .B(n44037), .Y(n59924) );
  INVX1 U64088 ( .A(n59728), .Y(n59726) );
  NAND2X1 U64089 ( .A(n59726), .B(n59729), .Y(n59921) );
  NOR2X1 U64090 ( .A(n59727), .B(n39824), .Y(n59734) );
  OR2X1 U64091 ( .A(n59924), .B(n59922), .Y(n59732) );
  NOR2X1 U64092 ( .A(n59728), .B(n59924), .Y(n59730) );
  NAND2X1 U64093 ( .A(n59730), .B(n59729), .Y(n59731) );
  NAND2X1 U64094 ( .A(n59732), .B(n59731), .Y(n59733) );
  INVX1 U64095 ( .A(n59932), .Y(n59930) );
  XNOR2X1 U64096 ( .A(n59931), .B(n59930), .Y(n59741) );
  INVX1 U64097 ( .A(n59736), .Y(n59740) );
  NAND2X1 U64098 ( .A(n59738), .B(n59737), .Y(n59739) );
  XNOR2X1 U64099 ( .A(n59741), .B(n40656), .Y(n59937) );
  INVX1 U64100 ( .A(n59937), .Y(n59938) );
  XNOR2X1 U64101 ( .A(n59742), .B(n59938), .Y(n59952) );
  INVX1 U64102 ( .A(n59952), .Y(n59950) );
  XNOR2X1 U64103 ( .A(n59951), .B(n59950), .Y(n59747) );
  INVX1 U64104 ( .A(n59744), .Y(n59746) );
  XNOR2X1 U64105 ( .A(n59747), .B(n40586), .Y(n59956) );
  NAND2X1 U64106 ( .A(n59749), .B(n59748), .Y(n59954) );
  NAND2X1 U64107 ( .A(n43952), .B(n43788), .Y(n59957) );
  NAND2X1 U64108 ( .A(n59954), .B(n59957), .Y(n59753) );
  INVX1 U64109 ( .A(n59754), .Y(n59752) );
  NAND2X1 U64110 ( .A(n59752), .B(n59755), .Y(n59953) );
  NOR2X1 U64111 ( .A(n59753), .B(n39745), .Y(n59760) );
  OR2X1 U64112 ( .A(n59957), .B(n59954), .Y(n59758) );
  NOR2X1 U64113 ( .A(n59754), .B(n59957), .Y(n59756) );
  NAND2X1 U64114 ( .A(n59756), .B(n59755), .Y(n59757) );
  NAND2X1 U64115 ( .A(n59758), .B(n59757), .Y(n59759) );
  NOR2X1 U64116 ( .A(n59760), .B(n59759), .Y(n59761) );
  XOR2X1 U64117 ( .A(n59956), .B(n59761), .Y(n59961) );
  INVX1 U64118 ( .A(n59961), .Y(n59963) );
  XNOR2X1 U64119 ( .A(n59962), .B(n59963), .Y(n59770) );
  NAND2X1 U64120 ( .A(n59763), .B(n59762), .Y(n59769) );
  NAND2X1 U64121 ( .A(n59769), .B(n59768), .Y(n59960) );
  XNOR2X1 U64122 ( .A(n59770), .B(n36685), .Y(n59969) );
  INVX1 U64123 ( .A(n59969), .Y(n59967) );
  XNOR2X1 U64124 ( .A(n59771), .B(n59967), .Y(n59860) );
  XNOR2X1 U64125 ( .A(n59773), .B(n59772), .Y(n59775) );
  XNOR2X1 U64126 ( .A(n59775), .B(n59774), .Y(n59841) );
  INVX1 U64127 ( .A(n59841), .Y(n59977) );
  XNOR2X1 U64128 ( .A(n59777), .B(n59776), .Y(n59779) );
  XNOR2X1 U64129 ( .A(n59779), .B(n59778), .Y(n59837) );
  INVX1 U64130 ( .A(n59837), .Y(n60044) );
  XNOR2X1 U64131 ( .A(n36419), .B(n41849), .Y(n59780) );
  XNOR2X1 U64132 ( .A(n59781), .B(n59780), .Y(n59827) );
  XNOR2X1 U64133 ( .A(n59782), .B(n41828), .Y(n59783) );
  XNOR2X1 U64134 ( .A(n59784), .B(n59783), .Y(n59817) );
  INVX1 U64135 ( .A(n59817), .Y(n60019) );
  XNOR2X1 U64136 ( .A(n59785), .B(n41794), .Y(n59786) );
  XNOR2X1 U64137 ( .A(n59789), .B(n59788), .Y(n59790) );
  XNOR2X1 U64138 ( .A(n59790), .B(n41759), .Y(n59799) );
  INVX1 U64139 ( .A(n59799), .Y(n60004) );
  INVX1 U64140 ( .A(n59996), .Y(n59991) );
  NAND2X1 U64141 ( .A(n59792), .B(n59791), .Y(n59794) );
  NAND2X1 U64142 ( .A(n59794), .B(n59793), .Y(n59992) );
  INVX1 U64143 ( .A(n59992), .Y(n59795) );
  NAND2X1 U64144 ( .A(n59991), .B(n59795), .Y(n59798) );
  NAND2X1 U64145 ( .A(n59996), .B(n59992), .Y(n59796) );
  NAND2X1 U64146 ( .A(n41761), .B(n59796), .Y(n59797) );
  NAND2X1 U64147 ( .A(n60004), .B(n60005), .Y(n59802) );
  NAND2X1 U64148 ( .A(n40625), .B(n59799), .Y(n59800) );
  NAND2X1 U64149 ( .A(n41780), .B(n59800), .Y(n59801) );
  NAND2X1 U64150 ( .A(n59802), .B(n59801), .Y(n59989) );
  XNOR2X1 U64151 ( .A(n39607), .B(n59803), .Y(n59804) );
  XNOR2X1 U64152 ( .A(n59804), .B(n41778), .Y(n59805) );
  NAND2X1 U64153 ( .A(n59989), .B(n59805), .Y(n59808) );
  INVX1 U64154 ( .A(n59805), .Y(n59988) );
  NAND2X1 U64155 ( .A(n41798), .B(n59806), .Y(n59807) );
  NAND2X1 U64156 ( .A(n59808), .B(n59807), .Y(n60011) );
  XNOR2X1 U64157 ( .A(n59810), .B(n41809), .Y(n59811) );
  XNOR2X1 U64158 ( .A(n59812), .B(n59811), .Y(n59813) );
  NAND2X1 U64159 ( .A(n59985), .B(n59813), .Y(n59816) );
  INVX1 U64160 ( .A(n59813), .Y(n59987) );
  NAND2X1 U64161 ( .A(n40659), .B(n59987), .Y(n59814) );
  NAND2X1 U64162 ( .A(n41830), .B(n59814), .Y(n59815) );
  NAND2X1 U64163 ( .A(n59816), .B(n59815), .Y(n60017) );
  NAND2X1 U64164 ( .A(n39392), .B(n59817), .Y(n59818) );
  XNOR2X1 U64165 ( .A(n59819), .B(n41839), .Y(n59820) );
  XNOR2X1 U64166 ( .A(n59821), .B(n59820), .Y(n59822) );
  INVX1 U64167 ( .A(n59822), .Y(n59984) );
  NAND2X1 U64168 ( .A(n59982), .B(n59984), .Y(n59826) );
  INVX1 U64169 ( .A(n59982), .Y(n59823) );
  NAND2X1 U64170 ( .A(n59823), .B(n59822), .Y(n59824) );
  NAND2X1 U64171 ( .A(n41858), .B(n59824), .Y(n59825) );
  NAND2X1 U64172 ( .A(n59826), .B(n59825), .Y(n60031) );
  INVX1 U64173 ( .A(n60031), .Y(n59828) );
  INVX1 U64174 ( .A(n59827), .Y(n60033) );
  NAND2X1 U64175 ( .A(n59828), .B(n60033), .Y(n59829) );
  XNOR2X1 U64176 ( .A(n59831), .B(n59830), .Y(n59833) );
  XNOR2X1 U64177 ( .A(n59833), .B(n59832), .Y(n59834) );
  INVX1 U64178 ( .A(n59834), .Y(n59979) );
  NAND2X1 U64179 ( .A(n43859), .B(n40468), .Y(n59980) );
  INVX1 U64180 ( .A(n59980), .Y(n59836) );
  NAND2X1 U64181 ( .A(n40649), .B(n59834), .Y(n59835) );
  NAND2X1 U64182 ( .A(n43962), .B(n40468), .Y(n60043) );
  INVX1 U64183 ( .A(n60043), .Y(n59839) );
  NAND2X1 U64184 ( .A(n39230), .B(n59837), .Y(n59838) );
  INVX1 U64185 ( .A(n59840), .Y(n59975) );
  INVX1 U64186 ( .A(n59976), .Y(n59842) );
  NAND2X1 U64187 ( .A(n59842), .B(n59841), .Y(n59843) );
  XNOR2X1 U64188 ( .A(n59845), .B(n59844), .Y(n59847) );
  XNOR2X1 U64189 ( .A(n59847), .B(n59846), .Y(n59849) );
  NAND2X1 U64190 ( .A(n43869), .B(n40461), .Y(n59973) );
  INVX1 U64191 ( .A(n59973), .Y(n59851) );
  INVX1 U64192 ( .A(n59849), .Y(n59972) );
  NAND2X1 U64193 ( .A(n36603), .B(n59972), .Y(n59850) );
  XNOR2X1 U64194 ( .A(n59853), .B(n59852), .Y(n59855) );
  XNOR2X1 U64195 ( .A(n59855), .B(n59854), .Y(n59857) );
  INVX1 U64196 ( .A(n59857), .Y(n60061) );
  NAND2X1 U64197 ( .A(n40462), .B(n43882), .Y(n60062) );
  INVX1 U64198 ( .A(n60062), .Y(n60057) );
  INVX1 U64199 ( .A(n59856), .Y(n60063) );
  NAND2X1 U64200 ( .A(n40461), .B(n43892), .Y(n60066) );
  INVX1 U64201 ( .A(n60066), .Y(n59862) );
  INVX1 U64202 ( .A(n59859), .Y(n60065) );
  INVX1 U64203 ( .A(n59860), .Y(n60067) );
  NAND2X1 U64204 ( .A(n43869), .B(n43788), .Y(n60193) );
  NAND2X1 U64205 ( .A(n43798), .B(n43853), .Y(n60208) );
  NAND2X1 U64206 ( .A(n38380), .B(n42708), .Y(n60663) );
  NAND2X1 U64207 ( .A(n43841), .B(n43795), .Y(n60260) );
  XNOR2X1 U64208 ( .A(n60260), .B(n40111), .Y(n59897) );
  INVX1 U64209 ( .A(n59868), .Y(n59871) );
  NAND2X1 U64210 ( .A(n40601), .B(n59869), .Y(n59870) );
  NAND2X1 U64211 ( .A(n39938), .B(n43776), .Y(n60252) );
  NAND2X1 U64212 ( .A(n43464), .B(n43479), .Y(n60254) );
  INVX1 U64213 ( .A(n60254), .Y(n60225) );
  XNOR2X1 U64214 ( .A(n60252), .B(n60225), .Y(n59878) );
  INVX1 U64215 ( .A(n59874), .Y(n59877) );
  NAND2X1 U64216 ( .A(n38444), .B(n59875), .Y(n59876) );
  XNOR2X1 U64217 ( .A(n59878), .B(n39194), .Y(n59895) );
  NAND2X1 U64218 ( .A(n70371), .B(n43472), .Y(n59884) );
  INVX1 U64219 ( .A(n59879), .Y(n59880) );
  XNOR2X1 U64220 ( .A(n59884), .B(n39617), .Y(n59894) );
  NAND2X1 U64221 ( .A(n41749), .B(n40577), .Y(n60607) );
  INVX1 U64222 ( .A(n60607), .Y(n60606) );
  NOR2X1 U64223 ( .A(n41749), .B(n40577), .Y(n59885) );
  NOR2X1 U64224 ( .A(n60606), .B(n59885), .Y(n59893) );
  INVX1 U64225 ( .A(n60240), .Y(n60942) );
  NAND2X1 U64226 ( .A(n36736), .B(n59886), .Y(n59888) );
  NOR2X1 U64227 ( .A(n36725), .B(n59888), .Y(n59889) );
  NAND2X1 U64228 ( .A(n70671), .B(n62659), .Y(n60228) );
  XNOR2X1 U64229 ( .A(n59893), .B(n59892), .Y(n60247) );
  INVX1 U64230 ( .A(n60247), .Y(n60246) );
  XNOR2X1 U64231 ( .A(n59894), .B(n60246), .Y(n60223) );
  INVX1 U64232 ( .A(n60223), .Y(n60253) );
  XNOR2X1 U64233 ( .A(n59895), .B(n60253), .Y(n59896) );
  XNOR2X1 U64234 ( .A(n60663), .B(n37377), .Y(n59907) );
  NAND2X1 U64235 ( .A(n59899), .B(n59898), .Y(n59906) );
  INVX1 U64236 ( .A(n59900), .Y(n59904) );
  NAND2X1 U64237 ( .A(n59902), .B(n59901), .Y(n59903) );
  NAND2X1 U64238 ( .A(n59904), .B(n59903), .Y(n59905) );
  NAND2X1 U64239 ( .A(n59906), .B(n59905), .Y(n60263) );
  INVX1 U64240 ( .A(n60263), .Y(n60262) );
  XNOR2X1 U64241 ( .A(n59907), .B(n60262), .Y(n60221) );
  INVX1 U64242 ( .A(n60221), .Y(n60218) );
  NAND2X1 U64243 ( .A(n42654), .B(n44037), .Y(n60216) );
  INVX1 U64244 ( .A(n60216), .Y(n60222) );
  INVX1 U64245 ( .A(n59913), .Y(n60215) );
  NAND2X1 U64246 ( .A(n60222), .B(n60215), .Y(n59915) );
  NAND2X1 U64247 ( .A(n59909), .B(n59908), .Y(n60212) );
  NOR2X1 U64248 ( .A(n59910), .B(n60213), .Y(n59919) );
  NOR2X1 U64249 ( .A(n60222), .B(n36734), .Y(n59912) );
  NAND2X1 U64250 ( .A(n60215), .B(n60212), .Y(n59911) );
  NAND2X1 U64251 ( .A(n60216), .B(n59913), .Y(n59914) );
  NAND2X1 U64252 ( .A(n40399), .B(n59914), .Y(n59917) );
  NAND2X1 U64253 ( .A(n59915), .B(n60212), .Y(n59916) );
  NOR2X1 U64254 ( .A(n59919), .B(n59918), .Y(n59920) );
  XNOR2X1 U64255 ( .A(n60218), .B(n59920), .Y(n60207) );
  INVX1 U64256 ( .A(n60207), .Y(n60209) );
  XNOR2X1 U64257 ( .A(n60208), .B(n60209), .Y(n59929) );
  NAND2X1 U64258 ( .A(n59922), .B(n59921), .Y(n59925) );
  INVX1 U64259 ( .A(n59926), .Y(n59923) );
  INVX1 U64260 ( .A(n59924), .Y(n59928) );
  NAND2X1 U64261 ( .A(n40375), .B(n59926), .Y(n59927) );
  XNOR2X1 U64262 ( .A(n59929), .B(n40663), .Y(n60205) );
  INVX1 U64263 ( .A(n59931), .Y(n59934) );
  NAND2X1 U64264 ( .A(n40656), .B(n59932), .Y(n59933) );
  XNOR2X1 U64265 ( .A(n37390), .B(n42181), .Y(n59935) );
  XNOR2X1 U64266 ( .A(n38728), .B(n59935), .Y(n60198) );
  NAND2X1 U64267 ( .A(n59937), .B(n59936), .Y(n60197) );
  NAND2X1 U64268 ( .A(n43962), .B(n42644), .Y(n60199) );
  NAND2X1 U64269 ( .A(n60199), .B(n60197), .Y(n59940) );
  INVX1 U64270 ( .A(n59941), .Y(n59939) );
  NAND2X1 U64271 ( .A(n36723), .B(n59938), .Y(n59942) );
  NOR2X1 U64272 ( .A(n59940), .B(n37371), .Y(n59947) );
  OR2X1 U64273 ( .A(n60199), .B(n60197), .Y(n59945) );
  NOR2X1 U64274 ( .A(n59941), .B(n60199), .Y(n59943) );
  NAND2X1 U64275 ( .A(n59943), .B(n59942), .Y(n59944) );
  NAND2X1 U64276 ( .A(n59945), .B(n59944), .Y(n59946) );
  NOR2X1 U64277 ( .A(n59947), .B(n59946), .Y(n59948) );
  XOR2X1 U64278 ( .A(n60198), .B(n59948), .Y(n60276) );
  NAND2X1 U64279 ( .A(n43724), .B(n43955), .Y(n60272) );
  NAND2X1 U64280 ( .A(n59950), .B(n59949), .Y(n60273) );
  NAND2X1 U64281 ( .A(n60273), .B(n60274), .Y(n60271) );
  NAND2X1 U64282 ( .A(n59954), .B(n59953), .Y(n59955) );
  NAND2X1 U64283 ( .A(n36489), .B(n59956), .Y(n60194) );
  NOR2X1 U64284 ( .A(n59956), .B(n59955), .Y(n59958) );
  OR2X1 U64285 ( .A(n59958), .B(n59957), .Y(n60195) );
  NAND2X1 U64286 ( .A(n60194), .B(n60195), .Y(n60192) );
  INVX1 U64287 ( .A(n59959), .Y(n60288) );
  XNOR2X1 U64288 ( .A(n60284), .B(n60288), .Y(n59966) );
  INVX1 U64289 ( .A(n59962), .Y(n59965) );
  INVX1 U64290 ( .A(n60283), .Y(n60286) );
  XNOR2X1 U64291 ( .A(n59966), .B(n60286), .Y(n60292) );
  NAND2X1 U64292 ( .A(n40474), .B(n43892), .Y(n60291) );
  NAND2X1 U64293 ( .A(n59967), .B(n36567), .Y(n60293) );
  NAND2X1 U64294 ( .A(n60293), .B(n60294), .Y(n60289) );
  XOR2X1 U64295 ( .A(n60291), .B(n60289), .Y(n59970) );
  XOR2X1 U64296 ( .A(n60292), .B(n59970), .Y(n60298) );
  INVX1 U64297 ( .A(n60298), .Y(n60300) );
  XNOR2X1 U64298 ( .A(n60299), .B(n60300), .Y(n59971) );
  XNOR2X1 U64299 ( .A(n59971), .B(n41944), .Y(n60188) );
  INVX1 U64300 ( .A(n60188), .Y(n60186) );
  XNOR2X1 U64301 ( .A(n60187), .B(n60186), .Y(n60075) );
  NAND2X1 U64302 ( .A(n43809), .B(n43891), .Y(n60080) );
  INVX1 U64303 ( .A(n60080), .Y(n60060) );
  XNOR2X1 U64304 ( .A(n59973), .B(n59972), .Y(n59974) );
  XNOR2X1 U64305 ( .A(n59974), .B(n36603), .Y(n60170) );
  INVX1 U64306 ( .A(n60170), .Y(n60053) );
  XNOR2X1 U64307 ( .A(n59976), .B(n59975), .Y(n59978) );
  XNOR2X1 U64308 ( .A(n59978), .B(n59977), .Y(n60052) );
  XNOR2X1 U64309 ( .A(n59980), .B(n59979), .Y(n59981) );
  XNOR2X1 U64310 ( .A(n40649), .B(n59981), .Y(n60089) );
  XNOR2X1 U64311 ( .A(n59982), .B(n41858), .Y(n59983) );
  XNOR2X1 U64312 ( .A(n59984), .B(n59983), .Y(n60026) );
  XNOR2X1 U64313 ( .A(n59985), .B(n41830), .Y(n59986) );
  XNOR2X1 U64314 ( .A(n59987), .B(n59986), .Y(n60015) );
  INVX1 U64315 ( .A(n60015), .Y(n60143) );
  XNOR2X1 U64316 ( .A(n59989), .B(n59988), .Y(n59990) );
  XNOR2X1 U64317 ( .A(n59990), .B(n41798), .Y(n60009) );
  INVX1 U64318 ( .A(n60009), .Y(n60133) );
  XNOR2X1 U64319 ( .A(n59992), .B(n59991), .Y(n59993) );
  XNOR2X1 U64320 ( .A(n59993), .B(n41761), .Y(n60002) );
  INVX1 U64321 ( .A(n60002), .Y(n60123) );
  NAND2X1 U64322 ( .A(n42715), .B(n43811), .Y(n60110) );
  INVX1 U64323 ( .A(n60112), .Y(n60107) );
  NAND2X1 U64324 ( .A(n59995), .B(n59994), .Y(n59997) );
  NAND2X1 U64325 ( .A(n59997), .B(n59996), .Y(n60108) );
  INVX1 U64326 ( .A(n60108), .Y(n59998) );
  NAND2X1 U64327 ( .A(n60107), .B(n59998), .Y(n60001) );
  NAND2X1 U64328 ( .A(n60112), .B(n60108), .Y(n59999) );
  NAND2X1 U64329 ( .A(n41769), .B(n59999), .Y(n60000) );
  NAND2X1 U64330 ( .A(n60001), .B(n60000), .Y(n60124) );
  NAND2X1 U64331 ( .A(n39632), .B(n60002), .Y(n60003) );
  XNOR2X1 U64332 ( .A(n60005), .B(n60004), .Y(n60006) );
  XNOR2X1 U64333 ( .A(n60006), .B(n41780), .Y(n60007) );
  INVX1 U64334 ( .A(n60007), .Y(n60105) );
  NAND2X1 U64335 ( .A(n39560), .B(n60009), .Y(n60010) );
  XNOR2X1 U64336 ( .A(n60011), .B(n41815), .Y(n60012) );
  XNOR2X1 U64337 ( .A(n36786), .B(n60012), .Y(n60013) );
  INVX1 U64338 ( .A(n60013), .Y(n60104) );
  NAND2X1 U64339 ( .A(n40635), .B(n60104), .Y(n60014) );
  NAND2X1 U64340 ( .A(n40053), .B(n60015), .Y(n60016) );
  XNOR2X1 U64341 ( .A(n60017), .B(n41843), .Y(n60018) );
  NAND2X1 U64342 ( .A(n37982), .B(n60020), .Y(n60024) );
  NAND2X1 U64343 ( .A(n44036), .B(n72820), .Y(n60100) );
  INVX1 U64344 ( .A(n60100), .Y(n60022) );
  NAND2X1 U64345 ( .A(n39458), .B(n38247), .Y(n60021) );
  NAND2X1 U64346 ( .A(n60022), .B(n60021), .Y(n60023) );
  NAND2X1 U64347 ( .A(n60024), .B(n60023), .Y(n60025) );
  NAND2X1 U64348 ( .A(n60026), .B(n60025), .Y(n60030) );
  NAND2X1 U64349 ( .A(n43850), .B(n43810), .Y(n60097) );
  INVX1 U64350 ( .A(n60097), .Y(n60028) );
  INVX1 U64351 ( .A(n60025), .Y(n60098) );
  INVX1 U64352 ( .A(n60026), .Y(n60096) );
  NAND2X1 U64353 ( .A(n60098), .B(n60096), .Y(n60027) );
  NAND2X1 U64354 ( .A(n60028), .B(n60027), .Y(n60029) );
  NAND2X1 U64355 ( .A(n60030), .B(n60029), .Y(n60034) );
  XNOR2X1 U64356 ( .A(n60031), .B(n41869), .Y(n60032) );
  XNOR2X1 U64357 ( .A(n60033), .B(n60032), .Y(n60035) );
  INVX1 U64358 ( .A(n60035), .Y(n60092) );
  NAND2X1 U64359 ( .A(n60034), .B(n60092), .Y(n60039) );
  NAND2X1 U64360 ( .A(n43859), .B(n72820), .Y(n60093) );
  INVX1 U64361 ( .A(n60093), .Y(n60037) );
  INVX1 U64362 ( .A(n60034), .Y(n60094) );
  NAND2X1 U64363 ( .A(n60094), .B(n60035), .Y(n60036) );
  NAND2X1 U64364 ( .A(n60037), .B(n60036), .Y(n60038) );
  NAND2X1 U64365 ( .A(n60039), .B(n60038), .Y(n60040) );
  INVX1 U64366 ( .A(n60040), .Y(n60091) );
  INVX1 U64367 ( .A(n60089), .Y(n60041) );
  NAND2X1 U64368 ( .A(n60091), .B(n60041), .Y(n60042) );
  XNOR2X1 U64369 ( .A(n39230), .B(n60043), .Y(n60045) );
  XNOR2X1 U64370 ( .A(n60045), .B(n60044), .Y(n60046) );
  NAND2X1 U64371 ( .A(n36477), .B(n60046), .Y(n60050) );
  NAND2X1 U64372 ( .A(n72820), .B(n43955), .Y(n60087) );
  INVX1 U64373 ( .A(n60087), .Y(n60048) );
  INVX1 U64374 ( .A(n60046), .Y(n60086) );
  NAND2X1 U64375 ( .A(n39397), .B(n60086), .Y(n60047) );
  NAND2X1 U64376 ( .A(n60048), .B(n60047), .Y(n60049) );
  NAND2X1 U64377 ( .A(n60050), .B(n60049), .Y(n60051) );
  NAND2X1 U64378 ( .A(n60052), .B(n60051), .Y(n60054) );
  NAND2X1 U64379 ( .A(n43869), .B(n43810), .Y(n60083) );
  INVX1 U64380 ( .A(n60051), .Y(n60084) );
  INVX1 U64381 ( .A(n60052), .Y(n60082) );
  NAND2X1 U64382 ( .A(n60054), .B(n60055), .Y(n60169) );
  XNOR2X1 U64383 ( .A(n60061), .B(n60063), .Y(n60058) );
  XNOR2X1 U64384 ( .A(n60062), .B(n60061), .Y(n60064) );
  XNOR2X1 U64385 ( .A(n60064), .B(n60063), .Y(n60079) );
  XNOR2X1 U64386 ( .A(n60066), .B(n60065), .Y(n60068) );
  XNOR2X1 U64387 ( .A(n60068), .B(n60067), .Y(n60070) );
  INVX1 U64388 ( .A(n60070), .Y(n60076) );
  NAND2X1 U64389 ( .A(n60069), .B(n60076), .Y(n60074) );
  NAND2X1 U64390 ( .A(n43898), .B(n43810), .Y(n60077) );
  INVX1 U64391 ( .A(n60077), .Y(n60072) );
  NAND2X1 U64392 ( .A(n36478), .B(n60070), .Y(n60071) );
  NAND2X1 U64393 ( .A(n60072), .B(n60071), .Y(n60073) );
  NAND2X1 U64394 ( .A(n60074), .B(n60073), .Y(n60185) );
  INVX1 U64395 ( .A(n60185), .Y(n60189) );
  XNOR2X1 U64396 ( .A(n60075), .B(n60189), .Y(n60306) );
  XNOR2X1 U64397 ( .A(n60077), .B(n60076), .Y(n60078) );
  XNOR2X1 U64398 ( .A(n60078), .B(n36478), .Y(n60416) );
  INVX1 U64399 ( .A(n60175), .Y(n60310) );
  XNOR2X1 U64400 ( .A(n60083), .B(n60082), .Y(n60085) );
  XNOR2X1 U64401 ( .A(n60085), .B(n60084), .Y(n60166) );
  INVX1 U64402 ( .A(n60166), .Y(n60317) );
  XNOR2X1 U64403 ( .A(n60087), .B(n60086), .Y(n60088) );
  XNOR2X1 U64404 ( .A(n60088), .B(n39397), .Y(n60442) );
  INVX1 U64405 ( .A(n60442), .Y(n60319) );
  XNOR2X1 U64406 ( .A(n60089), .B(n41895), .Y(n60090) );
  XNOR2X1 U64407 ( .A(n60091), .B(n60090), .Y(n60322) );
  INVX1 U64408 ( .A(n60322), .Y(n60161) );
  XNOR2X1 U64409 ( .A(n60093), .B(n60092), .Y(n60095) );
  XNOR2X1 U64410 ( .A(n60095), .B(n60094), .Y(n60388) );
  XNOR2X1 U64411 ( .A(n60097), .B(n60096), .Y(n60099) );
  XNOR2X1 U64412 ( .A(n60099), .B(n60098), .Y(n60326) );
  INVX1 U64413 ( .A(n60326), .Y(n60152) );
  XNOR2X1 U64414 ( .A(n60100), .B(n38247), .Y(n60101) );
  XNOR2X1 U64415 ( .A(n60102), .B(n41835), .Y(n60103) );
  XNOR2X1 U64416 ( .A(n60104), .B(n60103), .Y(n60138) );
  INVX1 U64417 ( .A(n60138), .Y(n60370) );
  XNOR2X1 U64418 ( .A(n37395), .B(n60105), .Y(n60106) );
  XNOR2X1 U64419 ( .A(n60106), .B(n41807), .Y(n60131) );
  INVX1 U64420 ( .A(n60131), .Y(n60361) );
  XNOR2X1 U64421 ( .A(n60108), .B(n60107), .Y(n60109) );
  XNOR2X1 U64422 ( .A(n60109), .B(n41769), .Y(n60118) );
  INVX1 U64423 ( .A(n60118), .Y(n60353) );
  NAND2X1 U64424 ( .A(n72825), .B(n42719), .Y(n60340) );
  NAND2X1 U64425 ( .A(n44070), .B(n43811), .Y(n60341) );
  INVX1 U64426 ( .A(n60342), .Y(n60337) );
  NAND2X1 U64427 ( .A(n60111), .B(n60110), .Y(n60113) );
  NAND2X1 U64428 ( .A(n60113), .B(n60112), .Y(n60338) );
  INVX1 U64429 ( .A(n60338), .Y(n60114) );
  NAND2X1 U64430 ( .A(n60337), .B(n60114), .Y(n60117) );
  NAND2X1 U64431 ( .A(n60342), .B(n60338), .Y(n60115) );
  NAND2X1 U64432 ( .A(n41772), .B(n60115), .Y(n60116) );
  NAND2X1 U64433 ( .A(n60117), .B(n60116), .Y(n60354) );
  NAND2X1 U64434 ( .A(n60353), .B(n60354), .Y(n60122) );
  INVX1 U64435 ( .A(n60354), .Y(n60119) );
  NAND2X1 U64436 ( .A(n60119), .B(n60118), .Y(n60120) );
  NAND2X1 U64437 ( .A(n41792), .B(n60120), .Y(n60121) );
  NAND2X1 U64438 ( .A(n60122), .B(n60121), .Y(n60335) );
  XNOR2X1 U64439 ( .A(n60124), .B(n60123), .Y(n60125) );
  XNOR2X1 U64440 ( .A(n60125), .B(n41785), .Y(n60126) );
  NAND2X1 U64441 ( .A(n60335), .B(n60126), .Y(n60130) );
  INVX1 U64442 ( .A(n60335), .Y(n60127) );
  INVX1 U64443 ( .A(n60126), .Y(n60334) );
  NAND2X1 U64444 ( .A(n60127), .B(n60334), .Y(n60128) );
  NAND2X1 U64445 ( .A(n41811), .B(n60128), .Y(n60129) );
  NAND2X1 U64446 ( .A(n38242), .B(n60131), .Y(n60132) );
  XNOR2X1 U64447 ( .A(n60134), .B(n60133), .Y(n60135) );
  XNOR2X1 U64448 ( .A(n60135), .B(n41819), .Y(n60136) );
  INVX1 U64449 ( .A(n60136), .Y(n60331) );
  NAND2X1 U64450 ( .A(n39685), .B(n60331), .Y(n60137) );
  INVX1 U64451 ( .A(n60368), .Y(n60139) );
  NAND2X1 U64452 ( .A(n60139), .B(n60138), .Y(n60140) );
  XNOR2X1 U64453 ( .A(n60141), .B(n41847), .Y(n60142) );
  XNOR2X1 U64454 ( .A(n60143), .B(n60142), .Y(n60144) );
  NAND2X1 U64455 ( .A(n39816), .B(n60144), .Y(n60148) );
  NAND2X1 U64456 ( .A(n43821), .B(n44037), .Y(n60329) );
  INVX1 U64457 ( .A(n60329), .Y(n60146) );
  INVX1 U64458 ( .A(n60144), .Y(n60328) );
  NAND2X1 U64459 ( .A(n40643), .B(n60328), .Y(n60145) );
  NAND2X1 U64460 ( .A(n60146), .B(n60145), .Y(n60147) );
  NAND2X1 U64461 ( .A(n60148), .B(n60147), .Y(n60149) );
  NAND2X1 U64462 ( .A(n43821), .B(n43853), .Y(n60378) );
  INVX1 U64463 ( .A(n60378), .Y(n60151) );
  INVX1 U64464 ( .A(n60149), .Y(n60379) );
  NAND2X1 U64465 ( .A(n60152), .B(n60154), .Y(n60156) );
  INVX1 U64466 ( .A(n60153), .Y(n60325) );
  NAND2X1 U64467 ( .A(n60156), .B(n60155), .Y(n60157) );
  NAND2X1 U64468 ( .A(n60388), .B(n60157), .Y(n60160) );
  INVX1 U64469 ( .A(n60388), .Y(n60158) );
  NAND2X1 U64470 ( .A(n60160), .B(n60159), .Y(n60162) );
  INVX1 U64471 ( .A(n60162), .Y(n60324) );
  NAND2X1 U64472 ( .A(n60324), .B(n60322), .Y(n60163) );
  NAND2X1 U64473 ( .A(n43869), .B(n43821), .Y(n60438) );
  INVX1 U64474 ( .A(n60438), .Y(n60165) );
  INVX1 U64475 ( .A(n60440), .Y(n60321) );
  NAND2X1 U64476 ( .A(n60317), .B(n39812), .Y(n60168) );
  NAND2X1 U64477 ( .A(n43821), .B(n43881), .Y(n60316) );
  NAND2X1 U64478 ( .A(n60168), .B(n60167), .Y(n60171) );
  NAND2X1 U64479 ( .A(n43821), .B(n43891), .Y(n60313) );
  INVX1 U64480 ( .A(n60313), .Y(n60174) );
  INVX1 U64481 ( .A(n60171), .Y(n60314) );
  INVX1 U64482 ( .A(n60172), .Y(n60312) );
  NAND2X1 U64483 ( .A(n60312), .B(n60314), .Y(n60173) );
  NAND2X1 U64484 ( .A(n60310), .B(n37983), .Y(n60179) );
  NAND2X1 U64485 ( .A(n43897), .B(n43821), .Y(n60309) );
  INVX1 U64486 ( .A(n60309), .Y(n60177) );
  NAND2X1 U64487 ( .A(n38486), .B(n60175), .Y(n60176) );
  NAND2X1 U64488 ( .A(n60177), .B(n60176), .Y(n60178) );
  NAND2X1 U64489 ( .A(n60179), .B(n60178), .Y(n60180) );
  INVX1 U64490 ( .A(n60180), .Y(n60418) );
  INVX1 U64491 ( .A(n60416), .Y(n60181) );
  NAND2X1 U64492 ( .A(n60418), .B(n60181), .Y(n60182) );
  NAND2X1 U64493 ( .A(n60306), .B(n60739), .Y(n60741) );
  NAND2X1 U64494 ( .A(n43911), .B(n43821), .Y(n60737) );
  INVX1 U64495 ( .A(n60737), .Y(n60740) );
  INVX1 U64496 ( .A(n60739), .Y(n60308) );
  INVX1 U64497 ( .A(n60306), .Y(n60738) );
  NAND2X1 U64498 ( .A(n60308), .B(n60738), .Y(n60183) );
  NAND2X1 U64499 ( .A(n60740), .B(n60183), .Y(n60184) );
  NAND2X1 U64500 ( .A(n60741), .B(n60184), .Y(n60735) );
  INVX1 U64501 ( .A(n60187), .Y(n60191) );
  NAND2X1 U64502 ( .A(n60189), .B(n60188), .Y(n60190) );
  INVX1 U64503 ( .A(n60573), .Y(n60893) );
  NAND2X1 U64504 ( .A(n40461), .B(n43905), .Y(n60729) );
  NAND2X1 U64505 ( .A(n43898), .B(n40475), .Y(n60723) );
  NAND2X1 U64506 ( .A(n43889), .B(n40487), .Y(n60720) );
  NAND2X1 U64507 ( .A(n43788), .B(n43881), .Y(n60918) );
  NAND2X1 U64508 ( .A(n38253), .B(n60192), .Y(n60915) );
  NAND2X1 U64509 ( .A(n60195), .B(n60194), .Y(n60196) );
  XNOR2X1 U64510 ( .A(n60918), .B(n41275), .Y(n60282) );
  NAND2X1 U64511 ( .A(n43724), .B(n43872), .Y(n60575) );
  NAND2X1 U64512 ( .A(n43952), .B(n42632), .Y(n60699) );
  NAND2X1 U64513 ( .A(n60198), .B(n60200), .Y(n60204) );
  INVX1 U64514 ( .A(n60199), .Y(n60202) );
  XNOR2X1 U64515 ( .A(n38728), .B(n42181), .Y(n60201) );
  NAND2X1 U64516 ( .A(n60204), .B(n60203), .Y(n60696) );
  NAND2X1 U64517 ( .A(n39900), .B(n60205), .Y(n60206) );
  INVX1 U64518 ( .A(n60208), .Y(n60211) );
  NAND2X1 U64519 ( .A(n40663), .B(n60209), .Y(n60210) );
  NAND2X1 U64520 ( .A(n40399), .B(n60213), .Y(n60214) );
  NOR2X1 U64521 ( .A(n60217), .B(n60216), .Y(n60220) );
  XNOR2X1 U64522 ( .A(n41678), .B(n41499), .Y(n60267) );
  NAND2X1 U64523 ( .A(n38378), .B(n43796), .Y(n60589) );
  INVX1 U64524 ( .A(n60589), .Y(n61018) );
  NAND2X1 U64525 ( .A(n43840), .B(n43776), .Y(n61010) );
  INVX1 U64526 ( .A(n61010), .Y(n60992) );
  XNOR2X1 U64527 ( .A(n61018), .B(n60992), .Y(n60251) );
  NAND2X1 U64528 ( .A(n39420), .B(n60223), .Y(n60632) );
  NAND2X1 U64529 ( .A(n39955), .B(n60253), .Y(n60224) );
  NAND2X1 U64530 ( .A(n60225), .B(n60224), .Y(n60630) );
  NAND2X1 U64531 ( .A(n60632), .B(n60630), .Y(n60637) );
  INVX1 U64532 ( .A(n60227), .Y(n60226) );
  NAND2X1 U64533 ( .A(n60228), .B(n60227), .Y(n60230) );
  XNOR2X1 U64534 ( .A(n39206), .B(n41749), .Y(n60229) );
  NAND2X1 U64535 ( .A(n39680), .B(n61193), .Y(n60232) );
  NAND2X1 U64536 ( .A(n71546), .B(n40390), .Y(n60231) );
  NAND2X1 U64537 ( .A(n60232), .B(n60231), .Y(n60233) );
  NOR2X1 U64538 ( .A(n60234), .B(n38211), .Y(n60237) );
  NOR2X1 U64539 ( .A(n38503), .B(n60235), .Y(n60236) );
  NOR2X1 U64540 ( .A(n60237), .B(n60236), .Y(n60239) );
  NAND2X1 U64541 ( .A(n42376), .B(n62895), .Y(n63194) );
  INVX1 U64542 ( .A(n63194), .Y(n62458) );
  NOR2X1 U64543 ( .A(n39192), .B(n44072), .Y(n60238) );
  NAND2X1 U64544 ( .A(n60239), .B(n60238), .Y(n60241) );
  NAND2X1 U64545 ( .A(n40522), .B(n71033), .Y(n60608) );
  INVX1 U64546 ( .A(n60608), .Y(n60605) );
  XNOR2X1 U64547 ( .A(n60241), .B(n60605), .Y(n60242) );
  XNOR2X1 U64548 ( .A(n39682), .B(n60242), .Y(n60618) );
  NAND2X1 U64549 ( .A(n70371), .B(n43466), .Y(n60244) );
  NAND2X1 U64550 ( .A(n63222), .B(n70671), .Y(n60622) );
  INVX1 U64551 ( .A(n60622), .Y(n60620) );
  XNOR2X1 U64552 ( .A(n60244), .B(n60620), .Y(n60245) );
  NAND2X1 U64553 ( .A(n39939), .B(n43479), .Y(n60635) );
  NOR2X1 U64554 ( .A(n43485), .B(n43476), .Y(n60249) );
  NAND2X1 U64555 ( .A(n39617), .B(n60247), .Y(n60248) );
  XNOR2X1 U64556 ( .A(n60635), .B(n40155), .Y(n60250) );
  INVX1 U64557 ( .A(n60648), .Y(n61009) );
  XNOR2X1 U64558 ( .A(n60251), .B(n61009), .Y(n60258) );
  INVX1 U64559 ( .A(n60252), .Y(n60645) );
  XNOR2X1 U64560 ( .A(n60254), .B(n60253), .Y(n60255) );
  XNOR2X1 U64561 ( .A(n39955), .B(n60255), .Y(n60643) );
  INVX1 U64562 ( .A(n60643), .Y(n60256) );
  NAND2X1 U64563 ( .A(n60645), .B(n38961), .Y(n61012) );
  NAND2X1 U64564 ( .A(n60256), .B(n38961), .Y(n61013) );
  NAND2X1 U64565 ( .A(n61012), .B(n38443), .Y(n60257) );
  NOR2X1 U64566 ( .A(n38240), .B(n60257), .Y(n60991) );
  XNOR2X1 U64567 ( .A(n60258), .B(n40009), .Y(n60660) );
  NAND2X1 U64568 ( .A(n60259), .B(n39271), .Y(n61008) );
  NAND2X1 U64569 ( .A(n61008), .B(n61007), .Y(n60588) );
  NAND2X1 U64570 ( .A(n44036), .B(n42709), .Y(n60664) );
  INVX1 U64571 ( .A(n60664), .Y(n60662) );
  XNOR2X1 U64572 ( .A(n60588), .B(n60662), .Y(n60261) );
  XNOR2X1 U64573 ( .A(n60660), .B(n60261), .Y(n60266) );
  NOR2X1 U64574 ( .A(n60264), .B(n40957), .Y(n60265) );
  XNOR2X1 U64575 ( .A(n60267), .B(n36787), .Y(n60268) );
  XNOR2X1 U64576 ( .A(n60584), .B(n60268), .Y(n60269) );
  XNOR2X1 U64577 ( .A(n39914), .B(n60269), .Y(n60683) );
  NAND2X1 U64578 ( .A(n40259), .B(n43964), .Y(n60687) );
  INVX1 U64579 ( .A(n60687), .Y(n60684) );
  XNOR2X1 U64580 ( .A(n60683), .B(n60684), .Y(n60270) );
  XNOR2X1 U64581 ( .A(n42835), .B(n60270), .Y(n60697) );
  INVX1 U64582 ( .A(n60697), .Y(n60694) );
  XNOR2X1 U64583 ( .A(n60575), .B(n36753), .Y(n60281) );
  NAND2X1 U64584 ( .A(n60276), .B(n60271), .Y(n60280) );
  INVX1 U64585 ( .A(n60272), .Y(n60278) );
  NAND2X1 U64586 ( .A(n60274), .B(n60273), .Y(n60275) );
  OR2X1 U64587 ( .A(n60276), .B(n60275), .Y(n60277) );
  NAND2X1 U64588 ( .A(n60278), .B(n60277), .Y(n60279) );
  NAND2X1 U64589 ( .A(n60280), .B(n60279), .Y(n60574) );
  INVX1 U64590 ( .A(n60574), .Y(n60577) );
  XNOR2X1 U64591 ( .A(n60281), .B(n60577), .Y(n60917) );
  INVX1 U64592 ( .A(n60917), .Y(n60708) );
  XNOR2X1 U64593 ( .A(n60282), .B(n60708), .Y(n60721) );
  INVX1 U64594 ( .A(n60721), .Y(n60719) );
  INVX1 U64595 ( .A(n60284), .Y(n60285) );
  NAND2X1 U64596 ( .A(n60286), .B(n60285), .Y(n60287) );
  XNOR2X1 U64597 ( .A(n60723), .B(n38289), .Y(n60297) );
  INVX1 U64598 ( .A(n60292), .Y(n60290) );
  INVX1 U64599 ( .A(n60291), .Y(n60296) );
  XNOR2X1 U64600 ( .A(n60297), .B(n39695), .Y(n60730) );
  INVX1 U64601 ( .A(n60730), .Y(n60728) );
  XNOR2X1 U64602 ( .A(n60729), .B(n60728), .Y(n60303) );
  INVX1 U64603 ( .A(n60299), .Y(n60301) );
  NAND2X1 U64604 ( .A(n60301), .B(n60300), .Y(n60302) );
  INVX1 U64605 ( .A(n60727), .Y(n60731) );
  XNOR2X1 U64606 ( .A(n60303), .B(n60731), .Y(n60571) );
  NAND2X1 U64607 ( .A(n43911), .B(n72820), .Y(n60570) );
  INVX1 U64608 ( .A(n60570), .Y(n60895) );
  XNOR2X1 U64609 ( .A(n60571), .B(n60895), .Y(n60304) );
  XNOR2X1 U64610 ( .A(n60893), .B(n60304), .Y(n60745) );
  XNOR2X1 U64611 ( .A(n60745), .B(n41977), .Y(n60305) );
  INVX1 U64612 ( .A(n60564), .Y(n60567) );
  XNOR2X1 U64613 ( .A(n60566), .B(n60567), .Y(n60428) );
  XNOR2X1 U64614 ( .A(n60306), .B(n60740), .Y(n60307) );
  XNOR2X1 U64615 ( .A(n60308), .B(n60307), .Y(n60425) );
  INVX1 U64616 ( .A(n60425), .Y(n60431) );
  XNOR2X1 U64617 ( .A(n60309), .B(n38486), .Y(n60311) );
  XNOR2X1 U64618 ( .A(n60311), .B(n60310), .Y(n60413) );
  XNOR2X1 U64619 ( .A(n60313), .B(n60312), .Y(n60315) );
  XNOR2X1 U64620 ( .A(n60315), .B(n60314), .Y(n60539) );
  INVX1 U64621 ( .A(n60539), .Y(n60407) );
  XNOR2X1 U64622 ( .A(n60316), .B(n40546), .Y(n60318) );
  XNOR2X1 U64623 ( .A(n60318), .B(n60317), .Y(n60532) );
  XNOR2X1 U64624 ( .A(n60438), .B(n60319), .Y(n60320) );
  XNOR2X1 U64625 ( .A(n60321), .B(n60320), .Y(n60401) );
  XNOR2X1 U64626 ( .A(n60322), .B(n41910), .Y(n60323) );
  XNOR2X1 U64627 ( .A(n60324), .B(n60323), .Y(n60523) );
  XNOR2X1 U64628 ( .A(n60326), .B(n60325), .Y(n60327) );
  XNOR2X1 U64629 ( .A(n36490), .B(n60327), .Y(n60512) );
  XNOR2X1 U64630 ( .A(n60329), .B(n60328), .Y(n60330) );
  XNOR2X1 U64631 ( .A(n60330), .B(n40643), .Y(n60503) );
  INVX1 U64632 ( .A(n60503), .Y(n60376) );
  XNOR2X1 U64633 ( .A(n60332), .B(n60331), .Y(n60333) );
  XNOR2X1 U64634 ( .A(n60333), .B(n41838), .Y(n60366) );
  INVX1 U64635 ( .A(n60366), .Y(n60494) );
  XNOR2X1 U64636 ( .A(n60335), .B(n60334), .Y(n60336) );
  XNOR2X1 U64637 ( .A(n60336), .B(n41811), .Y(n60359) );
  INVX1 U64638 ( .A(n60359), .Y(n60484) );
  XNOR2X1 U64639 ( .A(n60338), .B(n60337), .Y(n60339) );
  XNOR2X1 U64640 ( .A(n60339), .B(n41772), .Y(n60348) );
  INVX1 U64641 ( .A(n60348), .Y(n60474) );
  NAND2X1 U64642 ( .A(n42719), .B(n72780), .Y(n60461) );
  NAND2X1 U64643 ( .A(n72825), .B(n73384), .Y(n60462) );
  INVX1 U64644 ( .A(n60463), .Y(n60458) );
  NAND2X1 U64645 ( .A(n60341), .B(n60340), .Y(n60343) );
  NAND2X1 U64646 ( .A(n60343), .B(n60342), .Y(n60459) );
  INVX1 U64647 ( .A(n60459), .Y(n60344) );
  NAND2X1 U64648 ( .A(n60458), .B(n60344), .Y(n60347) );
  NAND2X1 U64649 ( .A(n60463), .B(n60459), .Y(n60345) );
  NAND2X1 U64650 ( .A(n41775), .B(n60345), .Y(n60346) );
  NAND2X1 U64651 ( .A(n60347), .B(n60346), .Y(n60475) );
  NAND2X1 U64652 ( .A(n60474), .B(n60475), .Y(n60352) );
  INVX1 U64653 ( .A(n60475), .Y(n60349) );
  NAND2X1 U64654 ( .A(n60349), .B(n60348), .Y(n60350) );
  NAND2X1 U64655 ( .A(n41793), .B(n60350), .Y(n60351) );
  NAND2X1 U64656 ( .A(n60352), .B(n60351), .Y(n60456) );
  XNOR2X1 U64657 ( .A(n60354), .B(n60353), .Y(n60355) );
  XNOR2X1 U64658 ( .A(n60355), .B(n41792), .Y(n60356) );
  INVX1 U64659 ( .A(n60456), .Y(n60357) );
  INVX1 U64660 ( .A(n60356), .Y(n60455) );
  NAND2X1 U64661 ( .A(n60357), .B(n60455), .Y(n60358) );
  NAND2X1 U64662 ( .A(n39601), .B(n60359), .Y(n60360) );
  XNOR2X1 U64663 ( .A(n60362), .B(n60361), .Y(n60363) );
  XNOR2X1 U64664 ( .A(n60363), .B(n41824), .Y(n60364) );
  INVX1 U64665 ( .A(n60364), .Y(n60453) );
  NAND2X1 U64666 ( .A(n38180), .B(n60366), .Y(n60367) );
  XNOR2X1 U64667 ( .A(n60368), .B(n41851), .Y(n60369) );
  XNOR2X1 U64668 ( .A(n60370), .B(n60369), .Y(n60371) );
  NAND2X1 U64669 ( .A(n60451), .B(n60371), .Y(n60375) );
  INVX1 U64670 ( .A(n60451), .Y(n60372) );
  INVX1 U64671 ( .A(n60371), .Y(n60450) );
  NAND2X1 U64672 ( .A(n60372), .B(n60450), .Y(n60373) );
  NAND2X1 U64673 ( .A(n41868), .B(n60373), .Y(n60374) );
  NAND2X1 U64674 ( .A(n60375), .B(n60374), .Y(n60377) );
  INVX1 U64675 ( .A(n60377), .Y(n60504) );
  XNOR2X1 U64676 ( .A(n60378), .B(n36749), .Y(n60380) );
  XNOR2X1 U64677 ( .A(n60380), .B(n60379), .Y(n60446) );
  NAND2X1 U64678 ( .A(n60448), .B(n60446), .Y(n60384) );
  NOR2X1 U64679 ( .A(n60446), .B(n60448), .Y(n60381) );
  NAND2X1 U64680 ( .A(n43859), .B(n43758), .Y(n60447) );
  OR2X1 U64681 ( .A(n60381), .B(n60447), .Y(n60382) );
  NAND2X1 U64682 ( .A(n60384), .B(n60382), .Y(n60511) );
  NAND2X1 U64683 ( .A(n43758), .B(n43964), .Y(n60513) );
  INVX1 U64684 ( .A(n60513), .Y(n60387) );
  INVX1 U64685 ( .A(n60382), .Y(n60383) );
  NOR2X1 U64686 ( .A(n60383), .B(n60512), .Y(n60385) );
  NAND2X1 U64687 ( .A(n60385), .B(n60384), .Y(n60386) );
  XNOR2X1 U64688 ( .A(n60388), .B(n41894), .Y(n60389) );
  XNOR2X1 U64689 ( .A(n36493), .B(n60389), .Y(n60390) );
  INVX1 U64690 ( .A(n60390), .Y(n60443) );
  NAND2X1 U64691 ( .A(n60444), .B(n60443), .Y(n60395) );
  INVX1 U64692 ( .A(n60444), .Y(n60391) );
  NAND2X1 U64693 ( .A(n60391), .B(n60390), .Y(n60392) );
  NAND2X1 U64694 ( .A(n41911), .B(n60392), .Y(n60393) );
  NAND2X1 U64695 ( .A(n60395), .B(n60393), .Y(n60522) );
  NAND2X1 U64696 ( .A(n43869), .B(n43758), .Y(n60524) );
  INVX1 U64697 ( .A(n60524), .Y(n60398) );
  INVX1 U64698 ( .A(n60393), .Y(n60394) );
  NOR2X1 U64699 ( .A(n60394), .B(n60523), .Y(n60396) );
  NAND2X1 U64700 ( .A(n60396), .B(n60395), .Y(n60397) );
  NAND2X1 U64701 ( .A(n60398), .B(n60397), .Y(n60399) );
  NAND2X1 U64702 ( .A(n60400), .B(n60399), .Y(n60436) );
  NAND2X1 U64703 ( .A(n60401), .B(n60436), .Y(n60403) );
  NAND2X1 U64704 ( .A(n43758), .B(n43881), .Y(n60437) );
  OR2X1 U64705 ( .A(n60402), .B(n60437), .Y(n60404) );
  NAND2X1 U64706 ( .A(n60403), .B(n60404), .Y(n60531) );
  NAND2X1 U64707 ( .A(n60404), .B(n60403), .Y(n60405) );
  OR2X1 U64708 ( .A(n60532), .B(n60405), .Y(n60406) );
  NAND2X1 U64709 ( .A(n60407), .B(n60408), .Y(n60411) );
  NAND2X1 U64710 ( .A(n38161), .B(n60539), .Y(n60409) );
  NAND2X1 U64711 ( .A(n41947), .B(n60409), .Y(n60410) );
  NAND2X1 U64712 ( .A(n60411), .B(n60410), .Y(n60412) );
  NAND2X1 U64713 ( .A(n43758), .B(n43905), .Y(n60546) );
  INVX1 U64714 ( .A(n60546), .Y(n60415) );
  INVX1 U64715 ( .A(n60413), .Y(n60545) );
  NAND2X1 U64716 ( .A(n36483), .B(n60545), .Y(n60414) );
  XNOR2X1 U64717 ( .A(n60416), .B(n41957), .Y(n60417) );
  XNOR2X1 U64718 ( .A(n60418), .B(n60417), .Y(n60419) );
  INVX1 U64719 ( .A(n60419), .Y(n60433) );
  NAND2X1 U64720 ( .A(n38566), .B(n60433), .Y(n60423) );
  NAND2X1 U64721 ( .A(n43911), .B(n43758), .Y(n60434) );
  INVX1 U64722 ( .A(n60434), .Y(n60421) );
  NAND2X1 U64723 ( .A(n39140), .B(n60419), .Y(n60420) );
  NAND2X1 U64724 ( .A(n60421), .B(n60420), .Y(n60422) );
  NAND2X1 U64725 ( .A(n60423), .B(n60422), .Y(n60424) );
  NAND2X1 U64726 ( .A(n43920), .B(n43758), .Y(n60430) );
  INVX1 U64727 ( .A(n60430), .Y(n60427) );
  INVX1 U64728 ( .A(n60424), .Y(n60429) );
  NAND2X1 U64729 ( .A(n60429), .B(n60425), .Y(n60426) );
  INVX1 U64730 ( .A(n60565), .Y(n60568) );
  XNOR2X1 U64731 ( .A(n60428), .B(n60568), .Y(n60749) );
  INVX1 U64732 ( .A(n60749), .Y(n60559) );
  XNOR2X1 U64733 ( .A(n60430), .B(n60429), .Y(n60432) );
  XNOR2X1 U64734 ( .A(n60432), .B(n60431), .Y(n60752) );
  XNOR2X1 U64735 ( .A(n60434), .B(n60433), .Y(n60435) );
  XNOR2X1 U64736 ( .A(n60435), .B(n39140), .Y(n60553) );
  XNOR2X1 U64737 ( .A(n60438), .B(n60437), .Y(n60439) );
  XOR2X1 U64738 ( .A(n39017), .B(n60439), .Y(n60441) );
  XNOR2X1 U64739 ( .A(n60444), .B(n60443), .Y(n60445) );
  XNOR2X1 U64740 ( .A(n60448), .B(n60447), .Y(n60449) );
  INVX1 U64741 ( .A(n60509), .Y(n60843) );
  XNOR2X1 U64742 ( .A(n60451), .B(n60450), .Y(n60452) );
  XNOR2X1 U64743 ( .A(n60452), .B(n41868), .Y(n60501) );
  INVX1 U64744 ( .A(n60501), .Y(n60781) );
  XNOR2X1 U64745 ( .A(n36789), .B(n60453), .Y(n60454) );
  XNOR2X1 U64746 ( .A(n60454), .B(n41840), .Y(n60490) );
  INVX1 U64747 ( .A(n60490), .Y(n60787) );
  XNOR2X1 U64748 ( .A(n60456), .B(n60455), .Y(n60457) );
  XNOR2X1 U64749 ( .A(n60457), .B(n41813), .Y(n60480) );
  INVX1 U64750 ( .A(n60480), .Y(n60792) );
  XNOR2X1 U64751 ( .A(n60459), .B(n60458), .Y(n60460) );
  XNOR2X1 U64752 ( .A(n60460), .B(n41775), .Y(n60469) );
  INVX1 U64753 ( .A(n60469), .Y(n60798) );
  NAND2X1 U64754 ( .A(n42715), .B(n72760), .Y(n60804) );
  NAND2X1 U64755 ( .A(n73384), .B(n72780), .Y(n60805) );
  INVX1 U64756 ( .A(n60806), .Y(n60801) );
  NAND2X1 U64757 ( .A(n60462), .B(n60461), .Y(n60464) );
  NAND2X1 U64758 ( .A(n60464), .B(n60463), .Y(n60802) );
  INVX1 U64759 ( .A(n60802), .Y(n60465) );
  NAND2X1 U64760 ( .A(n60801), .B(n60465), .Y(n60468) );
  NAND2X1 U64761 ( .A(n60802), .B(n60806), .Y(n60466) );
  NAND2X1 U64762 ( .A(n41776), .B(n60466), .Y(n60467) );
  NAND2X1 U64763 ( .A(n60468), .B(n60467), .Y(n60799) );
  NAND2X1 U64764 ( .A(n60798), .B(n60799), .Y(n60473) );
  INVX1 U64765 ( .A(n60799), .Y(n60470) );
  NAND2X1 U64766 ( .A(n60470), .B(n60469), .Y(n60471) );
  NAND2X1 U64767 ( .A(n41796), .B(n60471), .Y(n60472) );
  NAND2X1 U64768 ( .A(n60473), .B(n60472), .Y(n60796) );
  XNOR2X1 U64769 ( .A(n60475), .B(n60474), .Y(n60476) );
  XNOR2X1 U64770 ( .A(n60476), .B(n41793), .Y(n60477) );
  INVX1 U64771 ( .A(n60796), .Y(n60478) );
  INVX1 U64772 ( .A(n60477), .Y(n60795) );
  NAND2X1 U64773 ( .A(n60478), .B(n60795), .Y(n60479) );
  NAND2X1 U64774 ( .A(n60792), .B(n60793), .Y(n60483) );
  NAND2X1 U64775 ( .A(n39172), .B(n60480), .Y(n60481) );
  NAND2X1 U64776 ( .A(n41829), .B(n60481), .Y(n60482) );
  NAND2X1 U64777 ( .A(n60483), .B(n60482), .Y(n60790) );
  XNOR2X1 U64778 ( .A(n60485), .B(n60484), .Y(n60486) );
  XNOR2X1 U64779 ( .A(n60486), .B(n41825), .Y(n60487) );
  INVX1 U64780 ( .A(n60790), .Y(n60488) );
  INVX1 U64781 ( .A(n60487), .Y(n60789) );
  NAND2X1 U64782 ( .A(n60488), .B(n60789), .Y(n60489) );
  NAND2X1 U64783 ( .A(n60787), .B(n60788), .Y(n60493) );
  NAND2X1 U64784 ( .A(n39454), .B(n60490), .Y(n60491) );
  NAND2X1 U64785 ( .A(n41856), .B(n60491), .Y(n60492) );
  NAND2X1 U64786 ( .A(n60493), .B(n60492), .Y(n60498) );
  XNOR2X1 U64787 ( .A(n60495), .B(n60494), .Y(n60496) );
  XNOR2X1 U64788 ( .A(n60496), .B(n41855), .Y(n60784) );
  INVX1 U64789 ( .A(n60497), .Y(n60783) );
  INVX1 U64790 ( .A(n60498), .Y(n60785) );
  INVX1 U64791 ( .A(n60784), .Y(n60499) );
  NAND2X1 U64792 ( .A(n60785), .B(n60499), .Y(n60500) );
  NAND2X1 U64793 ( .A(n60501), .B(n40611), .Y(n60502) );
  XNOR2X1 U64794 ( .A(n60503), .B(n41878), .Y(n60505) );
  XNOR2X1 U64795 ( .A(n60505), .B(n60504), .Y(n60506) );
  INVX1 U64796 ( .A(n60779), .Y(n60507) );
  INVX1 U64797 ( .A(n60506), .Y(n60778) );
  NAND2X1 U64798 ( .A(n60507), .B(n60778), .Y(n60508) );
  NAND2X1 U64799 ( .A(n40067), .B(n60509), .Y(n60510) );
  INVX1 U64800 ( .A(n60514), .Y(n60775) );
  NAND2X1 U64801 ( .A(n60776), .B(n60775), .Y(n60517) );
  NAND2X1 U64802 ( .A(n36361), .B(n60514), .Y(n60515) );
  NAND2X1 U64803 ( .A(n41912), .B(n60515), .Y(n60516) );
  NAND2X1 U64804 ( .A(n60517), .B(n60516), .Y(n60518) );
  NAND2X1 U64805 ( .A(n60519), .B(n60518), .Y(n60521) );
  NAND2X1 U64806 ( .A(n43870), .B(n43736), .Y(n60772) );
  INVX1 U64807 ( .A(n60518), .Y(n60773) );
  NAND2X1 U64808 ( .A(n60521), .B(n60520), .Y(n60525) );
  NAND2X1 U64809 ( .A(n43736), .B(n43881), .Y(n60770) );
  INVX1 U64810 ( .A(n60770), .Y(n60527) );
  NAND2X1 U64811 ( .A(n37400), .B(n60768), .Y(n60530) );
  NAND2X1 U64812 ( .A(n41942), .B(n60528), .Y(n60529) );
  NAND2X1 U64813 ( .A(n60530), .B(n60529), .Y(n60534) );
  XNOR2X1 U64814 ( .A(n60532), .B(n41938), .Y(n60533) );
  NAND2X1 U64815 ( .A(n60534), .B(n36784), .Y(n60538) );
  NAND2X1 U64816 ( .A(n43897), .B(n43737), .Y(n60765) );
  INVX1 U64817 ( .A(n60765), .Y(n60536) );
  INVX1 U64818 ( .A(n60534), .Y(n60766) );
  NAND2X1 U64819 ( .A(n60536), .B(n60535), .Y(n60537) );
  NAND2X1 U64820 ( .A(n60538), .B(n60537), .Y(n60541) );
  XNOR2X1 U64821 ( .A(n60539), .B(n41947), .Y(n60540) );
  XNOR2X1 U64822 ( .A(n38161), .B(n60540), .Y(n60542) );
  NAND2X1 U64823 ( .A(n43735), .B(n43905), .Y(n60762) );
  INVX1 U64824 ( .A(n60762), .Y(n60544) );
  INVX1 U64825 ( .A(n60541), .Y(n60763) );
  INVX1 U64826 ( .A(n60542), .Y(n60761) );
  NAND2X1 U64827 ( .A(n60763), .B(n60761), .Y(n60543) );
  XNOR2X1 U64828 ( .A(n60546), .B(n60545), .Y(n60547) );
  XNOR2X1 U64829 ( .A(n60547), .B(n36483), .Y(n60549) );
  INVX1 U64830 ( .A(n60549), .Y(n60758) );
  NAND2X1 U64831 ( .A(n60548), .B(n60758), .Y(n60551) );
  NAND2X1 U64832 ( .A(n43911), .B(n43737), .Y(n60759) );
  NAND2X1 U64833 ( .A(n60551), .B(n60550), .Y(n60552) );
  NAND2X1 U64834 ( .A(n60553), .B(n60552), .Y(n60555) );
  NAND2X1 U64835 ( .A(n43920), .B(n43737), .Y(n60755) );
  INVX1 U64836 ( .A(n60552), .Y(n60756) );
  INVX1 U64837 ( .A(n60553), .Y(n60754) );
  NAND2X1 U64838 ( .A(n60555), .B(n60554), .Y(n60556) );
  INVX1 U64839 ( .A(n60752), .Y(n60557) );
  NAND2X1 U64840 ( .A(n36512), .B(n60557), .Y(n60558) );
  NAND2X1 U64841 ( .A(n60559), .B(n60560), .Y(n60563) );
  INVX1 U64842 ( .A(n60560), .Y(n60751) );
  NAND2X1 U64843 ( .A(n42006), .B(n60561), .Y(n60562) );
  NAND2X1 U64844 ( .A(n60563), .B(n60562), .Y(n60882) );
  NAND2X1 U64845 ( .A(n60565), .B(n60564), .Y(n61082) );
  NAND2X1 U64846 ( .A(n61082), .B(n61085), .Y(n61080) );
  NAND2X1 U64847 ( .A(n43758), .B(n43936), .Y(n61081) );
  NAND2X1 U64848 ( .A(n43926), .B(n43821), .Y(n60888) );
  XNOR2X1 U64849 ( .A(n60730), .B(n60727), .Y(n60569) );
  XOR2X1 U64850 ( .A(n60729), .B(n60569), .Y(n60892) );
  NOR2X1 U64851 ( .A(n60892), .B(n60570), .Y(n60572) );
  NAND2X1 U64852 ( .A(n43910), .B(n40464), .Y(n60900) );
  NAND2X1 U64853 ( .A(n43897), .B(n40488), .Y(n61074) );
  NAND2X1 U64854 ( .A(n43724), .B(n43881), .Y(n61256) );
  NAND2X1 U64855 ( .A(n36753), .B(n60574), .Y(n60581) );
  INVX1 U64856 ( .A(n60575), .Y(n60579) );
  NAND2X1 U64857 ( .A(n60577), .B(n60576), .Y(n60578) );
  NAND2X1 U64858 ( .A(n60579), .B(n60578), .Y(n60580) );
  NAND2X1 U64859 ( .A(n60581), .B(n60580), .Y(n60925) );
  XNOR2X1 U64860 ( .A(n61256), .B(n39341), .Y(n60707) );
  NAND2X1 U64861 ( .A(n43798), .B(n43964), .Y(n61044) );
  NAND2X1 U64862 ( .A(n39914), .B(n40620), .Y(n60583) );
  XNOR2X1 U64863 ( .A(n39219), .B(n61044), .Y(n60682) );
  NAND2X1 U64864 ( .A(n42658), .B(n43862), .Y(n61036) );
  XNOR2X1 U64865 ( .A(n61036), .B(n38957), .Y(n60681) );
  NAND2X1 U64866 ( .A(n44035), .B(n43796), .Y(n61006) );
  XNOR2X1 U64867 ( .A(n61010), .B(n61009), .Y(n60586) );
  XNOR2X1 U64868 ( .A(n40009), .B(n60586), .Y(n60587) );
  NOR2X1 U64869 ( .A(n60587), .B(n60589), .Y(n60592) );
  INVX1 U64870 ( .A(n60588), .Y(n60661) );
  OR2X1 U64871 ( .A(n60661), .B(n60589), .Y(n60590) );
  NAND2X1 U64872 ( .A(n61019), .B(n60590), .Y(n60591) );
  NOR2X1 U64873 ( .A(n60592), .B(n60591), .Y(n61002) );
  NAND2X1 U64874 ( .A(n43840), .B(n43479), .Y(n60985) );
  NAND2X1 U64875 ( .A(n39942), .B(n43483), .Y(n61203) );
  XNOR2X1 U64876 ( .A(n60617), .B(n60620), .Y(n60593) );
  XNOR2X1 U64877 ( .A(n38856), .B(n60593), .Y(n60597) );
  INVX1 U64878 ( .A(n60597), .Y(n60594) );
  NOR2X1 U64879 ( .A(n40614), .B(n60594), .Y(n60595) );
  XNOR2X1 U64880 ( .A(n61203), .B(n39614), .Y(n60629) );
  NAND2X1 U64881 ( .A(n62659), .B(n71297), .Y(n60939) );
  NAND2X1 U64882 ( .A(n60945), .B(n63194), .Y(n60598) );
  NAND2X1 U64883 ( .A(n60958), .B(n61185), .Y(n60599) );
  INVX1 U64884 ( .A(n60935), .Y(n61173) );
  NAND2X1 U64885 ( .A(n60598), .B(n60599), .Y(n60936) );
  INVX1 U64886 ( .A(n60936), .Y(n60600) );
  NOR2X1 U64887 ( .A(n61173), .B(n60600), .Y(n60601) );
  XNOR2X1 U64888 ( .A(n60939), .B(n60601), .Y(n60604) );
  NAND2X1 U64889 ( .A(n37361), .B(n71546), .Y(n60602) );
  NOR2X1 U64890 ( .A(n43499), .B(n60602), .Y(n60603) );
  XNOR2X1 U64891 ( .A(n60604), .B(n60603), .Y(n61148) );
  NAND2X1 U64892 ( .A(n60606), .B(n60605), .Y(n60970) );
  NAND2X1 U64893 ( .A(n60970), .B(n61147), .Y(n60609) );
  NAND2X1 U64894 ( .A(n60608), .B(n60607), .Y(n60610) );
  NAND2X1 U64895 ( .A(n39682), .B(n60610), .Y(n60969) );
  NOR2X1 U64896 ( .A(n60609), .B(n60611), .Y(n60615) );
  OR2X1 U64897 ( .A(n61147), .B(n60970), .Y(n60613) );
  INVX1 U64898 ( .A(n61147), .Y(n60972) );
  NAND2X1 U64899 ( .A(n60611), .B(n60972), .Y(n60612) );
  NAND2X1 U64900 ( .A(n60613), .B(n60612), .Y(n60614) );
  NOR2X1 U64901 ( .A(n60615), .B(n60614), .Y(n60616) );
  XOR2X1 U64902 ( .A(n61148), .B(n60616), .Y(n60934) );
  NAND2X1 U64903 ( .A(n43464), .B(n43488), .Y(n60932) );
  NAND2X1 U64904 ( .A(n60932), .B(n39681), .Y(n60621) );
  INVX1 U64905 ( .A(n60617), .Y(n60619) );
  NAND2X1 U64906 ( .A(n60619), .B(n60618), .Y(n60623) );
  NOR2X1 U64907 ( .A(n39571), .B(n60621), .Y(n60628) );
  OR2X1 U64908 ( .A(n60932), .B(n60930), .Y(n60626) );
  NOR2X1 U64909 ( .A(n60622), .B(n60932), .Y(n60624) );
  NAND2X1 U64910 ( .A(n60624), .B(n60623), .Y(n60625) );
  NAND2X1 U64911 ( .A(n60626), .B(n60625), .Y(n60627) );
  INVX1 U64912 ( .A(n39238), .Y(n60975) );
  XNOR2X1 U64913 ( .A(n60629), .B(n60975), .Y(n60986) );
  INVX1 U64914 ( .A(n60986), .Y(n60982) );
  XNOR2X1 U64915 ( .A(n60985), .B(n60982), .Y(n60642) );
  INVX1 U64916 ( .A(n60630), .Y(n60634) );
  NAND2X1 U64917 ( .A(n60632), .B(n60638), .Y(n60633) );
  NOR2X1 U64918 ( .A(n60634), .B(n60633), .Y(n60636) );
  NOR2X1 U64919 ( .A(n60636), .B(n60635), .Y(n60641) );
  INVX1 U64920 ( .A(n60637), .Y(n60639) );
  NOR2X1 U64921 ( .A(n60639), .B(n60638), .Y(n60640) );
  XNOR2X1 U64922 ( .A(n60642), .B(n38517), .Y(n60998) );
  NAND2X1 U64923 ( .A(n39892), .B(n60643), .Y(n60644) );
  NAND2X1 U64924 ( .A(n60645), .B(n60644), .Y(n60646) );
  NAND2X1 U64925 ( .A(n60646), .B(n61013), .Y(n60649) );
  INVX1 U64926 ( .A(n60652), .Y(n60647) );
  NOR2X1 U64927 ( .A(n61010), .B(n60647), .Y(n60651) );
  NAND2X1 U64928 ( .A(n60649), .B(n60648), .Y(n60993) );
  NAND2X1 U64929 ( .A(n38379), .B(n43776), .Y(n60997) );
  NAND2X1 U64930 ( .A(n60993), .B(n60997), .Y(n60650) );
  NOR2X1 U64931 ( .A(n60651), .B(n60650), .Y(n60657) );
  OR2X1 U64932 ( .A(n60997), .B(n60993), .Y(n60655) );
  NOR2X1 U64933 ( .A(n61010), .B(n60997), .Y(n60653) );
  NAND2X1 U64934 ( .A(n60653), .B(n60652), .Y(n60654) );
  NAND2X1 U64935 ( .A(n60655), .B(n60654), .Y(n60656) );
  INVX1 U64936 ( .A(n61032), .Y(n61029) );
  NOR2X1 U64937 ( .A(n60662), .B(n40957), .Y(n60659) );
  NAND2X1 U64938 ( .A(n41359), .B(n60665), .Y(n60658) );
  NAND2X1 U64939 ( .A(n60659), .B(n60658), .Y(n60674) );
  NAND2X1 U64940 ( .A(n60674), .B(n60672), .Y(n61026) );
  INVX1 U64941 ( .A(n61026), .Y(n60670) );
  NAND2X1 U64942 ( .A(n40957), .B(n60662), .Y(n60668) );
  NOR2X1 U64943 ( .A(n60664), .B(n60663), .Y(n60666) );
  NAND2X1 U64944 ( .A(n60666), .B(n60665), .Y(n60667) );
  NAND2X1 U64945 ( .A(n60668), .B(n60667), .Y(n60671) );
  INVX1 U64946 ( .A(n60671), .Y(n61027) );
  NAND2X1 U64947 ( .A(n43851), .B(n42708), .Y(n61028) );
  NAND2X1 U64948 ( .A(n61027), .B(n61028), .Y(n60669) );
  NOR2X1 U64949 ( .A(n60670), .B(n60669), .Y(n60679) );
  INVX1 U64950 ( .A(n61028), .Y(n61033) );
  NAND2X1 U64951 ( .A(n61033), .B(n60671), .Y(n60677) );
  INVX1 U64952 ( .A(n60672), .Y(n60673) );
  NOR2X1 U64953 ( .A(n60673), .B(n61028), .Y(n60675) );
  NAND2X1 U64954 ( .A(n60675), .B(n60674), .Y(n60676) );
  NAND2X1 U64955 ( .A(n60677), .B(n60676), .Y(n60678) );
  NOR2X1 U64956 ( .A(n60679), .B(n60678), .Y(n60680) );
  XNOR2X1 U64957 ( .A(n61029), .B(n60680), .Y(n61035) );
  INVX1 U64958 ( .A(n61035), .Y(n61037) );
  XNOR2X1 U64959 ( .A(n60681), .B(n61037), .Y(n61045) );
  INVX1 U64960 ( .A(n61045), .Y(n61043) );
  XNOR2X1 U64961 ( .A(n60682), .B(n61043), .Y(n61056) );
  INVX1 U64962 ( .A(n61056), .Y(n61052) );
  NAND2X1 U64963 ( .A(n40260), .B(n43954), .Y(n61055) );
  NAND2X1 U64964 ( .A(n61049), .B(n61055), .Y(n60686) );
  NAND2X1 U64965 ( .A(n42835), .B(n60683), .Y(n60688) );
  NAND2X1 U64966 ( .A(n60684), .B(n60688), .Y(n61048) );
  INVX1 U64967 ( .A(n61048), .Y(n60685) );
  NOR2X1 U64968 ( .A(n60686), .B(n60685), .Y(n60693) );
  OR2X1 U64969 ( .A(n61055), .B(n61049), .Y(n60691) );
  NOR2X1 U64970 ( .A(n60687), .B(n61055), .Y(n60689) );
  NAND2X1 U64971 ( .A(n60689), .B(n60688), .Y(n60690) );
  NAND2X1 U64972 ( .A(n60691), .B(n60690), .Y(n60692) );
  INVX1 U64973 ( .A(n60699), .Y(n60695) );
  NAND2X1 U64974 ( .A(n39205), .B(n60694), .Y(n60700) );
  NAND2X1 U64975 ( .A(n60695), .B(n60700), .Y(n61061) );
  NAND2X1 U64976 ( .A(n60697), .B(n60696), .Y(n61062) );
  NAND2X1 U64977 ( .A(n43869), .B(n42632), .Y(n61060) );
  NAND2X1 U64978 ( .A(n61062), .B(n61060), .Y(n60698) );
  NOR2X1 U64979 ( .A(n39336), .B(n60698), .Y(n60705) );
  INVX1 U64980 ( .A(n61060), .Y(n61067) );
  NOR2X1 U64981 ( .A(n60699), .B(n61060), .Y(n60701) );
  NAND2X1 U64982 ( .A(n60701), .B(n60700), .Y(n60702) );
  NAND2X1 U64983 ( .A(n60703), .B(n60702), .Y(n60704) );
  NOR2X1 U64984 ( .A(n60705), .B(n60704), .Y(n60706) );
  XNOR2X1 U64985 ( .A(n61063), .B(n60706), .Y(n60926) );
  INVX1 U64986 ( .A(n60926), .Y(n60927) );
  XNOR2X1 U64987 ( .A(n60707), .B(n60927), .Y(n60921) );
  INVX1 U64988 ( .A(n60921), .Y(n60913) );
  INVX1 U64989 ( .A(n60918), .Y(n60709) );
  NAND2X1 U64990 ( .A(n60709), .B(n60712), .Y(n60910) );
  NOR2X1 U64991 ( .A(n39713), .B(n60710), .Y(n60717) );
  INVX1 U64992 ( .A(n60711), .Y(n60924) );
  NAND2X1 U64993 ( .A(n39569), .B(n60924), .Y(n60715) );
  NOR2X1 U64994 ( .A(n60918), .B(n60711), .Y(n60713) );
  NAND2X1 U64995 ( .A(n60713), .B(n60712), .Y(n60714) );
  NAND2X1 U64996 ( .A(n60715), .B(n60714), .Y(n60716) );
  NOR2X1 U64997 ( .A(n60717), .B(n60716), .Y(n60718) );
  XNOR2X1 U64998 ( .A(n60913), .B(n60718), .Y(n61075) );
  INVX1 U64999 ( .A(n61075), .Y(n61072) );
  XNOR2X1 U65000 ( .A(n61074), .B(n61072), .Y(n60722) );
  XNOR2X1 U65001 ( .A(n60722), .B(n36686), .Y(n60907) );
  NAND2X1 U65002 ( .A(n40476), .B(n43905), .Y(n60904) );
  NAND2X1 U65003 ( .A(n36568), .B(n60724), .Y(n60903) );
  NAND2X1 U65004 ( .A(n60902), .B(n60903), .Y(n60725) );
  XNOR2X1 U65005 ( .A(n60907), .B(n60726), .Y(n60901) );
  INVX1 U65006 ( .A(n60901), .Y(n60899) );
  INVX1 U65007 ( .A(n60729), .Y(n60733) );
  NAND2X1 U65008 ( .A(n43920), .B(n43810), .Y(n61105) );
  INVX1 U65009 ( .A(n61105), .Y(n60896) );
  XNOR2X1 U65010 ( .A(n61108), .B(n60896), .Y(n60734) );
  INVX1 U65011 ( .A(n60889), .Y(n60886) );
  INVX1 U65012 ( .A(n60745), .Y(n60736) );
  NOR2X1 U65013 ( .A(n60738), .B(n60737), .Y(n60744) );
  NAND2X1 U65014 ( .A(n60740), .B(n60739), .Y(n60742) );
  NAND2X1 U65015 ( .A(n60742), .B(n60741), .Y(n60743) );
  NOR2X1 U65016 ( .A(n60744), .B(n60743), .Y(n60746) );
  NAND2X1 U65017 ( .A(n60746), .B(n60745), .Y(n60747) );
  XNOR2X1 U65018 ( .A(n60884), .B(n42015), .Y(n60748) );
  XNOR2X1 U65019 ( .A(n36628), .B(n60748), .Y(n61431) );
  XNOR2X1 U65020 ( .A(n60749), .B(n42006), .Y(n60750) );
  XNOR2X1 U65021 ( .A(n60751), .B(n60750), .Y(n61302) );
  XNOR2X1 U65022 ( .A(n60752), .B(n41991), .Y(n60753) );
  XNOR2X1 U65023 ( .A(n36512), .B(n60753), .Y(n61304) );
  INVX1 U65024 ( .A(n61304), .Y(n60875) );
  XNOR2X1 U65025 ( .A(n60755), .B(n60754), .Y(n60757) );
  XNOR2X1 U65026 ( .A(n60757), .B(n60756), .Y(n61306) );
  INVX1 U65027 ( .A(n61306), .Y(n60872) );
  XNOR2X1 U65028 ( .A(n60759), .B(n60758), .Y(n60760) );
  XNOR2X1 U65029 ( .A(n60760), .B(n38268), .Y(n61308) );
  XNOR2X1 U65030 ( .A(n60762), .B(n60761), .Y(n60764) );
  XNOR2X1 U65031 ( .A(n60764), .B(n60763), .Y(n61310) );
  INVX1 U65032 ( .A(n61310), .Y(n60867) );
  XNOR2X1 U65033 ( .A(n60765), .B(n36784), .Y(n60767) );
  XNOR2X1 U65034 ( .A(n60767), .B(n60766), .Y(n61313) );
  XNOR2X1 U65035 ( .A(n60768), .B(n37400), .Y(n60769) );
  XNOR2X1 U65036 ( .A(n60769), .B(n41942), .Y(n61316) );
  XNOR2X1 U65037 ( .A(n60770), .B(n37403), .Y(n60771) );
  XNOR2X1 U65038 ( .A(n60771), .B(n36460), .Y(n61318) );
  XNOR2X1 U65039 ( .A(n60772), .B(n38244), .Y(n60774) );
  XNOR2X1 U65040 ( .A(n60774), .B(n60773), .Y(n61320) );
  INVX1 U65041 ( .A(n61320), .Y(n60850) );
  XNOR2X1 U65042 ( .A(n60776), .B(n60775), .Y(n60777) );
  XNOR2X1 U65043 ( .A(n60777), .B(n41912), .Y(n61322) );
  XNOR2X1 U65044 ( .A(n60779), .B(n60778), .Y(n60780) );
  XNOR2X1 U65045 ( .A(n60780), .B(n41889), .Y(n61327) );
  INVX1 U65046 ( .A(n61327), .Y(n60840) );
  XNOR2X1 U65047 ( .A(n39694), .B(n60781), .Y(n60782) );
  XNOR2X1 U65048 ( .A(n60782), .B(n41879), .Y(n61329) );
  XNOR2X1 U65049 ( .A(n60784), .B(n60783), .Y(n60786) );
  XNOR2X1 U65050 ( .A(n60786), .B(n60785), .Y(n61331) );
  INVX1 U65051 ( .A(n61331), .Y(n60835) );
  XNOR2X1 U65052 ( .A(n60790), .B(n60789), .Y(n60791) );
  XNOR2X1 U65053 ( .A(n60791), .B(n41841), .Y(n61335) );
  INVX1 U65054 ( .A(n61335), .Y(n60830) );
  XNOR2X1 U65055 ( .A(n60793), .B(n60792), .Y(n60794) );
  XNOR2X1 U65056 ( .A(n60794), .B(n41829), .Y(n61339) );
  XNOR2X1 U65057 ( .A(n60796), .B(n60795), .Y(n60797) );
  XNOR2X1 U65058 ( .A(n60797), .B(n41814), .Y(n61341) );
  INVX1 U65059 ( .A(n61341), .Y(n60820) );
  XNOR2X1 U65060 ( .A(n60799), .B(n60798), .Y(n60800) );
  XNOR2X1 U65061 ( .A(n60800), .B(n41796), .Y(n61344) );
  XNOR2X1 U65062 ( .A(n60802), .B(n60801), .Y(n60803) );
  XNOR2X1 U65063 ( .A(n60803), .B(n41776), .Y(n61347) );
  INVX1 U65064 ( .A(n61347), .Y(n60812) );
  NAND2X1 U65065 ( .A(n42719), .B(n43782), .Y(n61352) );
  NAND2X1 U65066 ( .A(n44070), .B(n72760), .Y(n61353) );
  INVX1 U65067 ( .A(n61354), .Y(n61349) );
  NAND2X1 U65068 ( .A(n60805), .B(n60804), .Y(n60807) );
  NAND2X1 U65069 ( .A(n60807), .B(n60806), .Y(n61350) );
  INVX1 U65070 ( .A(n61350), .Y(n60808) );
  NAND2X1 U65071 ( .A(n61349), .B(n60808), .Y(n60811) );
  NAND2X1 U65072 ( .A(n61350), .B(n61354), .Y(n60809) );
  NAND2X1 U65073 ( .A(n41781), .B(n60809), .Y(n60810) );
  NAND2X1 U65074 ( .A(n60811), .B(n60810), .Y(n60813) );
  NAND2X1 U65075 ( .A(n60812), .B(n60813), .Y(n60816) );
  INVX1 U65076 ( .A(n60813), .Y(n61346) );
  NAND2X1 U65077 ( .A(n61346), .B(n61347), .Y(n60814) );
  NAND2X1 U65078 ( .A(n41799), .B(n60814), .Y(n60815) );
  NAND2X1 U65079 ( .A(n60816), .B(n60815), .Y(n60817) );
  INVX1 U65080 ( .A(n60817), .Y(n61343) );
  INVX1 U65081 ( .A(n61344), .Y(n60818) );
  NAND2X1 U65082 ( .A(n61343), .B(n60818), .Y(n60819) );
  NAND2X1 U65083 ( .A(n60820), .B(n60821), .Y(n60824) );
  NAND2X1 U65084 ( .A(n38915), .B(n61341), .Y(n60822) );
  NAND2X1 U65085 ( .A(n41831), .B(n60822), .Y(n60823) );
  NAND2X1 U65086 ( .A(n60824), .B(n60823), .Y(n60825) );
  NAND2X1 U65087 ( .A(n61339), .B(n60825), .Y(n60829) );
  INVX1 U65088 ( .A(n60825), .Y(n61338) );
  INVX1 U65089 ( .A(n61339), .Y(n60826) );
  NAND2X1 U65090 ( .A(n61338), .B(n60826), .Y(n60827) );
  NAND2X1 U65091 ( .A(n41844), .B(n60827), .Y(n60828) );
  NAND2X1 U65092 ( .A(n60829), .B(n60828), .Y(n60831) );
  INVX1 U65093 ( .A(n60831), .Y(n61337) );
  NAND2X1 U65094 ( .A(n61337), .B(n61335), .Y(n60832) );
  NAND2X1 U65095 ( .A(n39675), .B(n38219), .Y(n60834) );
  NAND2X1 U65096 ( .A(n39149), .B(n61331), .Y(n60837) );
  INVX1 U65097 ( .A(n61329), .Y(n60838) );
  NAND2X1 U65098 ( .A(n40243), .B(n60838), .Y(n60839) );
  NAND2X1 U65099 ( .A(n39098), .B(n61327), .Y(n60841) );
  XNOR2X1 U65100 ( .A(n38618), .B(n41901), .Y(n60842) );
  XNOR2X1 U65101 ( .A(n60843), .B(n60842), .Y(n60844) );
  INVX1 U65102 ( .A(n61324), .Y(n60845) );
  INVX1 U65103 ( .A(n60844), .Y(n61326) );
  NAND2X1 U65104 ( .A(n60845), .B(n61326), .Y(n60846) );
  INVX1 U65105 ( .A(n61322), .Y(n60848) );
  NAND2X1 U65106 ( .A(n40632), .B(n60848), .Y(n60849) );
  NAND2X1 U65107 ( .A(n60850), .B(n60851), .Y(n60854) );
  NAND2X1 U65108 ( .A(n39441), .B(n61320), .Y(n60852) );
  NAND2X1 U65109 ( .A(n41932), .B(n60852), .Y(n60853) );
  NAND2X1 U65110 ( .A(n60854), .B(n60853), .Y(n60855) );
  INVX1 U65111 ( .A(n61318), .Y(n60856) );
  NAND2X1 U65112 ( .A(n38150), .B(n60856), .Y(n60857) );
  NAND2X1 U65113 ( .A(n61316), .B(n60858), .Y(n60862) );
  INVX1 U65114 ( .A(n61316), .Y(n60859) );
  NAND2X1 U65115 ( .A(n36461), .B(n60859), .Y(n60860) );
  NAND2X1 U65116 ( .A(n41953), .B(n60860), .Y(n60861) );
  NAND2X1 U65117 ( .A(n60862), .B(n60861), .Y(n60863) );
  NAND2X1 U65118 ( .A(n61313), .B(n60863), .Y(n60866) );
  INVX1 U65119 ( .A(n60863), .Y(n61315) );
  NAND2X1 U65120 ( .A(n41962), .B(n60864), .Y(n60865) );
  NAND2X1 U65121 ( .A(n60866), .B(n60865), .Y(n60868) );
  INVX1 U65122 ( .A(n60868), .Y(n61312) );
  NAND2X1 U65123 ( .A(n61312), .B(n61310), .Y(n60869) );
  INVX1 U65124 ( .A(n61308), .Y(n60870) );
  NAND2X1 U65125 ( .A(n40357), .B(n60870), .Y(n60871) );
  NAND2X1 U65126 ( .A(n37888), .B(n61306), .Y(n60874) );
  NAND2X1 U65127 ( .A(n40549), .B(n61304), .Y(n60876) );
  INVX1 U65128 ( .A(n61302), .Y(n60878) );
  NAND2X1 U65129 ( .A(n39999), .B(n60878), .Y(n60879) );
  INVX1 U65130 ( .A(n61431), .Y(n60880) );
  NAND2X1 U65131 ( .A(n60880), .B(n37891), .Y(n60881) );
  INVX1 U65132 ( .A(n60884), .Y(n60883) );
  NAND2X1 U65133 ( .A(n36628), .B(n60884), .Y(n60885) );
  NAND2X1 U65134 ( .A(n43758), .B(n43944), .Y(n62356) );
  NAND2X1 U65135 ( .A(n43821), .B(n43935), .Y(n61101) );
  INVX1 U65136 ( .A(n60888), .Y(n60891) );
  NAND2X1 U65137 ( .A(n39387), .B(n60889), .Y(n60890) );
  XNOR2X1 U65138 ( .A(n61101), .B(n38645), .Y(n61079) );
  NAND2X1 U65139 ( .A(n61108), .B(n61110), .Y(n60898) );
  NAND2X1 U65140 ( .A(n60893), .B(n60892), .Y(n60894) );
  NAND2X1 U65141 ( .A(n60896), .B(n61106), .Y(n60897) );
  NAND2X1 U65142 ( .A(n60898), .B(n60897), .Y(n61117) );
  NAND2X1 U65143 ( .A(n43919), .B(n40465), .Y(n61103) );
  NAND2X1 U65144 ( .A(n43926), .B(n72820), .Y(n61109) );
  XNOR2X1 U65145 ( .A(n61103), .B(n61109), .Y(n61078) );
  NAND2X1 U65146 ( .A(n38472), .B(n60899), .Y(n61290) );
  NAND2X1 U65147 ( .A(n61290), .B(n61289), .Y(n61295) );
  NAND2X1 U65148 ( .A(n43910), .B(n40470), .Y(n61285) );
  NAND2X1 U65149 ( .A(n60903), .B(n60902), .Y(n60906) );
  NOR2X1 U65150 ( .A(n60907), .B(n60906), .Y(n60905) );
  INVX1 U65151 ( .A(n60906), .Y(n60909) );
  INVX1 U65152 ( .A(n60907), .Y(n60908) );
  XNOR2X1 U65153 ( .A(n61285), .B(n38885), .Y(n61076) );
  NAND2X1 U65154 ( .A(n40489), .B(n43905), .Y(n61275) );
  NAND2X1 U65155 ( .A(n60911), .B(n60910), .Y(n60912) );
  NAND2X1 U65156 ( .A(n60915), .B(n60914), .Y(n60916) );
  NOR2X1 U65157 ( .A(n60917), .B(n60916), .Y(n60919) );
  NOR2X1 U65158 ( .A(n60919), .B(n60918), .Y(n60920) );
  NOR2X1 U65159 ( .A(n39569), .B(n60920), .Y(n60922) );
  NAND2X1 U65160 ( .A(n60922), .B(n60921), .Y(n60923) );
  NAND2X1 U65161 ( .A(n43724), .B(n43891), .Y(n61255) );
  XNOR2X1 U65162 ( .A(n61255), .B(n41930), .Y(n60929) );
  NAND2X1 U65163 ( .A(n60926), .B(n60925), .Y(n61254) );
  INVX1 U65164 ( .A(n61256), .Y(n60928) );
  NAND2X1 U65165 ( .A(n39341), .B(n60927), .Y(n61257) );
  NAND2X1 U65166 ( .A(n60928), .B(n61257), .Y(n61251) );
  XNOR2X1 U65167 ( .A(n60929), .B(n42841), .Y(n61069) );
  NAND2X1 U65168 ( .A(n43879), .B(n42632), .Y(n61240) );
  NAND2X1 U65169 ( .A(n40259), .B(n43872), .Y(n61121) );
  NAND2X1 U65170 ( .A(n43798), .B(n43954), .Y(n61234) );
  NAND2X1 U65171 ( .A(n42659), .B(n43964), .Y(n61128) );
  NAND2X1 U65172 ( .A(n43859), .B(n42714), .Y(n61226) );
  NAND2X1 U65173 ( .A(n43851), .B(n43796), .Y(n61221) );
  NAND2X1 U65174 ( .A(n44036), .B(n43776), .Y(n61131) );
  NAND2X1 U65175 ( .A(n38380), .B(n43479), .Y(n61217) );
  INVX1 U65176 ( .A(n60934), .Y(n60931) );
  NAND2X1 U65177 ( .A(n60933), .B(n60931), .Y(n61141) );
  NAND2X1 U65178 ( .A(n61141), .B(n61142), .Y(n61137) );
  NAND2X1 U65179 ( .A(n60935), .B(n60936), .Y(n60940) );
  NOR2X1 U65180 ( .A(n60940), .B(n60937), .Y(n60938) );
  OR2X1 U65181 ( .A(n60939), .B(n60940), .Y(n60941) );
  NAND2X1 U65182 ( .A(n40393), .B(n43496), .Y(n61161) );
  NOR2X1 U65183 ( .A(n43469), .B(n60942), .Y(n60943) );
  XNOR2X1 U65184 ( .A(n61161), .B(n60943), .Y(n60944) );
  XNOR2X1 U65185 ( .A(n36720), .B(n60944), .Y(n60968) );
  NAND2X1 U65186 ( .A(n39650), .B(n39604), .Y(n60945) );
  NOR2X1 U65187 ( .A(n46366), .B(n40019), .Y(n60947) );
  NAND2X1 U65188 ( .A(n42383), .B(n42227), .Y(n60946) );
  NAND2X1 U65189 ( .A(n60950), .B(n38831), .Y(n60954) );
  NAND2X1 U65190 ( .A(n60952), .B(n60951), .Y(n60953) );
  NOR2X1 U65191 ( .A(n60954), .B(n60953), .Y(n60955) );
  NOR2X1 U65192 ( .A(n39192), .B(n60955), .Y(n60957) );
  NAND2X1 U65193 ( .A(n60957), .B(n60956), .Y(n61196) );
  NAND2X1 U65194 ( .A(n61169), .B(n61196), .Y(n61171) );
  NAND2X1 U65195 ( .A(n44069), .B(n61193), .Y(n60965) );
  NOR2X1 U65196 ( .A(n60959), .B(n60953), .Y(n60963) );
  NOR2X1 U65197 ( .A(n60961), .B(n60960), .Y(n60962) );
  OR2X1 U65198 ( .A(n60963), .B(n60962), .Y(n60964) );
  NOR2X1 U65199 ( .A(n60965), .B(n60964), .Y(n60966) );
  XNOR2X1 U65200 ( .A(n61171), .B(n60967), .Y(n61162) );
  INVX1 U65201 ( .A(n61162), .Y(n61165) );
  XNOR2X1 U65202 ( .A(n60968), .B(n61165), .Y(n61136) );
  NAND2X1 U65203 ( .A(n39940), .B(n43487), .Y(n61139) );
  NAND2X1 U65204 ( .A(n60970), .B(n60969), .Y(n60971) );
  NAND2X1 U65205 ( .A(n60972), .B(n60971), .Y(n61150) );
  XNOR2X1 U65206 ( .A(n61135), .B(n61139), .Y(n60973) );
  NOR2X1 U65207 ( .A(n61203), .B(n40496), .Y(n60977) );
  NAND2X1 U65208 ( .A(n43841), .B(n43484), .Y(n62423) );
  NAND2X1 U65209 ( .A(n39061), .B(n62423), .Y(n60976) );
  NOR2X1 U65210 ( .A(n60977), .B(n60976), .Y(n60981) );
  OR2X1 U65211 ( .A(n62423), .B(n39061), .Y(n60979) );
  NAND2X1 U65212 ( .A(n60979), .B(n60978), .Y(n60980) );
  INVX1 U65213 ( .A(n61216), .Y(n61218) );
  XNOR2X1 U65214 ( .A(n61217), .B(n61218), .Y(n60990) );
  NOR2X1 U65215 ( .A(n38516), .B(n60985), .Y(n60984) );
  NOR2X1 U65216 ( .A(n60982), .B(n38517), .Y(n60983) );
  NOR2X1 U65217 ( .A(n60983), .B(n60984), .Y(n60989) );
  INVX1 U65218 ( .A(n60985), .Y(n60987) );
  NAND2X1 U65219 ( .A(n60987), .B(n60986), .Y(n60988) );
  XNOR2X1 U65220 ( .A(n60990), .B(n40595), .Y(n61132) );
  INVX1 U65221 ( .A(n61132), .Y(n61129) );
  XNOR2X1 U65222 ( .A(n61131), .B(n61129), .Y(n61001) );
  NOR2X1 U65223 ( .A(n41278), .B(n60997), .Y(n60996) );
  NOR2X1 U65224 ( .A(n41278), .B(n60998), .Y(n60995) );
  NOR2X1 U65225 ( .A(n60996), .B(n60995), .Y(n61000) );
  OR2X1 U65226 ( .A(n60998), .B(n60997), .Y(n60999) );
  NAND2X1 U65227 ( .A(n60999), .B(n61000), .Y(n61130) );
  XNOR2X1 U65228 ( .A(n61001), .B(n38693), .Y(n61220) );
  INVX1 U65229 ( .A(n61220), .Y(n61222) );
  XNOR2X1 U65230 ( .A(n61221), .B(n61222), .Y(n61025) );
  NOR2X1 U65231 ( .A(n61002), .B(n61003), .Y(n61005) );
  NOR2X1 U65232 ( .A(n61003), .B(n61006), .Y(n61004) );
  NOR2X1 U65233 ( .A(n61005), .B(n61004), .Y(n61024) );
  INVX1 U65234 ( .A(n61006), .Y(n61022) );
  XNOR2X1 U65235 ( .A(n60586), .B(n61014), .Y(n61015) );
  NAND2X1 U65236 ( .A(n61016), .B(n61015), .Y(n61017) );
  NAND2X1 U65237 ( .A(n61018), .B(n61017), .Y(n61020) );
  NAND2X1 U65238 ( .A(n61020), .B(n61019), .Y(n61021) );
  NAND2X1 U65239 ( .A(n61022), .B(n61021), .Y(n61023) );
  NAND2X1 U65240 ( .A(n61024), .B(n61023), .Y(n61219) );
  NOR2X1 U65241 ( .A(n40945), .B(n61028), .Y(n61031) );
  NOR2X1 U65242 ( .A(n40945), .B(n61029), .Y(n61030) );
  NAND2X1 U65243 ( .A(n61035), .B(n61034), .Y(n61041) );
  INVX1 U65244 ( .A(n61036), .Y(n61039) );
  NAND2X1 U65245 ( .A(n39863), .B(n61037), .Y(n61038) );
  NAND2X1 U65246 ( .A(n61039), .B(n61038), .Y(n61040) );
  NAND2X1 U65247 ( .A(n61041), .B(n61040), .Y(n61126) );
  INVX1 U65248 ( .A(n61235), .Y(n61233) );
  INVX1 U65249 ( .A(n61044), .Y(n61047) );
  NAND2X1 U65250 ( .A(n39219), .B(n61045), .Y(n61046) );
  INVX1 U65251 ( .A(n61120), .Y(n61122) );
  XNOR2X1 U65252 ( .A(n61121), .B(n61122), .Y(n61059) );
  NAND2X1 U65253 ( .A(n61049), .B(n61048), .Y(n61050) );
  INVX1 U65254 ( .A(n61050), .Y(n61051) );
  NOR2X1 U65255 ( .A(n61052), .B(n61051), .Y(n61053) );
  NOR2X1 U65256 ( .A(n61054), .B(n61053), .Y(n61058) );
  NAND2X1 U65257 ( .A(n42823), .B(n61056), .Y(n61057) );
  NAND2X1 U65258 ( .A(n61058), .B(n61057), .Y(n61119) );
  INVX1 U65259 ( .A(n61119), .Y(n61123) );
  XNOR2X1 U65260 ( .A(n61059), .B(n61123), .Y(n62384) );
  XNOR2X1 U65261 ( .A(n61240), .B(n36455), .Y(n61068) );
  NOR2X1 U65262 ( .A(n61063), .B(n61060), .Y(n61065) );
  NAND2X1 U65263 ( .A(n61062), .B(n61061), .Y(n61066) );
  XNOR2X1 U65264 ( .A(n61068), .B(n39215), .Y(n61263) );
  INVX1 U65265 ( .A(n61263), .Y(n61247) );
  XNOR2X1 U65266 ( .A(n61069), .B(n61247), .Y(n61070) );
  XNOR2X1 U65267 ( .A(n36743), .B(n61070), .Y(n61273) );
  INVX1 U65268 ( .A(n61273), .Y(n61071) );
  NAND2X1 U65269 ( .A(n61073), .B(n61072), .Y(n61268) );
  NAND2X1 U65270 ( .A(n61268), .B(n61269), .Y(n61272) );
  INVX1 U65271 ( .A(n61286), .Y(n61284) );
  XNOR2X1 U65272 ( .A(n61076), .B(n61284), .Y(n61296) );
  INVX1 U65273 ( .A(n61296), .Y(n61291) );
  XNOR2X1 U65274 ( .A(n61295), .B(n61291), .Y(n61077) );
  INVX1 U65275 ( .A(n61100), .Y(n61102) );
  XNOR2X1 U65276 ( .A(n61079), .B(n61102), .Y(n61098) );
  INVX1 U65277 ( .A(n61098), .Y(n61097) );
  XNOR2X1 U65278 ( .A(n62356), .B(n61097), .Y(n61091) );
  NAND2X1 U65279 ( .A(n61084), .B(n61080), .Y(n61090) );
  INVX1 U65280 ( .A(n61081), .Y(n61088) );
  INVX1 U65281 ( .A(n61082), .Y(n61083) );
  NOR2X1 U65282 ( .A(n61084), .B(n61083), .Y(n61086) );
  NAND2X1 U65283 ( .A(n61086), .B(n61085), .Y(n61087) );
  NAND2X1 U65284 ( .A(n61088), .B(n61087), .Y(n61089) );
  XNOR2X1 U65285 ( .A(n61091), .B(n39505), .Y(n61094) );
  XNOR2X1 U65286 ( .A(n61094), .B(n42025), .Y(n61092) );
  INVX1 U65287 ( .A(n61094), .Y(n61095) );
  NAND2X1 U65288 ( .A(n39873), .B(n61095), .Y(n61096) );
  NAND2X1 U65289 ( .A(n43735), .B(n43985), .Y(n62343) );
  INVX1 U65290 ( .A(n62356), .Y(n61099) );
  NAND2X1 U65291 ( .A(n39505), .B(n61098), .Y(n62357) );
  NAND2X1 U65292 ( .A(n61100), .B(n36607), .Y(n63033) );
  NAND2X1 U65293 ( .A(n43810), .B(n43935), .Y(n62367) );
  INVX1 U65294 ( .A(n61103), .Y(n61294) );
  XNOR2X1 U65295 ( .A(n61296), .B(n61294), .Y(n61104) );
  NOR2X1 U65296 ( .A(n61116), .B(n61109), .Y(n61115) );
  NOR2X1 U65297 ( .A(n61105), .B(n61109), .Y(n61107) );
  NAND2X1 U65298 ( .A(n61107), .B(n61106), .Y(n61113) );
  NOR2X1 U65299 ( .A(n36443), .B(n61109), .Y(n61111) );
  NAND2X1 U65300 ( .A(n61111), .B(n61110), .Y(n61112) );
  NAND2X1 U65301 ( .A(n61113), .B(n61112), .Y(n61114) );
  INVX1 U65302 ( .A(n61116), .Y(n61118) );
  XNOR2X1 U65303 ( .A(n62367), .B(n39393), .Y(n61297) );
  NAND2X1 U65304 ( .A(n43926), .B(n40467), .Y(n62537) );
  NAND2X1 U65305 ( .A(n43919), .B(n40470), .Y(n62527) );
  NAND2X1 U65306 ( .A(n43890), .B(n42638), .Y(n62383) );
  INVX1 U65307 ( .A(n61121), .Y(n61125) );
  INVX1 U65308 ( .A(n62397), .Y(n62391) );
  NAND2X1 U65309 ( .A(n43860), .B(n43796), .Y(n62499) );
  INVX1 U65310 ( .A(n61131), .Y(n61134) );
  NAND2X1 U65311 ( .A(n38693), .B(n61132), .Y(n61133) );
  NAND2X1 U65312 ( .A(n43851), .B(n43776), .Y(n62492) );
  NAND2X1 U65313 ( .A(n44036), .B(n43479), .Y(n62488) );
  INVX1 U65314 ( .A(n61140), .Y(n61138) );
  NAND2X1 U65315 ( .A(n61138), .B(n61137), .Y(n61146) );
  INVX1 U65316 ( .A(n61139), .Y(n61144) );
  NAND2X1 U65317 ( .A(n61144), .B(n61143), .Y(n61145) );
  NAND2X1 U65318 ( .A(n61146), .B(n61145), .Y(n62480) );
  NAND2X1 U65319 ( .A(n43841), .B(n43486), .Y(n62479) );
  NOR2X1 U65320 ( .A(n61148), .B(n61147), .Y(n61151) );
  NOR2X1 U65321 ( .A(n36663), .B(n36664), .Y(n61152) );
  NAND2X1 U65322 ( .A(n43492), .B(n43466), .Y(n61156) );
  NOR2X1 U65323 ( .A(n61152), .B(n61156), .Y(n61155) );
  INVX1 U65324 ( .A(n61161), .Y(n61166) );
  XNOR2X1 U65325 ( .A(n61162), .B(n61166), .Y(n61153) );
  XNOR2X1 U65326 ( .A(n38233), .B(n61153), .Y(n61157) );
  NOR2X1 U65327 ( .A(n61155), .B(n61154), .Y(n61160) );
  INVX1 U65328 ( .A(n61156), .Y(n61158) );
  NAND2X1 U65329 ( .A(n61158), .B(n61157), .Y(n61159) );
  NOR2X1 U65330 ( .A(n61161), .B(n38233), .Y(n61164) );
  NOR2X1 U65331 ( .A(n61162), .B(n38233), .Y(n61163) );
  NOR2X1 U65332 ( .A(n61164), .B(n61163), .Y(n61168) );
  NAND2X1 U65333 ( .A(n61166), .B(n61165), .Y(n61167) );
  NAND2X1 U65334 ( .A(n61168), .B(n61167), .Y(n62474) );
  NOR2X1 U65335 ( .A(n43503), .B(n43459), .Y(n61170) );
  INVX1 U65336 ( .A(n61171), .Y(n61172) );
  NAND2X1 U65337 ( .A(n43471), .B(n43502), .Y(n62440) );
  INVX1 U65338 ( .A(n62905), .Y(n61175) );
  NAND2X1 U65339 ( .A(opcode_instr_w_48), .B(n61174), .Y(n64087) );
  NOR2X1 U65340 ( .A(n61175), .B(n64087), .Y(n61176) );
  NAND2X1 U65341 ( .A(n42392), .B(n61177), .Y(n61180) );
  NAND2X1 U65342 ( .A(n42392), .B(n61178), .Y(n61179) );
  OR2X1 U65343 ( .A(n43453), .B(n64087), .Y(n61181) );
  NOR2X1 U65344 ( .A(n61182), .B(n61181), .Y(n61184) );
  NOR2X1 U65345 ( .A(n64087), .B(n62902), .Y(n61183) );
  NOR2X1 U65346 ( .A(n61184), .B(n61183), .Y(n61186) );
  NAND2X1 U65347 ( .A(n42234), .B(n61186), .Y(n63830) );
  NAND2X1 U65348 ( .A(n63830), .B(n40383), .Y(n63555) );
  NAND2X1 U65349 ( .A(n42383), .B(n42227), .Y(n62443) );
  NOR2X1 U65350 ( .A(n42225), .B(n62443), .Y(n61191) );
  NAND2X1 U65351 ( .A(n40383), .B(n61192), .Y(n61194) );
  NAND2X1 U65352 ( .A(n61195), .B(n61194), .Y(n62465) );
  NAND2X1 U65353 ( .A(n63555), .B(n62465), .Y(n61199) );
  NAND2X1 U65354 ( .A(n39868), .B(n38527), .Y(n61197) );
  XNOR2X1 U65355 ( .A(n61197), .B(n39641), .Y(n61198) );
  XNOR2X1 U65356 ( .A(n61199), .B(n61198), .Y(n62442) );
  XOR2X1 U65357 ( .A(n62440), .B(n62442), .Y(n61200) );
  XNOR2X1 U65358 ( .A(n62439), .B(n61200), .Y(n62473) );
  NAND2X1 U65359 ( .A(n43464), .B(n43497), .Y(n62469) );
  XNOR2X1 U65360 ( .A(n62473), .B(n62469), .Y(n61201) );
  XNOR2X1 U65361 ( .A(n62474), .B(n61201), .Y(n62433) );
  NAND2X1 U65362 ( .A(n43493), .B(n39939), .Y(n62432) );
  XNOR2X1 U65363 ( .A(n62433), .B(n62432), .Y(n61202) );
  NAND2X1 U65364 ( .A(n61204), .B(n39061), .Y(n61206) );
  INVX1 U65365 ( .A(n61205), .Y(n62424) );
  NAND2X1 U65366 ( .A(n39899), .B(n62424), .Y(n61209) );
  NOR2X1 U65367 ( .A(n62423), .B(n41388), .Y(n61208) );
  NAND2X1 U65368 ( .A(n61206), .B(n61205), .Y(n62425) );
  NAND2X1 U65369 ( .A(n38384), .B(n38312), .Y(n62427) );
  NAND2X1 U65370 ( .A(n62425), .B(n62427), .Y(n61207) );
  NOR2X1 U65371 ( .A(n61208), .B(n61207), .Y(n61214) );
  OR2X1 U65372 ( .A(n62427), .B(n62425), .Y(n61212) );
  NOR2X1 U65373 ( .A(n62423), .B(n62427), .Y(n61210) );
  NAND2X1 U65374 ( .A(n61210), .B(n61209), .Y(n61211) );
  NAND2X1 U65375 ( .A(n61212), .B(n61211), .Y(n61213) );
  INVX1 U65376 ( .A(n62500), .Y(n62503) );
  XNOR2X1 U65377 ( .A(n62499), .B(n62503), .Y(n61225) );
  INVX1 U65378 ( .A(n61221), .Y(n61224) );
  XNOR2X1 U65379 ( .A(n61225), .B(n40082), .Y(n62420) );
  NAND2X1 U65380 ( .A(n43798), .B(n43872), .Y(n63009) );
  INVX1 U65381 ( .A(n63009), .Y(n62405) );
  NAND2X1 U65382 ( .A(n43963), .B(n42714), .Y(n62416) );
  INVX1 U65383 ( .A(n62416), .Y(n62409) );
  XNOR2X1 U65384 ( .A(n62405), .B(n41253), .Y(n61230) );
  INVX1 U65385 ( .A(n61226), .Y(n61229) );
  NAND2X1 U65386 ( .A(n39859), .B(n61227), .Y(n61228) );
  XNOR2X1 U65387 ( .A(n61230), .B(n38638), .Y(n61231) );
  XNOR2X1 U65388 ( .A(n62420), .B(n61231), .Y(n61232) );
  XNOR2X1 U65389 ( .A(n37388), .B(n61232), .Y(n62392) );
  INVX1 U65390 ( .A(n61234), .Y(n61237) );
  NAND2X1 U65391 ( .A(n38684), .B(n61235), .Y(n61236) );
  NAND2X1 U65392 ( .A(n40260), .B(n43881), .Y(n62393) );
  XNOR2X1 U65393 ( .A(n62392), .B(n61238), .Y(n61239) );
  XNOR2X1 U65394 ( .A(n62391), .B(n61239), .Y(n62380) );
  INVX1 U65395 ( .A(n62380), .Y(n62382) );
  XNOR2X1 U65396 ( .A(n62383), .B(n62382), .Y(n61246) );
  NOR2X1 U65397 ( .A(n62384), .B(n61240), .Y(n61244) );
  NAND2X1 U65398 ( .A(n61241), .B(n36455), .Y(n62387) );
  INVX1 U65399 ( .A(n61240), .Y(n62386) );
  NAND2X1 U65400 ( .A(n62386), .B(n61241), .Y(n61242) );
  NAND2X1 U65401 ( .A(n62387), .B(n61242), .Y(n61243) );
  NOR2X1 U65402 ( .A(n61244), .B(n61243), .Y(n61245) );
  XNOR2X1 U65403 ( .A(n61246), .B(n61245), .Y(n62514) );
  NOR2X1 U65404 ( .A(n42841), .B(n61255), .Y(n61249) );
  INVX1 U65405 ( .A(n61255), .Y(n61250) );
  NAND2X1 U65406 ( .A(n61254), .B(n61255), .Y(n61253) );
  INVX1 U65407 ( .A(n61251), .Y(n61252) );
  NOR2X1 U65408 ( .A(n61253), .B(n61252), .Y(n61262) );
  OR2X1 U65409 ( .A(n61255), .B(n61254), .Y(n61260) );
  NOR2X1 U65410 ( .A(n61256), .B(n61255), .Y(n61258) );
  NAND2X1 U65411 ( .A(n61258), .B(n61257), .Y(n61259) );
  NAND2X1 U65412 ( .A(n61260), .B(n61259), .Y(n61261) );
  INVX1 U65413 ( .A(n61267), .Y(n61264) );
  NAND2X1 U65414 ( .A(n36743), .B(n61264), .Y(n61265) );
  NAND2X1 U65415 ( .A(n43788), .B(n43905), .Y(n62376) );
  INVX1 U65416 ( .A(n61275), .Y(n61271) );
  NAND2X1 U65417 ( .A(n61269), .B(n61268), .Y(n61270) );
  OR2X1 U65418 ( .A(n61273), .B(n61270), .Y(n61276) );
  NAND2X1 U65419 ( .A(n61271), .B(n61276), .Y(n62519) );
  NAND2X1 U65420 ( .A(n61273), .B(n61272), .Y(n62520) );
  NAND2X1 U65421 ( .A(n43910), .B(n40482), .Y(n62522) );
  NOR2X1 U65422 ( .A(n39429), .B(n61274), .Y(n61281) );
  NOR2X1 U65423 ( .A(n61275), .B(n62522), .Y(n61277) );
  NAND2X1 U65424 ( .A(n61277), .B(n61276), .Y(n61278) );
  NAND2X1 U65425 ( .A(n61279), .B(n61278), .Y(n61280) );
  NOR2X1 U65426 ( .A(n61281), .B(n61280), .Y(n61282) );
  XNOR2X1 U65427 ( .A(n61282), .B(n62850), .Y(n62528) );
  INVX1 U65428 ( .A(n62528), .Y(n62526) );
  INVX1 U65429 ( .A(n61285), .Y(n61288) );
  NAND2X1 U65430 ( .A(n38885), .B(n61286), .Y(n61287) );
  INVX1 U65431 ( .A(n62538), .Y(n62534) );
  INVX1 U65432 ( .A(n62368), .Y(n62372) );
  XNOR2X1 U65433 ( .A(n61297), .B(n62372), .Y(n63034) );
  NAND2X1 U65434 ( .A(n43821), .B(n43944), .Y(n63032) );
  XNOR2X1 U65435 ( .A(n62363), .B(n62364), .Y(n61298) );
  NAND2X1 U65436 ( .A(n43758), .B(n43974), .Y(n62355) );
  INVX1 U65437 ( .A(n62355), .Y(n62345) );
  XNOR2X1 U65438 ( .A(n61298), .B(n62345), .Y(n62342) );
  XNOR2X1 U65439 ( .A(n62559), .B(n42052), .Y(n61299) );
  XNOR2X1 U65440 ( .A(n39666), .B(n61299), .Y(n62340) );
  XNOR2X1 U65441 ( .A(n61300), .B(n42039), .Y(n61301) );
  XNOR2X1 U65442 ( .A(n37394), .B(n61301), .Y(n61440) );
  XNOR2X1 U65443 ( .A(n61302), .B(n42016), .Y(n61303) );
  XNOR2X1 U65444 ( .A(n39999), .B(n61303), .Y(n61443) );
  INVX1 U65445 ( .A(n61443), .Y(n61428) );
  XNOR2X1 U65446 ( .A(n61304), .B(n42007), .Y(n61305) );
  XNOR2X1 U65447 ( .A(n40549), .B(n61305), .Y(n61445) );
  XNOR2X1 U65448 ( .A(n61306), .B(n41993), .Y(n61307) );
  XNOR2X1 U65449 ( .A(n61308), .B(n41982), .Y(n61309) );
  XNOR2X1 U65450 ( .A(n40357), .B(n61309), .Y(n61449) );
  INVX1 U65451 ( .A(n61449), .Y(n61422) );
  XNOR2X1 U65452 ( .A(n61310), .B(n41972), .Y(n61311) );
  XNOR2X1 U65453 ( .A(n61312), .B(n61311), .Y(n61451) );
  XNOR2X1 U65454 ( .A(n61313), .B(n41962), .Y(n61314) );
  XNOR2X1 U65455 ( .A(n61315), .B(n61314), .Y(n61453) );
  INVX1 U65456 ( .A(n61453), .Y(n61417) );
  XNOR2X1 U65457 ( .A(n61316), .B(n41953), .Y(n61317) );
  XNOR2X1 U65458 ( .A(n36461), .B(n61317), .Y(n61455) );
  XNOR2X1 U65459 ( .A(n61318), .B(n38150), .Y(n61319) );
  XNOR2X1 U65460 ( .A(n41943), .B(n61319), .Y(n61457) );
  INVX1 U65461 ( .A(n61457), .Y(n61412) );
  XNOR2X1 U65462 ( .A(n61320), .B(n38149), .Y(n61321) );
  XNOR2X1 U65463 ( .A(n41932), .B(n61321), .Y(n61459) );
  XNOR2X1 U65464 ( .A(n61322), .B(n41921), .Y(n61323) );
  XNOR2X1 U65465 ( .A(n40632), .B(n61323), .Y(n61461) );
  INVX1 U65466 ( .A(n61461), .Y(n61405) );
  XNOR2X1 U65467 ( .A(n61324), .B(n41913), .Y(n61325) );
  XNOR2X1 U65468 ( .A(n61326), .B(n61325), .Y(n61463) );
  INVX1 U65469 ( .A(n61463), .Y(n61401) );
  XNOR2X1 U65470 ( .A(n61327), .B(n39098), .Y(n61328) );
  XNOR2X1 U65471 ( .A(n41902), .B(n61328), .Y(n61466) );
  XNOR2X1 U65472 ( .A(n61329), .B(n40243), .Y(n61330) );
  XNOR2X1 U65473 ( .A(n41890), .B(n61330), .Y(n61468) );
  INVX1 U65474 ( .A(n61468), .Y(n61394) );
  XNOR2X1 U65475 ( .A(n61331), .B(n39149), .Y(n61332) );
  XNOR2X1 U65476 ( .A(n41881), .B(n61332), .Y(n61470) );
  XNOR2X1 U65477 ( .A(n61333), .B(n39675), .Y(n61334) );
  XNOR2X1 U65478 ( .A(n41870), .B(n61334), .Y(n61473) );
  INVX1 U65479 ( .A(n61473), .Y(n61389) );
  XNOR2X1 U65480 ( .A(n61335), .B(n41857), .Y(n61336) );
  XNOR2X1 U65481 ( .A(n61337), .B(n61336), .Y(n61476) );
  XNOR2X1 U65482 ( .A(n61339), .B(n61338), .Y(n61340) );
  XNOR2X1 U65483 ( .A(n41844), .B(n61340), .Y(n61479) );
  INVX1 U65484 ( .A(n61479), .Y(n61380) );
  XNOR2X1 U65485 ( .A(n61341), .B(n38915), .Y(n61342) );
  XNOR2X1 U65486 ( .A(n41831), .B(n61342), .Y(n61482) );
  XNOR2X1 U65487 ( .A(n61344), .B(n61343), .Y(n61345) );
  XNOR2X1 U65488 ( .A(n41816), .B(n61345), .Y(n61486) );
  INVX1 U65489 ( .A(n61486), .Y(n61369) );
  XNOR2X1 U65490 ( .A(n61347), .B(n61346), .Y(n61348) );
  XNOR2X1 U65491 ( .A(n41799), .B(n61348), .Y(n61489) );
  XNOR2X1 U65492 ( .A(n61350), .B(n61349), .Y(n61351) );
  XNOR2X1 U65493 ( .A(n41781), .B(n61351), .Y(n61492) );
  INVX1 U65494 ( .A(n61492), .Y(n61359) );
  NAND2X1 U65495 ( .A(n42715), .B(n72810), .Y(n61497) );
  NAND2X1 U65496 ( .A(n44070), .B(n43780), .Y(n61498) );
  INVX1 U65497 ( .A(n61499), .Y(n61494) );
  NAND2X1 U65498 ( .A(n61353), .B(n61352), .Y(n61355) );
  NAND2X1 U65499 ( .A(n61355), .B(n61354), .Y(n61495) );
  NAND2X1 U65500 ( .A(n61494), .B(n40354), .Y(n61358) );
  NAND2X1 U65501 ( .A(n61499), .B(n61495), .Y(n61356) );
  NAND2X1 U65502 ( .A(n41790), .B(n61356), .Y(n61357) );
  NAND2X1 U65503 ( .A(n61358), .B(n61357), .Y(n61360) );
  NAND2X1 U65504 ( .A(n61359), .B(n61360), .Y(n61363) );
  INVX1 U65505 ( .A(n61360), .Y(n61491) );
  NAND2X1 U65506 ( .A(n61491), .B(n61492), .Y(n61361) );
  NAND2X1 U65507 ( .A(n41806), .B(n61361), .Y(n61362) );
  NAND2X1 U65508 ( .A(n61363), .B(n61362), .Y(n61364) );
  NAND2X1 U65509 ( .A(n61489), .B(n61364), .Y(n61368) );
  INVX1 U65510 ( .A(n61364), .Y(n61488) );
  INVX1 U65511 ( .A(n61489), .Y(n61365) );
  NAND2X1 U65512 ( .A(n61488), .B(n61365), .Y(n61366) );
  NAND2X1 U65513 ( .A(n41818), .B(n61366), .Y(n61367) );
  NAND2X1 U65514 ( .A(n61368), .B(n61367), .Y(n61370) );
  NAND2X1 U65515 ( .A(n61369), .B(n61370), .Y(n61373) );
  INVX1 U65516 ( .A(n61370), .Y(n61485) );
  NAND2X1 U65517 ( .A(n61485), .B(n61486), .Y(n61371) );
  NAND2X1 U65518 ( .A(n41834), .B(n61371), .Y(n61372) );
  NAND2X1 U65519 ( .A(n61373), .B(n61372), .Y(n61375) );
  NAND2X1 U65520 ( .A(n61482), .B(n61375), .Y(n61379) );
  INVX1 U65521 ( .A(n61374), .Y(n61481) );
  INVX1 U65522 ( .A(n61375), .Y(n61484) );
  INVX1 U65523 ( .A(n61482), .Y(n61376) );
  NAND2X1 U65524 ( .A(n61484), .B(n61376), .Y(n61377) );
  NAND2X1 U65525 ( .A(n61481), .B(n61377), .Y(n61378) );
  NAND2X1 U65526 ( .A(n61379), .B(n61378), .Y(n61381) );
  NAND2X1 U65527 ( .A(n61380), .B(n61381), .Y(n61384) );
  INVX1 U65528 ( .A(n61381), .Y(n61478) );
  NAND2X1 U65529 ( .A(n61478), .B(n61479), .Y(n61382) );
  NAND2X1 U65530 ( .A(n41863), .B(n61382), .Y(n61383) );
  NAND2X1 U65531 ( .A(n61384), .B(n61383), .Y(n61385) );
  NAND2X1 U65532 ( .A(n61476), .B(n61385), .Y(n61388) );
  INVX1 U65533 ( .A(n61385), .Y(n61475) );
  NAND2X1 U65534 ( .A(n41873), .B(n61386), .Y(n61387) );
  NAND2X1 U65535 ( .A(n61388), .B(n61387), .Y(n61390) );
  INVX1 U65536 ( .A(n61390), .Y(n61472) );
  NAND2X1 U65537 ( .A(n61472), .B(n61473), .Y(n61391) );
  INVX1 U65538 ( .A(n61470), .Y(n61392) );
  NAND2X1 U65539 ( .A(n39547), .B(n61392), .Y(n61393) );
  NAND2X1 U65540 ( .A(n61394), .B(n39184), .Y(n61397) );
  NAND2X1 U65541 ( .A(n39463), .B(n61468), .Y(n61395) );
  NAND2X1 U65542 ( .A(n41905), .B(n61395), .Y(n61396) );
  NAND2X1 U65543 ( .A(n61397), .B(n61396), .Y(n61398) );
  INVX1 U65544 ( .A(n61398), .Y(n61465) );
  INVX1 U65545 ( .A(n61466), .Y(n61399) );
  NAND2X1 U65546 ( .A(n61465), .B(n61399), .Y(n61400) );
  NAND2X1 U65547 ( .A(n61401), .B(n38146), .Y(n61404) );
  NAND2X1 U65548 ( .A(n39375), .B(n61463), .Y(n61402) );
  NAND2X1 U65549 ( .A(n41926), .B(n61402), .Y(n61403) );
  NAND2X1 U65550 ( .A(n61404), .B(n61403), .Y(n61406) );
  NAND2X1 U65551 ( .A(n36346), .B(n61461), .Y(n61407) );
  NAND2X1 U65552 ( .A(n61459), .B(n39634), .Y(n61411) );
  INVX1 U65553 ( .A(n61459), .Y(n61408) );
  NAND2X1 U65554 ( .A(n39813), .B(n61408), .Y(n61409) );
  NAND2X1 U65555 ( .A(n41948), .B(n61409), .Y(n61410) );
  NAND2X1 U65556 ( .A(n61411), .B(n61410), .Y(n61413) );
  NAND2X1 U65557 ( .A(n36394), .B(n61457), .Y(n61414) );
  NAND2X1 U65558 ( .A(n38746), .B(n61453), .Y(n61419) );
  INVX1 U65559 ( .A(n61451), .Y(n61420) );
  NAND2X1 U65560 ( .A(n40608), .B(n61420), .Y(n61421) );
  NAND2X1 U65561 ( .A(n61447), .B(n36456), .Y(n61425) );
  NAND2X1 U65562 ( .A(n61425), .B(n61424), .Y(n61426) );
  INVX1 U65563 ( .A(n61445), .Y(n61427) );
  NAND2X1 U65564 ( .A(n36579), .B(n61443), .Y(n61430) );
  XNOR2X1 U65565 ( .A(n61431), .B(n42027), .Y(n61432) );
  XNOR2X1 U65566 ( .A(n37891), .B(n61432), .Y(n61441) );
  INVX1 U65567 ( .A(n61441), .Y(n61433) );
  NAND2X1 U65568 ( .A(n61433), .B(n39482), .Y(n61435) );
  NAND2X1 U65569 ( .A(n61434), .B(n61435), .Y(n61439) );
  NAND2X1 U65570 ( .A(n61435), .B(n61434), .Y(n61436) );
  OR2X1 U65571 ( .A(n61440), .B(n61436), .Y(n61437) );
  XNOR2X1 U65572 ( .A(n62340), .B(n38925), .Y(n61438) );
  XNOR2X1 U65573 ( .A(n42064), .B(n61438), .Y(n62338) );
  INVX1 U65574 ( .A(n61589), .Y(n61584) );
  XNOR2X1 U65575 ( .A(n61441), .B(n40073), .Y(n61442) );
  XNOR2X1 U65576 ( .A(n42043), .B(n61442), .Y(n61591) );
  XNOR2X1 U65577 ( .A(n61443), .B(n36579), .Y(n61444) );
  XNOR2X1 U65578 ( .A(n42031), .B(n61444), .Y(n61594) );
  XNOR2X1 U65579 ( .A(n61445), .B(n37925), .Y(n61446) );
  XNOR2X1 U65580 ( .A(n42019), .B(n61446), .Y(n61596) );
  INVX1 U65581 ( .A(n61596), .Y(n61574) );
  XNOR2X1 U65582 ( .A(n37947), .B(n61447), .Y(n61448) );
  XNOR2X1 U65583 ( .A(n42010), .B(n61448), .Y(n61598) );
  INVX1 U65584 ( .A(n61598), .Y(n61572) );
  XNOR2X1 U65585 ( .A(n61449), .B(n40230), .Y(n61450) );
  XNOR2X1 U65586 ( .A(n41997), .B(n61450), .Y(n61601) );
  XNOR2X1 U65587 ( .A(n61451), .B(n40608), .Y(n61452) );
  XNOR2X1 U65588 ( .A(n41986), .B(n61452), .Y(n61603) );
  INVX1 U65589 ( .A(n61603), .Y(n61565) );
  XNOR2X1 U65590 ( .A(n61453), .B(n38746), .Y(n61454) );
  XNOR2X1 U65591 ( .A(n41976), .B(n61454), .Y(n61605) );
  XNOR2X1 U65592 ( .A(n61455), .B(n40011), .Y(n61456) );
  XNOR2X1 U65593 ( .A(n41965), .B(n61456), .Y(n61607) );
  XNOR2X1 U65594 ( .A(n61457), .B(n36394), .Y(n61458) );
  XNOR2X1 U65595 ( .A(n41956), .B(n61458), .Y(n61609) );
  XNOR2X1 U65596 ( .A(n61459), .B(n39813), .Y(n61460) );
  XNOR2X1 U65597 ( .A(n41948), .B(n61460), .Y(n61611) );
  INVX1 U65598 ( .A(n61611), .Y(n61554) );
  XNOR2X1 U65599 ( .A(n61461), .B(n36346), .Y(n61462) );
  XNOR2X1 U65600 ( .A(n41936), .B(n61462), .Y(n61614) );
  XNOR2X1 U65601 ( .A(n61463), .B(n39375), .Y(n61464) );
  XNOR2X1 U65602 ( .A(n41926), .B(n61464), .Y(n61616) );
  XNOR2X1 U65603 ( .A(n61466), .B(n61465), .Y(n61467) );
  XNOR2X1 U65604 ( .A(n41916), .B(n61467), .Y(n61618) );
  INVX1 U65605 ( .A(n61618), .Y(n61545) );
  XNOR2X1 U65606 ( .A(n39463), .B(n61468), .Y(n61469) );
  XNOR2X1 U65607 ( .A(n41905), .B(n61469), .Y(n61621) );
  XNOR2X1 U65608 ( .A(n61470), .B(n39547), .Y(n61471) );
  XNOR2X1 U65609 ( .A(n41893), .B(n61471), .Y(n61623) );
  INVX1 U65610 ( .A(n61623), .Y(n61538) );
  XNOR2X1 U65611 ( .A(n61473), .B(n61472), .Y(n61474) );
  XNOR2X1 U65612 ( .A(n41884), .B(n61474), .Y(n61625) );
  XNOR2X1 U65613 ( .A(n61476), .B(n61475), .Y(n61477) );
  XNOR2X1 U65614 ( .A(n41873), .B(n61477), .Y(n61628) );
  INVX1 U65615 ( .A(n61628), .Y(n61530) );
  XNOR2X1 U65616 ( .A(n61479), .B(n61478), .Y(n61480) );
  XNOR2X1 U65617 ( .A(n41863), .B(n61480), .Y(n61631) );
  XNOR2X1 U65618 ( .A(n61482), .B(n61481), .Y(n61483) );
  XNOR2X1 U65619 ( .A(n61484), .B(n61483), .Y(n61634) );
  INVX1 U65620 ( .A(n61634), .Y(n61522) );
  XNOR2X1 U65621 ( .A(n61486), .B(n61485), .Y(n61487) );
  XNOR2X1 U65622 ( .A(n41834), .B(n61487), .Y(n61636) );
  XNOR2X1 U65623 ( .A(n61489), .B(n61488), .Y(n61490) );
  XNOR2X1 U65624 ( .A(n41818), .B(n61490), .Y(n61638) );
  INVX1 U65625 ( .A(n61638), .Y(n61514) );
  XNOR2X1 U65626 ( .A(n61492), .B(n61491), .Y(n61493) );
  XNOR2X1 U65627 ( .A(n41806), .B(n61493), .Y(n61642) );
  XNOR2X1 U65628 ( .A(n61495), .B(n61494), .Y(n61496) );
  XNOR2X1 U65629 ( .A(n41790), .B(n61496), .Y(n61644) );
  INVX1 U65630 ( .A(n61644), .Y(n61504) );
  NAND2X1 U65631 ( .A(n42715), .B(n43743), .Y(n61649) );
  NAND2X1 U65632 ( .A(n73384), .B(n72810), .Y(n61650) );
  INVX1 U65633 ( .A(n61651), .Y(n61646) );
  INVX1 U65634 ( .A(n61647), .Y(n61500) );
  NAND2X1 U65635 ( .A(n61646), .B(n61500), .Y(n61503) );
  NAND2X1 U65636 ( .A(n61651), .B(n61647), .Y(n61501) );
  NAND2X1 U65637 ( .A(n41789), .B(n61501), .Y(n61502) );
  NAND2X1 U65638 ( .A(n61503), .B(n61502), .Y(n61505) );
  NAND2X1 U65639 ( .A(n61504), .B(n61505), .Y(n61508) );
  NAND2X1 U65640 ( .A(n36397), .B(n61644), .Y(n61506) );
  NAND2X1 U65641 ( .A(n41810), .B(n61506), .Y(n61507) );
  NAND2X1 U65642 ( .A(n61508), .B(n61507), .Y(n61509) );
  NAND2X1 U65643 ( .A(n61642), .B(n61509), .Y(n61513) );
  INVX1 U65644 ( .A(n61509), .Y(n61641) );
  INVX1 U65645 ( .A(n61642), .Y(n61510) );
  NAND2X1 U65646 ( .A(n61641), .B(n61510), .Y(n61511) );
  NAND2X1 U65647 ( .A(n41822), .B(n61511), .Y(n61512) );
  NAND2X1 U65648 ( .A(n61513), .B(n61512), .Y(n61515) );
  INVX1 U65649 ( .A(n61515), .Y(n61640) );
  NAND2X1 U65650 ( .A(n61640), .B(n61638), .Y(n61516) );
  NAND2X1 U65651 ( .A(n61636), .B(n61517), .Y(n61521) );
  INVX1 U65652 ( .A(n61636), .Y(n61518) );
  NAND2X1 U65653 ( .A(n38761), .B(n61518), .Y(n61519) );
  NAND2X1 U65654 ( .A(n41852), .B(n61519), .Y(n61520) );
  NAND2X1 U65655 ( .A(n61521), .B(n61520), .Y(n61523) );
  NAND2X1 U65656 ( .A(n61522), .B(n61523), .Y(n61526) );
  INVX1 U65657 ( .A(n61523), .Y(n61633) );
  NAND2X1 U65658 ( .A(n61633), .B(n61634), .Y(n61524) );
  NAND2X1 U65659 ( .A(n41867), .B(n61524), .Y(n61525) );
  NAND2X1 U65660 ( .A(n61526), .B(n61525), .Y(n61527) );
  INVX1 U65661 ( .A(n61527), .Y(n61630) );
  INVX1 U65662 ( .A(n61631), .Y(n61528) );
  NAND2X1 U65663 ( .A(n61630), .B(n61528), .Y(n61529) );
  NAND2X1 U65664 ( .A(n61530), .B(n61531), .Y(n61534) );
  INVX1 U65665 ( .A(n61531), .Y(n61627) );
  NAND2X1 U65666 ( .A(n41888), .B(n61532), .Y(n61533) );
  NAND2X1 U65667 ( .A(n61534), .B(n61533), .Y(n61535) );
  INVX1 U65668 ( .A(n61625), .Y(n61536) );
  NAND2X1 U65669 ( .A(n38993), .B(n61536), .Y(n61537) );
  NAND2X1 U65670 ( .A(n61538), .B(n39183), .Y(n61541) );
  NAND2X1 U65671 ( .A(n39400), .B(n61623), .Y(n61539) );
  NAND2X1 U65672 ( .A(n41909), .B(n61539), .Y(n61540) );
  NAND2X1 U65673 ( .A(n61541), .B(n61540), .Y(n61542) );
  INVX1 U65674 ( .A(n61542), .Y(n61620) );
  INVX1 U65675 ( .A(n61621), .Y(n61543) );
  NAND2X1 U65676 ( .A(n61620), .B(n61543), .Y(n61544) );
  NAND2X1 U65677 ( .A(n61618), .B(n39642), .Y(n61546) );
  NAND2X1 U65678 ( .A(n61616), .B(n38102), .Y(n61550) );
  INVX1 U65679 ( .A(n61616), .Y(n61547) );
  NAND2X1 U65680 ( .A(n38453), .B(n61547), .Y(n61548) );
  NAND2X1 U65681 ( .A(n41941), .B(n61548), .Y(n61549) );
  NAND2X1 U65682 ( .A(n61550), .B(n61549), .Y(n61551) );
  INVX1 U65683 ( .A(n61551), .Y(n61613) );
  INVX1 U65684 ( .A(n61614), .Y(n61552) );
  NAND2X1 U65685 ( .A(n61613), .B(n61552), .Y(n61553) );
  NAND2X1 U65686 ( .A(n39830), .B(n61611), .Y(n61555) );
  INVX1 U65687 ( .A(n61609), .Y(n61557) );
  NAND2X1 U65688 ( .A(n38017), .B(n61557), .Y(n61558) );
  NAND2X1 U65689 ( .A(n61607), .B(n39847), .Y(n61562) );
  INVX1 U65690 ( .A(n61607), .Y(n61559) );
  NAND2X1 U65691 ( .A(n40030), .B(n61559), .Y(n61560) );
  NAND2X1 U65692 ( .A(n41981), .B(n61560), .Y(n61561) );
  NAND2X1 U65693 ( .A(n61562), .B(n61561), .Y(n61563) );
  NAND2X1 U65694 ( .A(n61565), .B(n40038), .Y(n61568) );
  NAND2X1 U65695 ( .A(n40108), .B(n61603), .Y(n61566) );
  NAND2X1 U65696 ( .A(n42003), .B(n61566), .Y(n61567) );
  NAND2X1 U65697 ( .A(n61568), .B(n61567), .Y(n61569) );
  INVX1 U65698 ( .A(n61569), .Y(n61600) );
  INVX1 U65699 ( .A(n61601), .Y(n61570) );
  NAND2X1 U65700 ( .A(n61600), .B(n61570), .Y(n61571) );
  NAND2X1 U65701 ( .A(n40238), .B(n61598), .Y(n61573) );
  NAND2X1 U65702 ( .A(n61574), .B(n61575), .Y(n61578) );
  NAND2X1 U65703 ( .A(n36553), .B(n61596), .Y(n61576) );
  NAND2X1 U65704 ( .A(n42038), .B(n61576), .Y(n61577) );
  NAND2X1 U65705 ( .A(n61578), .B(n61577), .Y(n61579) );
  INVX1 U65706 ( .A(n61579), .Y(n61593) );
  INVX1 U65707 ( .A(n61594), .Y(n61580) );
  NAND2X1 U65708 ( .A(n61593), .B(n61580), .Y(n61581) );
  INVX1 U65709 ( .A(n61591), .Y(n61583) );
  INVX1 U65710 ( .A(n61585), .Y(n61588) );
  XNOR2X1 U65711 ( .A(n62338), .B(n40314), .Y(n61587) );
  XNOR2X1 U65712 ( .A(n42082), .B(n61587), .Y(n62564) );
  XNOR2X1 U65713 ( .A(n61589), .B(n61588), .Y(n61590) );
  XNOR2X1 U65714 ( .A(n42074), .B(n61590), .Y(n61751) );
  XNOR2X1 U65715 ( .A(n61591), .B(n36556), .Y(n61592) );
  XNOR2X1 U65716 ( .A(n42063), .B(n61592), .Y(n61754) );
  INVX1 U65717 ( .A(n61754), .Y(n61743) );
  XNOR2X1 U65718 ( .A(n61594), .B(n61593), .Y(n61595) );
  XNOR2X1 U65719 ( .A(n42051), .B(n61595), .Y(n61757) );
  INVX1 U65720 ( .A(n61757), .Y(n61739) );
  XNOR2X1 U65721 ( .A(n61596), .B(n36553), .Y(n61597) );
  XNOR2X1 U65722 ( .A(n42038), .B(n61597), .Y(n61759) );
  XNOR2X1 U65723 ( .A(n61598), .B(n38688), .Y(n61599) );
  XNOR2X1 U65724 ( .A(n42024), .B(n61599), .Y(n61762) );
  XNOR2X1 U65725 ( .A(n61601), .B(n61600), .Y(n61602) );
  XNOR2X1 U65726 ( .A(n42014), .B(n61602), .Y(n61765) );
  INVX1 U65727 ( .A(n61765), .Y(n61730) );
  XNOR2X1 U65728 ( .A(n61603), .B(n38675), .Y(n61604) );
  XNOR2X1 U65729 ( .A(n42003), .B(n61604), .Y(n61768) );
  XNOR2X1 U65730 ( .A(n61605), .B(n36395), .Y(n61606) );
  XNOR2X1 U65731 ( .A(n41990), .B(n61606), .Y(n61771) );
  INVX1 U65732 ( .A(n61771), .Y(n61724) );
  XNOR2X1 U65733 ( .A(n61607), .B(n40030), .Y(n61608) );
  XNOR2X1 U65734 ( .A(n41981), .B(n61608), .Y(n61773) );
  INVX1 U65735 ( .A(n61773), .Y(n61721) );
  XNOR2X1 U65736 ( .A(n61609), .B(n38017), .Y(n61610) );
  XNOR2X1 U65737 ( .A(n41971), .B(n61610), .Y(n61775) );
  INVX1 U65738 ( .A(n61775), .Y(n61716) );
  XNOR2X1 U65739 ( .A(n61611), .B(n39830), .Y(n61612) );
  XNOR2X1 U65740 ( .A(n41961), .B(n61612), .Y(n61777) );
  XNOR2X1 U65741 ( .A(n61614), .B(n61613), .Y(n61615) );
  XNOR2X1 U65742 ( .A(n41952), .B(n61615), .Y(n61780) );
  INVX1 U65743 ( .A(n61780), .Y(n61709) );
  XNOR2X1 U65744 ( .A(n61616), .B(n38453), .Y(n61617) );
  XNOR2X1 U65745 ( .A(n41941), .B(n61617), .Y(n61783) );
  INVX1 U65746 ( .A(n61783), .Y(n61706) );
  XNOR2X1 U65747 ( .A(n61618), .B(n39642), .Y(n61619) );
  XNOR2X1 U65748 ( .A(n41931), .B(n61619), .Y(n61786) );
  XNOR2X1 U65749 ( .A(n61621), .B(n61620), .Y(n61622) );
  XNOR2X1 U65750 ( .A(n41920), .B(n61622), .Y(n61789) );
  INVX1 U65751 ( .A(n61789), .Y(n61698) );
  XNOR2X1 U65752 ( .A(n61623), .B(n39400), .Y(n61624) );
  XNOR2X1 U65753 ( .A(n41909), .B(n61624), .Y(n61792) );
  XNOR2X1 U65754 ( .A(n61625), .B(n38993), .Y(n61626) );
  XNOR2X1 U65755 ( .A(n41899), .B(n61626), .Y(n61795) );
  INVX1 U65756 ( .A(n61795), .Y(n61691) );
  XNOR2X1 U65757 ( .A(n61628), .B(n61627), .Y(n61629) );
  XNOR2X1 U65758 ( .A(n41888), .B(n61629), .Y(n61798) );
  XNOR2X1 U65759 ( .A(n61631), .B(n61630), .Y(n61632) );
  XNOR2X1 U65760 ( .A(n41877), .B(n61632), .Y(n61801) );
  INVX1 U65761 ( .A(n61801), .Y(n61682) );
  XNOR2X1 U65762 ( .A(n61634), .B(n61633), .Y(n61635) );
  XNOR2X1 U65763 ( .A(n41867), .B(n61635), .Y(n61804) );
  XNOR2X1 U65764 ( .A(n61636), .B(n38761), .Y(n61637) );
  XNOR2X1 U65765 ( .A(n41852), .B(n61637), .Y(n61807) );
  INVX1 U65766 ( .A(n61807), .Y(n61673) );
  XNOR2X1 U65767 ( .A(n61638), .B(n41837), .Y(n61639) );
  XNOR2X1 U65768 ( .A(n61640), .B(n61639), .Y(n61810) );
  XNOR2X1 U65769 ( .A(n61642), .B(n61641), .Y(n61643) );
  XNOR2X1 U65770 ( .A(n41822), .B(n61643), .Y(n61812) );
  INVX1 U65771 ( .A(n61812), .Y(n61665) );
  XNOR2X1 U65772 ( .A(n61644), .B(n36397), .Y(n61645) );
  XNOR2X1 U65773 ( .A(n41810), .B(n61645), .Y(n61815) );
  XNOR2X1 U65774 ( .A(n61647), .B(n61646), .Y(n61648) );
  XNOR2X1 U65775 ( .A(n41789), .B(n61648), .Y(n61819) );
  INVX1 U65776 ( .A(n61819), .Y(n61656) );
  NAND2X1 U65777 ( .A(n42715), .B(n43765), .Y(n61824) );
  NAND2X1 U65778 ( .A(n40390), .B(n43743), .Y(n61825) );
  INVX1 U65779 ( .A(n61826), .Y(n61821) );
  NAND2X1 U65780 ( .A(n61650), .B(n61649), .Y(n61652) );
  NAND2X1 U65781 ( .A(n61651), .B(n61652), .Y(n61822) );
  NAND2X1 U65782 ( .A(n61821), .B(n37405), .Y(n61655) );
  NAND2X1 U65783 ( .A(n61822), .B(n61826), .Y(n61653) );
  NAND2X1 U65784 ( .A(n41804), .B(n61653), .Y(n61654) );
  NAND2X1 U65785 ( .A(n61655), .B(n61654), .Y(n61657) );
  NAND2X1 U65786 ( .A(n61656), .B(n61657), .Y(n61660) );
  INVX1 U65787 ( .A(n61657), .Y(n61818) );
  NAND2X1 U65788 ( .A(n61818), .B(n61819), .Y(n61658) );
  NAND2X1 U65789 ( .A(n41817), .B(n61658), .Y(n61659) );
  NAND2X1 U65790 ( .A(n61660), .B(n61659), .Y(n61662) );
  INVX1 U65791 ( .A(n61661), .Y(n61814) );
  INVX1 U65792 ( .A(n61662), .Y(n61817) );
  INVX1 U65793 ( .A(n61815), .Y(n61663) );
  NAND2X1 U65794 ( .A(n61817), .B(n61663), .Y(n61664) );
  NAND2X1 U65795 ( .A(n61665), .B(n61666), .Y(n61669) );
  NAND2X1 U65796 ( .A(n41845), .B(n61667), .Y(n61668) );
  NAND2X1 U65797 ( .A(n61669), .B(n61668), .Y(n61670) );
  INVX1 U65798 ( .A(n61670), .Y(n61809) );
  INVX1 U65799 ( .A(n61810), .Y(n61671) );
  NAND2X1 U65800 ( .A(n61809), .B(n61671), .Y(n61672) );
  NAND2X1 U65801 ( .A(n61673), .B(n61674), .Y(n61677) );
  INVX1 U65802 ( .A(n61674), .Y(n61806) );
  NAND2X1 U65803 ( .A(n41871), .B(n61675), .Y(n61676) );
  NAND2X1 U65804 ( .A(n61677), .B(n61676), .Y(n61678) );
  NAND2X1 U65805 ( .A(n61804), .B(n61678), .Y(n61681) );
  INVX1 U65806 ( .A(n61678), .Y(n61803) );
  INVX1 U65807 ( .A(n61804), .Y(n61679) );
  NAND2X1 U65808 ( .A(n61681), .B(n61680), .Y(n61683) );
  NAND2X1 U65809 ( .A(n61682), .B(n61683), .Y(n61685) );
  INVX1 U65810 ( .A(n61683), .Y(n61800) );
  NAND2X1 U65811 ( .A(n61685), .B(n61684), .Y(n61686) );
  NAND2X1 U65812 ( .A(n61798), .B(n61686), .Y(n61690) );
  INVX1 U65813 ( .A(n61686), .Y(n61797) );
  INVX1 U65814 ( .A(n61798), .Y(n61687) );
  NAND2X1 U65815 ( .A(n61797), .B(n61687), .Y(n61688) );
  NAND2X1 U65816 ( .A(n41903), .B(n61688), .Y(n61689) );
  NAND2X1 U65817 ( .A(n61690), .B(n61689), .Y(n61692) );
  NAND2X1 U65818 ( .A(n61691), .B(n61692), .Y(n61695) );
  INVX1 U65819 ( .A(n61692), .Y(n61794) );
  NAND2X1 U65820 ( .A(n61794), .B(n61795), .Y(n61693) );
  NAND2X1 U65821 ( .A(n41914), .B(n61693), .Y(n61694) );
  NAND2X1 U65822 ( .A(n61695), .B(n61694), .Y(n61696) );
  INVX1 U65823 ( .A(n61696), .Y(n61791) );
  NAND2X1 U65824 ( .A(n61698), .B(n61699), .Y(n61702) );
  INVX1 U65825 ( .A(n61699), .Y(n61788) );
  NAND2X1 U65826 ( .A(n41933), .B(n61700), .Y(n61701) );
  NAND2X1 U65827 ( .A(n61702), .B(n61701), .Y(n61703) );
  INVX1 U65828 ( .A(n61703), .Y(n61785) );
  INVX1 U65829 ( .A(n61786), .Y(n61704) );
  NAND2X1 U65830 ( .A(n61785), .B(n61704), .Y(n61705) );
  INVX1 U65831 ( .A(n61707), .Y(n61782) );
  INVX1 U65832 ( .A(n61710), .Y(n61779) );
  NAND2X1 U65833 ( .A(n61777), .B(n61712), .Y(n61715) );
  INVX1 U65834 ( .A(n61777), .Y(n61713) );
  NAND2X1 U65835 ( .A(n61715), .B(n61714), .Y(n61717) );
  NAND2X1 U65836 ( .A(n61716), .B(n61717), .Y(n61720) );
  NAND2X1 U65837 ( .A(n36416), .B(n61775), .Y(n61718) );
  NAND2X1 U65838 ( .A(n41984), .B(n61718), .Y(n61719) );
  NAND2X1 U65839 ( .A(n61720), .B(n61719), .Y(n61722) );
  NAND2X1 U65840 ( .A(n61724), .B(n61725), .Y(n61727) );
  INVX1 U65841 ( .A(n61725), .Y(n61770) );
  NAND2X1 U65842 ( .A(n61727), .B(n61726), .Y(n61728) );
  INVX1 U65843 ( .A(n61728), .Y(n61767) );
  INVX1 U65844 ( .A(n61768), .Y(n61729) );
  NAND2X1 U65845 ( .A(n61730), .B(n61731), .Y(n61733) );
  INVX1 U65846 ( .A(n61731), .Y(n61764) );
  NAND2X1 U65847 ( .A(n61733), .B(n61732), .Y(n61734) );
  INVX1 U65848 ( .A(n61734), .Y(n61761) );
  INVX1 U65849 ( .A(n61759), .Y(n61737) );
  NAND2X1 U65850 ( .A(n36347), .B(n61737), .Y(n61738) );
  NAND2X1 U65851 ( .A(n61739), .B(n61740), .Y(n61742) );
  INVX1 U65852 ( .A(n61740), .Y(n61756) );
  NAND2X1 U65853 ( .A(n61742), .B(n61741), .Y(n61744) );
  NAND2X1 U65854 ( .A(n61743), .B(n61744), .Y(n61747) );
  INVX1 U65855 ( .A(n61744), .Y(n61753) );
  NAND2X1 U65856 ( .A(n61754), .B(n61753), .Y(n61745) );
  NAND2X1 U65857 ( .A(n42076), .B(n61745), .Y(n61746) );
  NAND2X1 U65858 ( .A(n61747), .B(n61746), .Y(n61748) );
  INVX1 U65859 ( .A(n61748), .Y(n61750) );
  XNOR2X1 U65860 ( .A(n62564), .B(n38250), .Y(n61749) );
  XNOR2X1 U65861 ( .A(n42095), .B(n61749), .Y(n62335) );
  XNOR2X1 U65862 ( .A(n61751), .B(n61750), .Y(n61752) );
  XNOR2X1 U65863 ( .A(n42086), .B(n61752), .Y(n61942) );
  INVX1 U65864 ( .A(n61942), .Y(n61937) );
  XNOR2X1 U65865 ( .A(n61754), .B(n61753), .Y(n61755) );
  XNOR2X1 U65866 ( .A(n42076), .B(n61755), .Y(n61945) );
  XNOR2X1 U65867 ( .A(n61757), .B(n61756), .Y(n61758) );
  XNOR2X1 U65868 ( .A(n42065), .B(n61758), .Y(n61947) );
  XNOR2X1 U65869 ( .A(n61759), .B(n36347), .Y(n61760) );
  XNOR2X1 U65870 ( .A(n42054), .B(n61760), .Y(n61949) );
  INVX1 U65871 ( .A(n61949), .Y(n61926) );
  XNOR2X1 U65872 ( .A(n61762), .B(n61761), .Y(n61763) );
  XNOR2X1 U65873 ( .A(n42042), .B(n61763), .Y(n61951) );
  INVX1 U65874 ( .A(n61951), .Y(n61921) );
  XNOR2X1 U65875 ( .A(n61765), .B(n61764), .Y(n61766) );
  XNOR2X1 U65876 ( .A(n42030), .B(n61766), .Y(n61953) );
  XNOR2X1 U65877 ( .A(n61768), .B(n61767), .Y(n61769) );
  XNOR2X1 U65878 ( .A(n42018), .B(n61769), .Y(n61956) );
  INVX1 U65879 ( .A(n61956), .Y(n61913) );
  XNOR2X1 U65880 ( .A(n61771), .B(n61770), .Y(n61772) );
  XNOR2X1 U65881 ( .A(n42008), .B(n61772), .Y(n61958) );
  XNOR2X1 U65882 ( .A(n61773), .B(n36418), .Y(n61774) );
  XNOR2X1 U65883 ( .A(n41995), .B(n61774), .Y(n61960) );
  XNOR2X1 U65884 ( .A(n61775), .B(n36416), .Y(n61776) );
  XNOR2X1 U65885 ( .A(n41984), .B(n61776), .Y(n61962) );
  XNOR2X1 U65886 ( .A(n61777), .B(n36413), .Y(n61778) );
  XNOR2X1 U65887 ( .A(n41974), .B(n61778), .Y(n61965) );
  INVX1 U65888 ( .A(n61965), .Y(n61898) );
  XNOR2X1 U65889 ( .A(n61780), .B(n61779), .Y(n61781) );
  XNOR2X1 U65890 ( .A(n41963), .B(n61781), .Y(n61967) );
  XNOR2X1 U65891 ( .A(n61783), .B(n61782), .Y(n61784) );
  XNOR2X1 U65892 ( .A(n41954), .B(n61784), .Y(n61969) );
  XNOR2X1 U65893 ( .A(n61786), .B(n61785), .Y(n61787) );
  XNOR2X1 U65894 ( .A(n41945), .B(n61787), .Y(n61972) );
  INVX1 U65895 ( .A(n61972), .Y(n61885) );
  XNOR2X1 U65896 ( .A(n61789), .B(n61788), .Y(n61790) );
  XNOR2X1 U65897 ( .A(n41933), .B(n61790), .Y(n61974) );
  XNOR2X1 U65898 ( .A(n61792), .B(n61791), .Y(n61793) );
  XNOR2X1 U65899 ( .A(n41924), .B(n61793), .Y(n61977) );
  INVX1 U65900 ( .A(n61977), .Y(n61878) );
  XNOR2X1 U65901 ( .A(n61795), .B(n61794), .Y(n61796) );
  XNOR2X1 U65902 ( .A(n41914), .B(n61796), .Y(n61980) );
  XNOR2X1 U65903 ( .A(n61798), .B(n61797), .Y(n61799) );
  XNOR2X1 U65904 ( .A(n41903), .B(n61799), .Y(n61983) );
  INVX1 U65905 ( .A(n61983), .Y(n61868) );
  XNOR2X1 U65906 ( .A(n61801), .B(n61800), .Y(n61802) );
  XNOR2X1 U65907 ( .A(n41891), .B(n61802), .Y(n61986) );
  XNOR2X1 U65908 ( .A(n61804), .B(n61803), .Y(n61805) );
  XNOR2X1 U65909 ( .A(n41882), .B(n61805), .Y(n61989) );
  INVX1 U65910 ( .A(n61989), .Y(n61858) );
  XNOR2X1 U65911 ( .A(n61807), .B(n61806), .Y(n61808) );
  XNOR2X1 U65912 ( .A(n41871), .B(n61808), .Y(n61992) );
  XNOR2X1 U65913 ( .A(n61810), .B(n61809), .Y(n61811) );
  XNOR2X1 U65914 ( .A(n41861), .B(n61811), .Y(n61994) );
  INVX1 U65915 ( .A(n61994), .Y(n61848) );
  XNOR2X1 U65916 ( .A(n61812), .B(n38445), .Y(n61813) );
  XNOR2X1 U65917 ( .A(n41845), .B(n61813), .Y(n61997) );
  XNOR2X1 U65918 ( .A(n61815), .B(n61814), .Y(n61816) );
  XNOR2X1 U65919 ( .A(n61817), .B(n61816), .Y(n61999) );
  INVX1 U65920 ( .A(n61999), .Y(n61840) );
  XNOR2X1 U65921 ( .A(n61819), .B(n61818), .Y(n61820) );
  XNOR2X1 U65922 ( .A(n41817), .B(n61820), .Y(n62002) );
  XNOR2X1 U65923 ( .A(n61822), .B(n61821), .Y(n61823) );
  XNOR2X1 U65924 ( .A(n41804), .B(n61823), .Y(n62004) );
  INVX1 U65925 ( .A(n62004), .Y(n61832) );
  NAND2X1 U65926 ( .A(n43802), .B(n42719), .Y(n62010) );
  NAND2X1 U65927 ( .A(n44070), .B(n43765), .Y(n62011) );
  INVX1 U65928 ( .A(n62012), .Y(n62007) );
  NAND2X1 U65929 ( .A(n61825), .B(n61824), .Y(n61827) );
  NAND2X1 U65930 ( .A(n61827), .B(n61826), .Y(n62008) );
  INVX1 U65931 ( .A(n62008), .Y(n61828) );
  NAND2X1 U65932 ( .A(n62007), .B(n61828), .Y(n61831) );
  NAND2X1 U65933 ( .A(n62012), .B(n62008), .Y(n61829) );
  NAND2X1 U65934 ( .A(n41820), .B(n61829), .Y(n61830) );
  NAND2X1 U65935 ( .A(n61831), .B(n61830), .Y(n61833) );
  NAND2X1 U65936 ( .A(n61832), .B(n61833), .Y(n61836) );
  INVX1 U65937 ( .A(n61833), .Y(n62006) );
  NAND2X1 U65938 ( .A(n62006), .B(n62004), .Y(n61834) );
  NAND2X1 U65939 ( .A(n41836), .B(n61834), .Y(n61835) );
  NAND2X1 U65940 ( .A(n61836), .B(n61835), .Y(n61837) );
  INVX1 U65941 ( .A(n61837), .Y(n62001) );
  INVX1 U65942 ( .A(n62002), .Y(n61838) );
  NAND2X1 U65943 ( .A(n62001), .B(n61838), .Y(n61839) );
  NAND2X1 U65944 ( .A(n61840), .B(n61841), .Y(n61844) );
  NAND2X1 U65945 ( .A(n38286), .B(n61999), .Y(n61842) );
  NAND2X1 U65946 ( .A(n41865), .B(n61842), .Y(n61843) );
  NAND2X1 U65947 ( .A(n61844), .B(n61843), .Y(n61845) );
  INVX1 U65948 ( .A(n61845), .Y(n61996) );
  INVX1 U65949 ( .A(n61997), .Y(n61846) );
  NAND2X1 U65950 ( .A(n61996), .B(n61846), .Y(n61847) );
  NAND2X1 U65951 ( .A(n61848), .B(n61849), .Y(n61852) );
  NAND2X1 U65952 ( .A(n36370), .B(n61994), .Y(n61850) );
  NAND2X1 U65953 ( .A(n41886), .B(n61850), .Y(n61851) );
  NAND2X1 U65954 ( .A(n61852), .B(n61851), .Y(n61853) );
  NAND2X1 U65955 ( .A(n61992), .B(n61853), .Y(n61857) );
  INVX1 U65956 ( .A(n61853), .Y(n61991) );
  INVX1 U65957 ( .A(n61992), .Y(n61854) );
  NAND2X1 U65958 ( .A(n61991), .B(n61854), .Y(n61855) );
  NAND2X1 U65959 ( .A(n41897), .B(n61855), .Y(n61856) );
  NAND2X1 U65960 ( .A(n61857), .B(n61856), .Y(n61859) );
  NAND2X1 U65961 ( .A(n61858), .B(n61859), .Y(n61862) );
  INVX1 U65962 ( .A(n61859), .Y(n61988) );
  NAND2X1 U65963 ( .A(n61988), .B(n61989), .Y(n61860) );
  NAND2X1 U65964 ( .A(n41907), .B(n61860), .Y(n61861) );
  NAND2X1 U65965 ( .A(n61862), .B(n61861), .Y(n61863) );
  NAND2X1 U65966 ( .A(n61986), .B(n61863), .Y(n61867) );
  INVX1 U65967 ( .A(n61863), .Y(n61985) );
  INVX1 U65968 ( .A(n61986), .Y(n61864) );
  NAND2X1 U65969 ( .A(n61985), .B(n61864), .Y(n61865) );
  NAND2X1 U65970 ( .A(n41919), .B(n61865), .Y(n61866) );
  NAND2X1 U65971 ( .A(n61867), .B(n61866), .Y(n61869) );
  NAND2X1 U65972 ( .A(n61868), .B(n61869), .Y(n61872) );
  INVX1 U65973 ( .A(n61869), .Y(n61982) );
  NAND2X1 U65974 ( .A(n61982), .B(n61983), .Y(n61870) );
  NAND2X1 U65975 ( .A(n41929), .B(n61870), .Y(n61871) );
  NAND2X1 U65976 ( .A(n61872), .B(n61871), .Y(n61873) );
  NAND2X1 U65977 ( .A(n61980), .B(n61873), .Y(n61877) );
  INVX1 U65978 ( .A(n61873), .Y(n61979) );
  INVX1 U65979 ( .A(n61980), .Y(n61874) );
  NAND2X1 U65980 ( .A(n61979), .B(n61874), .Y(n61875) );
  NAND2X1 U65981 ( .A(n41939), .B(n61875), .Y(n61876) );
  NAND2X1 U65982 ( .A(n61877), .B(n61876), .Y(n61879) );
  INVX1 U65983 ( .A(n61879), .Y(n61976) );
  NAND2X1 U65984 ( .A(n61976), .B(n61977), .Y(n61880) );
  NAND2X1 U65985 ( .A(n61974), .B(n36377), .Y(n61884) );
  INVX1 U65986 ( .A(n61974), .Y(n61881) );
  NAND2X1 U65987 ( .A(n38429), .B(n61881), .Y(n61882) );
  NAND2X1 U65988 ( .A(n41960), .B(n61882), .Y(n61883) );
  NAND2X1 U65989 ( .A(n61884), .B(n61883), .Y(n61886) );
  INVX1 U65990 ( .A(n61886), .Y(n61971) );
  NAND2X1 U65991 ( .A(n61971), .B(n61972), .Y(n61887) );
  NAND2X1 U65992 ( .A(n61969), .B(n61888), .Y(n61892) );
  INVX1 U65993 ( .A(n61969), .Y(n61889) );
  NAND2X1 U65994 ( .A(n41980), .B(n61890), .Y(n61891) );
  NAND2X1 U65995 ( .A(n61892), .B(n61891), .Y(n61893) );
  NAND2X1 U65996 ( .A(n61967), .B(n61893), .Y(n61897) );
  INVX1 U65997 ( .A(n61967), .Y(n61894) );
  NAND2X1 U65998 ( .A(n36440), .B(n61894), .Y(n61895) );
  NAND2X1 U65999 ( .A(n41989), .B(n61895), .Y(n61896) );
  NAND2X1 U66000 ( .A(n61897), .B(n61896), .Y(n61899) );
  INVX1 U66001 ( .A(n61899), .Y(n61964) );
  NAND2X1 U66002 ( .A(n61964), .B(n61965), .Y(n61900) );
  NAND2X1 U66003 ( .A(n61962), .B(n61901), .Y(n61905) );
  INVX1 U66004 ( .A(n61962), .Y(n61902) );
  NAND2X1 U66005 ( .A(n42013), .B(n61903), .Y(n61904) );
  NAND2X1 U66006 ( .A(n61905), .B(n61904), .Y(n61906) );
  INVX1 U66007 ( .A(n61960), .Y(n61907) );
  NAND2X1 U66008 ( .A(n36382), .B(n61907), .Y(n61908) );
  NAND2X1 U66009 ( .A(n61958), .B(n38132), .Y(n61912) );
  INVX1 U66010 ( .A(n61958), .Y(n61909) );
  NAND2X1 U66011 ( .A(n38306), .B(n61909), .Y(n61910) );
  NAND2X1 U66012 ( .A(n42037), .B(n61910), .Y(n61911) );
  NAND2X1 U66013 ( .A(n61912), .B(n61911), .Y(n61914) );
  INVX1 U66014 ( .A(n61914), .Y(n61955) );
  NAND2X1 U66015 ( .A(n61955), .B(n61956), .Y(n61915) );
  NAND2X1 U66016 ( .A(n61953), .B(n61916), .Y(n61920) );
  INVX1 U66017 ( .A(n61953), .Y(n61917) );
  NAND2X1 U66018 ( .A(n42060), .B(n61918), .Y(n61919) );
  NAND2X1 U66019 ( .A(n61920), .B(n61919), .Y(n61922) );
  NAND2X1 U66020 ( .A(n61921), .B(n61922), .Y(n61925) );
  NAND2X1 U66021 ( .A(n37950), .B(n61951), .Y(n61923) );
  NAND2X1 U66022 ( .A(n42072), .B(n61923), .Y(n61924) );
  NAND2X1 U66023 ( .A(n61925), .B(n61924), .Y(n61927) );
  NAND2X1 U66024 ( .A(n36396), .B(n61949), .Y(n61928) );
  NAND2X1 U66025 ( .A(n61947), .B(n61929), .Y(n61933) );
  INVX1 U66026 ( .A(n61947), .Y(n61930) );
  NAND2X1 U66027 ( .A(n42092), .B(n61931), .Y(n61932) );
  NAND2X1 U66028 ( .A(n61933), .B(n61932), .Y(n61934) );
  INVX1 U66029 ( .A(n61934), .Y(n61944) );
  INVX1 U66030 ( .A(n61945), .Y(n61935) );
  NAND2X1 U66031 ( .A(n61944), .B(n61935), .Y(n61936) );
  NAND2X1 U66032 ( .A(n61937), .B(n37958), .Y(n61940) );
  NAND2X1 U66033 ( .A(n38056), .B(n61942), .Y(n61938) );
  NAND2X1 U66034 ( .A(n42105), .B(n61938), .Y(n61939) );
  NAND2X1 U66035 ( .A(n61940), .B(n61939), .Y(n62333) );
  XNOR2X1 U66036 ( .A(n62335), .B(n37951), .Y(n61941) );
  XNOR2X1 U66037 ( .A(n42112), .B(n61941), .Y(n62571) );
  XNOR2X1 U66038 ( .A(n61942), .B(n38056), .Y(n61943) );
  XNOR2X1 U66039 ( .A(n42105), .B(n61943), .Y(n62133) );
  XNOR2X1 U66040 ( .A(n61945), .B(n61944), .Y(n61946) );
  XNOR2X1 U66041 ( .A(n42099), .B(n61946), .Y(n62135) );
  INVX1 U66042 ( .A(n62135), .Y(n62124) );
  XNOR2X1 U66043 ( .A(n61947), .B(n39472), .Y(n61948) );
  XNOR2X1 U66044 ( .A(n42092), .B(n61948), .Y(n62137) );
  XNOR2X1 U66045 ( .A(n61949), .B(n36396), .Y(n61950) );
  XNOR2X1 U66046 ( .A(n42081), .B(n61950), .Y(n62139) );
  XNOR2X1 U66047 ( .A(n61951), .B(n37950), .Y(n61952) );
  XNOR2X1 U66048 ( .A(n42072), .B(n61952), .Y(n62141) );
  XNOR2X1 U66049 ( .A(n61953), .B(n39289), .Y(n61954) );
  XNOR2X1 U66050 ( .A(n42060), .B(n61954), .Y(n62144) );
  INVX1 U66051 ( .A(n62144), .Y(n62112) );
  XNOR2X1 U66052 ( .A(n61956), .B(n61955), .Y(n61957) );
  XNOR2X1 U66053 ( .A(n42050), .B(n61957), .Y(n62146) );
  XNOR2X1 U66054 ( .A(n61958), .B(n38306), .Y(n61959) );
  XNOR2X1 U66055 ( .A(n42037), .B(n61959), .Y(n62149) );
  INVX1 U66056 ( .A(n62149), .Y(n62104) );
  XNOR2X1 U66057 ( .A(n61960), .B(n36382), .Y(n61961) );
  XNOR2X1 U66058 ( .A(n42023), .B(n61961), .Y(n62152) );
  INVX1 U66059 ( .A(n62152), .Y(n62099) );
  XNOR2X1 U66060 ( .A(n61962), .B(n39062), .Y(n61963) );
  XNOR2X1 U66061 ( .A(n42013), .B(n61963), .Y(n62155) );
  INVX1 U66062 ( .A(n62155), .Y(n62094) );
  XNOR2X1 U66063 ( .A(n61965), .B(n61964), .Y(n61966) );
  XNOR2X1 U66064 ( .A(n42002), .B(n61966), .Y(n62158) );
  XNOR2X1 U66065 ( .A(n61967), .B(n36440), .Y(n61968) );
  XNOR2X1 U66066 ( .A(n41989), .B(n61968), .Y(n62161) );
  INVX1 U66067 ( .A(n62161), .Y(n62085) );
  XNOR2X1 U66068 ( .A(n61969), .B(n38814), .Y(n61970) );
  XNOR2X1 U66069 ( .A(n41980), .B(n61970), .Y(n62163) );
  INVX1 U66070 ( .A(n62163), .Y(n62080) );
  XNOR2X1 U66071 ( .A(n61972), .B(n61971), .Y(n61973) );
  XNOR2X1 U66072 ( .A(n41970), .B(n61973), .Y(n62165) );
  XNOR2X1 U66073 ( .A(n61974), .B(n38429), .Y(n61975) );
  XNOR2X1 U66074 ( .A(n41960), .B(n61975), .Y(n62168) );
  INVX1 U66075 ( .A(n62168), .Y(n62073) );
  XNOR2X1 U66076 ( .A(n61977), .B(n61976), .Y(n61978) );
  XNOR2X1 U66077 ( .A(n41951), .B(n61978), .Y(n62171) );
  XNOR2X1 U66078 ( .A(n61980), .B(n61979), .Y(n61981) );
  XNOR2X1 U66079 ( .A(n41939), .B(n61981), .Y(n62174) );
  INVX1 U66080 ( .A(n62174), .Y(n62063) );
  XNOR2X1 U66081 ( .A(n61983), .B(n61982), .Y(n61984) );
  XNOR2X1 U66082 ( .A(n41929), .B(n61984), .Y(n62177) );
  XNOR2X1 U66083 ( .A(n61986), .B(n61985), .Y(n61987) );
  XNOR2X1 U66084 ( .A(n41919), .B(n61987), .Y(n62179) );
  INVX1 U66085 ( .A(n62179), .Y(n62053) );
  XNOR2X1 U66086 ( .A(n61989), .B(n61988), .Y(n61990) );
  XNOR2X1 U66087 ( .A(n41907), .B(n61990), .Y(n62182) );
  XNOR2X1 U66088 ( .A(n61992), .B(n61991), .Y(n61993) );
  XNOR2X1 U66089 ( .A(n41897), .B(n61993), .Y(n62185) );
  INVX1 U66090 ( .A(n62185), .Y(n62046) );
  XNOR2X1 U66091 ( .A(n61994), .B(n36370), .Y(n61995) );
  XNOR2X1 U66092 ( .A(n41886), .B(n61995), .Y(n62188) );
  XNOR2X1 U66093 ( .A(n61997), .B(n61996), .Y(n61998) );
  XNOR2X1 U66094 ( .A(n41875), .B(n61998), .Y(n62191) );
  INVX1 U66095 ( .A(n62191), .Y(n62036) );
  XNOR2X1 U66096 ( .A(n61999), .B(n38286), .Y(n62000) );
  XNOR2X1 U66097 ( .A(n41865), .B(n62000), .Y(n62194) );
  XNOR2X1 U66098 ( .A(n62002), .B(n62001), .Y(n62003) );
  XNOR2X1 U66099 ( .A(n41850), .B(n62003), .Y(n62197) );
  INVX1 U66100 ( .A(n62197), .Y(n62026) );
  XNOR2X1 U66101 ( .A(n62004), .B(n41836), .Y(n62005) );
  XNOR2X1 U66102 ( .A(n62006), .B(n62005), .Y(n62200) );
  XNOR2X1 U66103 ( .A(n62008), .B(n62007), .Y(n62009) );
  XNOR2X1 U66104 ( .A(n41820), .B(n62009), .Y(n62202) );
  INVX1 U66105 ( .A(n62202), .Y(n62016) );
  NAND2X1 U66106 ( .A(n42717), .B(n72823), .Y(n62207) );
  NAND2X1 U66107 ( .A(n43802), .B(n44070), .Y(n62208) );
  INVX1 U66108 ( .A(n62209), .Y(n62206) );
  NAND2X1 U66109 ( .A(n62011), .B(n62010), .Y(n62013) );
  INVX1 U66110 ( .A(n62014), .Y(n62204) );
  NAND2X1 U66111 ( .A(n62209), .B(n38112), .Y(n62015) );
  NAND2X1 U66112 ( .A(n62016), .B(n62017), .Y(n62020) );
  NAND2X1 U66113 ( .A(n38040), .B(n62202), .Y(n62018) );
  NAND2X1 U66114 ( .A(n41848), .B(n62018), .Y(n62019) );
  NAND2X1 U66115 ( .A(n62020), .B(n62019), .Y(n62021) );
  NAND2X1 U66116 ( .A(n62200), .B(n62021), .Y(n62025) );
  INVX1 U66117 ( .A(n62021), .Y(n62199) );
  INVX1 U66118 ( .A(n62200), .Y(n62022) );
  NAND2X1 U66119 ( .A(n62199), .B(n62022), .Y(n62023) );
  NAND2X1 U66120 ( .A(n41864), .B(n62023), .Y(n62024) );
  NAND2X1 U66121 ( .A(n62025), .B(n62024), .Y(n62027) );
  NAND2X1 U66122 ( .A(n62026), .B(n62027), .Y(n62030) );
  INVX1 U66123 ( .A(n62027), .Y(n62196) );
  NAND2X1 U66124 ( .A(n62196), .B(n62197), .Y(n62028) );
  NAND2X1 U66125 ( .A(n41874), .B(n62028), .Y(n62029) );
  NAND2X1 U66126 ( .A(n62030), .B(n62029), .Y(n62031) );
  NAND2X1 U66127 ( .A(n62194), .B(n62031), .Y(n62035) );
  INVX1 U66128 ( .A(n62031), .Y(n62193) );
  INVX1 U66129 ( .A(n62194), .Y(n62032) );
  NAND2X1 U66130 ( .A(n62193), .B(n62032), .Y(n62033) );
  NAND2X1 U66131 ( .A(n41885), .B(n62033), .Y(n62034) );
  NAND2X1 U66132 ( .A(n62035), .B(n62034), .Y(n62037) );
  NAND2X1 U66133 ( .A(n62036), .B(n62037), .Y(n62040) );
  INVX1 U66134 ( .A(n62037), .Y(n62190) );
  NAND2X1 U66135 ( .A(n62190), .B(n62191), .Y(n62038) );
  NAND2X1 U66136 ( .A(n41896), .B(n62038), .Y(n62039) );
  NAND2X1 U66137 ( .A(n62040), .B(n62039), .Y(n62041) );
  NAND2X1 U66138 ( .A(n62188), .B(n62041), .Y(n62045) );
  INVX1 U66139 ( .A(n62041), .Y(n62187) );
  INVX1 U66140 ( .A(n62188), .Y(n62042) );
  NAND2X1 U66141 ( .A(n62187), .B(n62042), .Y(n62043) );
  NAND2X1 U66142 ( .A(n41906), .B(n62043), .Y(n62044) );
  NAND2X1 U66143 ( .A(n62045), .B(n62044), .Y(n62047) );
  NAND2X1 U66144 ( .A(n62046), .B(n62047), .Y(n62050) );
  INVX1 U66145 ( .A(n62047), .Y(n62184) );
  NAND2X1 U66146 ( .A(n62184), .B(n62185), .Y(n62048) );
  NAND2X1 U66147 ( .A(n41917), .B(n62048), .Y(n62049) );
  NAND2X1 U66148 ( .A(n62050), .B(n62049), .Y(n62051) );
  INVX1 U66149 ( .A(n62051), .Y(n62181) );
  INVX1 U66150 ( .A(n62182), .Y(n62052) );
  NAND2X1 U66151 ( .A(n62053), .B(n62054), .Y(n62057) );
  NAND2X1 U66152 ( .A(n36398), .B(n62179), .Y(n62055) );
  NAND2X1 U66153 ( .A(n41937), .B(n62055), .Y(n62056) );
  NAND2X1 U66154 ( .A(n62057), .B(n62056), .Y(n62058) );
  NAND2X1 U66155 ( .A(n62177), .B(n62058), .Y(n62062) );
  INVX1 U66156 ( .A(n62058), .Y(n62176) );
  INVX1 U66157 ( .A(n62177), .Y(n62059) );
  NAND2X1 U66158 ( .A(n62176), .B(n62059), .Y(n62060) );
  NAND2X1 U66159 ( .A(n41949), .B(n62060), .Y(n62061) );
  NAND2X1 U66160 ( .A(n62062), .B(n62061), .Y(n62064) );
  NAND2X1 U66161 ( .A(n62063), .B(n62064), .Y(n62067) );
  INVX1 U66162 ( .A(n62064), .Y(n62173) );
  NAND2X1 U66163 ( .A(n62173), .B(n62174), .Y(n62065) );
  NAND2X1 U66164 ( .A(n41958), .B(n62065), .Y(n62066) );
  NAND2X1 U66165 ( .A(n62067), .B(n62066), .Y(n62068) );
  NAND2X1 U66166 ( .A(n62171), .B(n62068), .Y(n62072) );
  INVX1 U66167 ( .A(n62068), .Y(n62170) );
  INVX1 U66168 ( .A(n62171), .Y(n62069) );
  NAND2X1 U66169 ( .A(n62170), .B(n62069), .Y(n62070) );
  NAND2X1 U66170 ( .A(n41968), .B(n62070), .Y(n62071) );
  NAND2X1 U66171 ( .A(n62072), .B(n62071), .Y(n62074) );
  INVX1 U66172 ( .A(n62074), .Y(n62167) );
  NAND2X1 U66173 ( .A(n62167), .B(n62168), .Y(n62075) );
  NAND2X1 U66174 ( .A(n62165), .B(n38113), .Y(n62079) );
  INVX1 U66175 ( .A(n62165), .Y(n62076) );
  NAND2X1 U66176 ( .A(n38276), .B(n62076), .Y(n62077) );
  NAND2X1 U66177 ( .A(n41987), .B(n62077), .Y(n62078) );
  NAND2X1 U66178 ( .A(n62079), .B(n62078), .Y(n62081) );
  NAND2X1 U66179 ( .A(n62080), .B(n62081), .Y(n62084) );
  NAND2X1 U66180 ( .A(n38063), .B(n62163), .Y(n62082) );
  NAND2X1 U66181 ( .A(n42000), .B(n62082), .Y(n62083) );
  NAND2X1 U66182 ( .A(n62084), .B(n62083), .Y(n62086) );
  NAND2X1 U66183 ( .A(n62085), .B(n62086), .Y(n62089) );
  INVX1 U66184 ( .A(n62086), .Y(n62160) );
  NAND2X1 U66185 ( .A(n62160), .B(n62161), .Y(n62087) );
  NAND2X1 U66186 ( .A(n42011), .B(n62087), .Y(n62088) );
  NAND2X1 U66187 ( .A(n62089), .B(n62088), .Y(n62090) );
  NAND2X1 U66188 ( .A(n62158), .B(n62090), .Y(n62093) );
  INVX1 U66189 ( .A(n62090), .Y(n62157) );
  NAND2X1 U66190 ( .A(n42021), .B(n62091), .Y(n62092) );
  NAND2X1 U66191 ( .A(n62093), .B(n62092), .Y(n62095) );
  NAND2X1 U66192 ( .A(n62094), .B(n62095), .Y(n62098) );
  INVX1 U66193 ( .A(n62095), .Y(n62154) );
  NAND2X1 U66194 ( .A(n62154), .B(n62155), .Y(n62096) );
  NAND2X1 U66195 ( .A(n42035), .B(n62096), .Y(n62097) );
  NAND2X1 U66196 ( .A(n62098), .B(n62097), .Y(n62100) );
  NAND2X1 U66197 ( .A(n62099), .B(n62100), .Y(n62103) );
  INVX1 U66198 ( .A(n62100), .Y(n62151) );
  NAND2X1 U66199 ( .A(n62151), .B(n62152), .Y(n62101) );
  NAND2X1 U66200 ( .A(n42048), .B(n62101), .Y(n62102) );
  NAND2X1 U66201 ( .A(n62103), .B(n62102), .Y(n62105) );
  INVX1 U66202 ( .A(n62105), .Y(n62148) );
  NAND2X1 U66203 ( .A(n62148), .B(n62149), .Y(n62106) );
  NAND2X1 U66204 ( .A(n62146), .B(n62107), .Y(n62111) );
  INVX1 U66205 ( .A(n62146), .Y(n62108) );
  NAND2X1 U66206 ( .A(n37964), .B(n62108), .Y(n62109) );
  NAND2X1 U66207 ( .A(n42071), .B(n62109), .Y(n62110) );
  NAND2X1 U66208 ( .A(n62111), .B(n62110), .Y(n62113) );
  INVX1 U66209 ( .A(n62113), .Y(n62143) );
  NAND2X1 U66210 ( .A(n62143), .B(n62144), .Y(n62114) );
  INVX1 U66211 ( .A(n62141), .Y(n62116) );
  INVX1 U66212 ( .A(n62139), .Y(n62118) );
  NAND2X1 U66213 ( .A(n38088), .B(n38086), .Y(n62119) );
  NAND2X1 U66214 ( .A(n37970), .B(n62120), .Y(n62123) );
  NAND2X1 U66215 ( .A(n42104), .B(n62121), .Y(n62122) );
  NAND2X1 U66216 ( .A(n62123), .B(n62122), .Y(n62125) );
  NAND2X1 U66217 ( .A(n37971), .B(n62135), .Y(n62126) );
  NAND2X1 U66218 ( .A(n62133), .B(n62127), .Y(n62131) );
  INVX1 U66219 ( .A(n62133), .Y(n62128) );
  NAND2X1 U66220 ( .A(n42116), .B(n62129), .Y(n62130) );
  NAND2X1 U66221 ( .A(n62131), .B(n62130), .Y(n62570) );
  INVX1 U66222 ( .A(n62570), .Y(n62573) );
  XNOR2X1 U66223 ( .A(n62571), .B(n62573), .Y(n62132) );
  XNOR2X1 U66224 ( .A(n42119), .B(n62132), .Y(n62577) );
  INVX1 U66225 ( .A(n62577), .Y(n62329) );
  XNOR2X1 U66226 ( .A(n62133), .B(n39074), .Y(n62134) );
  XNOR2X1 U66227 ( .A(n42116), .B(n62134), .Y(n62580) );
  INVX1 U66228 ( .A(n62580), .Y(n62326) );
  XNOR2X1 U66229 ( .A(n62135), .B(n37971), .Y(n62136) );
  XNOR2X1 U66230 ( .A(n42110), .B(n62136), .Y(n62582) );
  XNOR2X1 U66231 ( .A(n62137), .B(n38090), .Y(n62138) );
  XNOR2X1 U66232 ( .A(n42104), .B(n62138), .Y(n62584) );
  XNOR2X1 U66233 ( .A(n62139), .B(n38519), .Y(n62140) );
  XNOR2X1 U66234 ( .A(n42098), .B(n62140), .Y(n62587) );
  INVX1 U66235 ( .A(n62587), .Y(n62318) );
  XNOR2X1 U66236 ( .A(n62141), .B(n38828), .Y(n62142) );
  XNOR2X1 U66237 ( .A(n42090), .B(n62142), .Y(n62589) );
  INVX1 U66238 ( .A(n62589), .Y(n62313) );
  XNOR2X1 U66239 ( .A(n62144), .B(n62143), .Y(n62145) );
  XNOR2X1 U66240 ( .A(n42080), .B(n62145), .Y(n62591) );
  XNOR2X1 U66241 ( .A(n62146), .B(n37964), .Y(n62147) );
  XNOR2X1 U66242 ( .A(n42071), .B(n62147), .Y(n62594) );
  INVX1 U66243 ( .A(n62594), .Y(n62306) );
  XNOR2X1 U66244 ( .A(n62149), .B(n62148), .Y(n62150) );
  XNOR2X1 U66245 ( .A(n42058), .B(n62150), .Y(n62596) );
  XNOR2X1 U66246 ( .A(n62152), .B(n62151), .Y(n62153) );
  XNOR2X1 U66247 ( .A(n42048), .B(n62153), .Y(n62598) );
  XNOR2X1 U66248 ( .A(n62155), .B(n62154), .Y(n62156) );
  XNOR2X1 U66249 ( .A(n42035), .B(n62156), .Y(n62600) );
  XNOR2X1 U66250 ( .A(n62158), .B(n62157), .Y(n62159) );
  XNOR2X1 U66251 ( .A(n42021), .B(n62159), .Y(n62603) );
  INVX1 U66252 ( .A(n62603), .Y(n62292) );
  XNOR2X1 U66253 ( .A(n62161), .B(n62160), .Y(n62162) );
  XNOR2X1 U66254 ( .A(n42011), .B(n62162), .Y(n62606) );
  XNOR2X1 U66255 ( .A(n62163), .B(n38063), .Y(n62164) );
  XNOR2X1 U66256 ( .A(n42000), .B(n62164), .Y(n62608) );
  XNOR2X1 U66257 ( .A(n62165), .B(n38276), .Y(n62166) );
  XNOR2X1 U66258 ( .A(n41987), .B(n62166), .Y(n62610) );
  INVX1 U66259 ( .A(n62610), .Y(n62277) );
  XNOR2X1 U66260 ( .A(n62168), .B(n62167), .Y(n62169) );
  XNOR2X1 U66261 ( .A(n41978), .B(n62169), .Y(n62613) );
  XNOR2X1 U66262 ( .A(n62171), .B(n62170), .Y(n62172) );
  XNOR2X1 U66263 ( .A(n41968), .B(n62172), .Y(n62616) );
  INVX1 U66264 ( .A(n62616), .Y(n62269) );
  XNOR2X1 U66265 ( .A(n62174), .B(n62173), .Y(n62175) );
  XNOR2X1 U66266 ( .A(n41958), .B(n62175), .Y(n62619) );
  XNOR2X1 U66267 ( .A(n62177), .B(n62176), .Y(n62178) );
  XNOR2X1 U66268 ( .A(n41949), .B(n62178), .Y(n62622) );
  INVX1 U66269 ( .A(n62622), .Y(n62259) );
  XNOR2X1 U66270 ( .A(n62179), .B(n36398), .Y(n62180) );
  XNOR2X1 U66271 ( .A(n41937), .B(n62180), .Y(n62625) );
  XNOR2X1 U66272 ( .A(n62182), .B(n62181), .Y(n62183) );
  XNOR2X1 U66273 ( .A(n41927), .B(n62183), .Y(n62628) );
  INVX1 U66274 ( .A(n62628), .Y(n62249) );
  XNOR2X1 U66275 ( .A(n62185), .B(n62184), .Y(n62186) );
  XNOR2X1 U66276 ( .A(n41917), .B(n62186), .Y(n62631) );
  XNOR2X1 U66277 ( .A(n62188), .B(n62187), .Y(n62189) );
  XNOR2X1 U66278 ( .A(n41906), .B(n62189), .Y(n62634) );
  INVX1 U66279 ( .A(n62634), .Y(n62239) );
  XNOR2X1 U66280 ( .A(n62191), .B(n62190), .Y(n62192) );
  XNOR2X1 U66281 ( .A(n41896), .B(n62192), .Y(n62637) );
  XNOR2X1 U66282 ( .A(n62194), .B(n62193), .Y(n62195) );
  XNOR2X1 U66283 ( .A(n41885), .B(n62195), .Y(n62640) );
  INVX1 U66284 ( .A(n62640), .Y(n62229) );
  XNOR2X1 U66285 ( .A(n62197), .B(n62196), .Y(n62198) );
  XNOR2X1 U66286 ( .A(n41874), .B(n62198), .Y(n62643) );
  XNOR2X1 U66287 ( .A(n62200), .B(n62199), .Y(n62201) );
  XNOR2X1 U66288 ( .A(n41864), .B(n62201), .Y(n62645) );
  INVX1 U66289 ( .A(n62645), .Y(n62219) );
  XNOR2X1 U66290 ( .A(n62202), .B(n38040), .Y(n62203) );
  XNOR2X1 U66291 ( .A(n41848), .B(n62203), .Y(n62647) );
  XNOR2X1 U66292 ( .A(n38112), .B(n62204), .Y(n62205) );
  XNOR2X1 U66293 ( .A(n62206), .B(n62205), .Y(n62649) );
  INVX1 U66294 ( .A(n62649), .Y(n62213) );
  NAND2X1 U66295 ( .A(n73384), .B(n38105), .Y(n62656) );
  INVX1 U66296 ( .A(n62657), .Y(n62651) );
  NAND2X1 U66297 ( .A(n62208), .B(n62207), .Y(n62210) );
  NAND2X1 U66298 ( .A(n62210), .B(n62209), .Y(n62652) );
  INVX1 U66299 ( .A(n62652), .Y(n62211) );
  NAND2X1 U66300 ( .A(n62657), .B(n62652), .Y(n62212) );
  NAND2X1 U66301 ( .A(n38034), .B(n62649), .Y(n62215) );
  INVX1 U66302 ( .A(n62647), .Y(n62217) );
  NAND2X1 U66303 ( .A(n36389), .B(n62217), .Y(n62218) );
  NAND2X1 U66304 ( .A(n62219), .B(n62220), .Y(n62223) );
  NAND2X1 U66305 ( .A(n36385), .B(n62645), .Y(n62221) );
  NAND2X1 U66306 ( .A(n41883), .B(n62221), .Y(n62222) );
  NAND2X1 U66307 ( .A(n62223), .B(n62222), .Y(n62224) );
  NAND2X1 U66308 ( .A(n62643), .B(n62224), .Y(n62228) );
  INVX1 U66309 ( .A(n62224), .Y(n62642) );
  INVX1 U66310 ( .A(n62643), .Y(n62225) );
  NAND2X1 U66311 ( .A(n62642), .B(n62225), .Y(n62226) );
  NAND2X1 U66312 ( .A(n41892), .B(n62226), .Y(n62227) );
  NAND2X1 U66313 ( .A(n62228), .B(n62227), .Y(n62230) );
  NAND2X1 U66314 ( .A(n62229), .B(n62230), .Y(n62233) );
  INVX1 U66315 ( .A(n62230), .Y(n62639) );
  NAND2X1 U66316 ( .A(n62639), .B(n62640), .Y(n62231) );
  NAND2X1 U66317 ( .A(n41904), .B(n62231), .Y(n62232) );
  NAND2X1 U66318 ( .A(n62233), .B(n62232), .Y(n62234) );
  NAND2X1 U66319 ( .A(n62637), .B(n62234), .Y(n62238) );
  INVX1 U66320 ( .A(n62234), .Y(n62636) );
  INVX1 U66321 ( .A(n62637), .Y(n62235) );
  NAND2X1 U66322 ( .A(n62636), .B(n62235), .Y(n62236) );
  NAND2X1 U66323 ( .A(n41915), .B(n62236), .Y(n62237) );
  NAND2X1 U66324 ( .A(n62238), .B(n62237), .Y(n62240) );
  NAND2X1 U66325 ( .A(n62239), .B(n62240), .Y(n62243) );
  INVX1 U66326 ( .A(n62240), .Y(n62633) );
  NAND2X1 U66327 ( .A(n62633), .B(n62634), .Y(n62241) );
  NAND2X1 U66328 ( .A(n41925), .B(n62241), .Y(n62242) );
  NAND2X1 U66329 ( .A(n62243), .B(n62242), .Y(n62244) );
  NAND2X1 U66330 ( .A(n62631), .B(n62244), .Y(n62248) );
  INVX1 U66331 ( .A(n62244), .Y(n62630) );
  INVX1 U66332 ( .A(n62631), .Y(n62245) );
  NAND2X1 U66333 ( .A(n62630), .B(n62245), .Y(n62246) );
  NAND2X1 U66334 ( .A(n41934), .B(n62246), .Y(n62247) );
  NAND2X1 U66335 ( .A(n62248), .B(n62247), .Y(n62250) );
  NAND2X1 U66336 ( .A(n62249), .B(n62250), .Y(n62253) );
  INVX1 U66337 ( .A(n62250), .Y(n62627) );
  NAND2X1 U66338 ( .A(n62627), .B(n62628), .Y(n62251) );
  NAND2X1 U66339 ( .A(n41946), .B(n62251), .Y(n62252) );
  NAND2X1 U66340 ( .A(n62253), .B(n62252), .Y(n62254) );
  NAND2X1 U66341 ( .A(n62625), .B(n62254), .Y(n62258) );
  INVX1 U66342 ( .A(n62254), .Y(n62624) );
  INVX1 U66343 ( .A(n62625), .Y(n62255) );
  NAND2X1 U66344 ( .A(n62624), .B(n62255), .Y(n62256) );
  NAND2X1 U66345 ( .A(n41955), .B(n62256), .Y(n62257) );
  NAND2X1 U66346 ( .A(n62258), .B(n62257), .Y(n62260) );
  NAND2X1 U66347 ( .A(n62259), .B(n62260), .Y(n62263) );
  INVX1 U66348 ( .A(n62260), .Y(n62621) );
  NAND2X1 U66349 ( .A(n62621), .B(n62622), .Y(n62261) );
  NAND2X1 U66350 ( .A(n41964), .B(n62261), .Y(n62262) );
  NAND2X1 U66351 ( .A(n62263), .B(n62262), .Y(n62264) );
  NAND2X1 U66352 ( .A(n62619), .B(n62264), .Y(n62268) );
  INVX1 U66353 ( .A(n62264), .Y(n62618) );
  INVX1 U66354 ( .A(n62619), .Y(n62265) );
  NAND2X1 U66355 ( .A(n62618), .B(n62265), .Y(n62266) );
  NAND2X1 U66356 ( .A(n41975), .B(n62266), .Y(n62267) );
  NAND2X1 U66357 ( .A(n62268), .B(n62267), .Y(n62270) );
  NAND2X1 U66358 ( .A(n62269), .B(n62270), .Y(n62273) );
  INVX1 U66359 ( .A(n62270), .Y(n62615) );
  NAND2X1 U66360 ( .A(n62615), .B(n62616), .Y(n62271) );
  NAND2X1 U66361 ( .A(n41985), .B(n62271), .Y(n62272) );
  NAND2X1 U66362 ( .A(n62273), .B(n62272), .Y(n62274) );
  INVX1 U66363 ( .A(n62274), .Y(n62612) );
  INVX1 U66364 ( .A(n62613), .Y(n62275) );
  NAND2X1 U66365 ( .A(n62612), .B(n62275), .Y(n62276) );
  NAND2X1 U66366 ( .A(n62277), .B(n62278), .Y(n62281) );
  NAND2X1 U66367 ( .A(n38237), .B(n62610), .Y(n62279) );
  NAND2X1 U66368 ( .A(n42009), .B(n62279), .Y(n62280) );
  NAND2X1 U66369 ( .A(n62281), .B(n62280), .Y(n62282) );
  NAND2X1 U66370 ( .A(n62608), .B(n62282), .Y(n62286) );
  INVX1 U66371 ( .A(n62608), .Y(n62283) );
  NAND2X1 U66372 ( .A(n38071), .B(n62283), .Y(n62284) );
  NAND2X1 U66373 ( .A(n42017), .B(n62284), .Y(n62285) );
  NAND2X1 U66374 ( .A(n62286), .B(n62285), .Y(n62287) );
  NAND2X1 U66375 ( .A(n62606), .B(n62287), .Y(n62291) );
  INVX1 U66376 ( .A(n62287), .Y(n62605) );
  INVX1 U66377 ( .A(n62606), .Y(n62288) );
  NAND2X1 U66378 ( .A(n62605), .B(n62288), .Y(n62289) );
  NAND2X1 U66379 ( .A(n42029), .B(n62289), .Y(n62290) );
  NAND2X1 U66380 ( .A(n62291), .B(n62290), .Y(n62293) );
  INVX1 U66381 ( .A(n62293), .Y(n62602) );
  NAND2X1 U66382 ( .A(n62602), .B(n62603), .Y(n62294) );
  INVX1 U66383 ( .A(n62600), .Y(n62296) );
  NAND2X1 U66384 ( .A(n36378), .B(n62296), .Y(n62297) );
  INVX1 U66385 ( .A(n62598), .Y(n62299) );
  NAND2X1 U66386 ( .A(n36364), .B(n62299), .Y(n62300) );
  NAND2X1 U66387 ( .A(n62596), .B(n62301), .Y(n62305) );
  INVX1 U66388 ( .A(n62596), .Y(n62302) );
  NAND2X1 U66389 ( .A(n36367), .B(n62302), .Y(n62303) );
  NAND2X1 U66390 ( .A(n42077), .B(n62303), .Y(n62304) );
  NAND2X1 U66391 ( .A(n62305), .B(n62304), .Y(n62307) );
  INVX1 U66392 ( .A(n62307), .Y(n62593) );
  NAND2X1 U66393 ( .A(n62593), .B(n62594), .Y(n62308) );
  NAND2X1 U66394 ( .A(n62591), .B(n37923), .Y(n62312) );
  INVX1 U66395 ( .A(n62591), .Y(n62309) );
  NAND2X1 U66396 ( .A(n38037), .B(n62309), .Y(n62310) );
  NAND2X1 U66397 ( .A(n42096), .B(n62310), .Y(n62311) );
  NAND2X1 U66398 ( .A(n62312), .B(n62311), .Y(n62314) );
  NAND2X1 U66399 ( .A(n62313), .B(n62314), .Y(n62317) );
  NAND2X1 U66400 ( .A(n38027), .B(n62589), .Y(n62315) );
  NAND2X1 U66401 ( .A(n42102), .B(n62315), .Y(n62316) );
  NAND2X1 U66402 ( .A(n62317), .B(n62316), .Y(n62319) );
  INVX1 U66403 ( .A(n62319), .Y(n62586) );
  NAND2X1 U66404 ( .A(n62586), .B(n62587), .Y(n62320) );
  INVX1 U66405 ( .A(n62584), .Y(n62321) );
  NAND2X1 U66406 ( .A(n38754), .B(n62321), .Y(n62322) );
  NAND2X1 U66407 ( .A(n62582), .B(n38081), .Y(n62325) );
  INVX1 U66408 ( .A(n62582), .Y(n62323) );
  NAND2X1 U66409 ( .A(n62325), .B(n62324), .Y(n62327) );
  NAND2X1 U66410 ( .A(n37924), .B(n62580), .Y(n62328) );
  NAND2X1 U66411 ( .A(n62329), .B(n38776), .Y(n62332) );
  NAND2X1 U66412 ( .A(n38906), .B(n62577), .Y(n62330) );
  NAND2X1 U66413 ( .A(n42128), .B(n62330), .Y(n62331) );
  AND2X1 U66414 ( .A(n62332), .B(n62331), .Y(n62808) );
  INVX1 U66415 ( .A(n62335), .Y(n62334) );
  NAND2X1 U66416 ( .A(n37951), .B(n62335), .Y(n62336) );
  INVX1 U66417 ( .A(n62338), .Y(n62337) );
  NAND2X1 U66418 ( .A(n38498), .B(n38497), .Y(n62339) );
  NAND2X1 U66419 ( .A(n62344), .B(n62342), .Y(n62351) );
  INVX1 U66420 ( .A(n62343), .Y(n62349) );
  XNOR2X1 U66421 ( .A(n62364), .B(n62345), .Y(n62347) );
  INVX1 U66422 ( .A(n62363), .Y(n62346) );
  NAND2X1 U66423 ( .A(n62349), .B(n62348), .Y(n62350) );
  NAND2X1 U66424 ( .A(n62351), .B(n62350), .Y(n62827) );
  XNOR2X1 U66425 ( .A(n63032), .B(n38598), .Y(n62352) );
  NOR2X1 U66426 ( .A(n62353), .B(n62355), .Y(n62362) );
  OR2X1 U66427 ( .A(n62355), .B(n62354), .Y(n62360) );
  NOR2X1 U66428 ( .A(n62356), .B(n62355), .Y(n62358) );
  NAND2X1 U66429 ( .A(n62358), .B(n62357), .Y(n62359) );
  NAND2X1 U66430 ( .A(n62360), .B(n62359), .Y(n62361) );
  NOR2X1 U66431 ( .A(n62362), .B(n62361), .Y(n62366) );
  NAND2X1 U66432 ( .A(n62364), .B(n62363), .Y(n62365) );
  INVX1 U66433 ( .A(n62367), .Y(n62370) );
  NAND2X1 U66434 ( .A(n39522), .B(n62368), .Y(n62369) );
  NAND2X1 U66435 ( .A(n62370), .B(n62369), .Y(n62374) );
  NAND2X1 U66436 ( .A(n62372), .B(n62371), .Y(n62373) );
  NAND2X1 U66437 ( .A(n62374), .B(n62373), .Y(n63029) );
  NAND2X1 U66438 ( .A(n72820), .B(n43944), .Y(n63372) );
  INVX1 U66439 ( .A(n38676), .Y(n62375) );
  NAND2X1 U66440 ( .A(n38676), .B(n62378), .Y(n62379) );
  NAND2X1 U66441 ( .A(n38912), .B(n38450), .Y(n62862) );
  INVX1 U66442 ( .A(n62383), .Y(n62381) );
  NAND2X1 U66443 ( .A(n39215), .B(n62384), .Y(n62385) );
  NAND2X1 U66444 ( .A(n62386), .B(n62385), .Y(n62388) );
  NAND2X1 U66445 ( .A(n62388), .B(n62387), .Y(n62389) );
  INVX1 U66446 ( .A(n63019), .Y(n63353) );
  NAND2X1 U66447 ( .A(n43896), .B(n42639), .Y(n63355) );
  NAND2X1 U66448 ( .A(n40259), .B(n43890), .Y(n63345) );
  INVX1 U66449 ( .A(n62404), .Y(n63008) );
  NOR2X1 U66450 ( .A(n62396), .B(n62393), .Y(n62394) );
  NOR2X1 U66451 ( .A(n62395), .B(n62394), .Y(n62400) );
  INVX1 U66452 ( .A(n62396), .Y(n62398) );
  NAND2X1 U66453 ( .A(n62398), .B(n62397), .Y(n62399) );
  NAND2X1 U66454 ( .A(n62400), .B(n62399), .Y(n62868) );
  XNOR2X1 U66455 ( .A(n63345), .B(n39563), .Y(n62510) );
  NAND2X1 U66456 ( .A(n43798), .B(n43880), .Y(n63014) );
  INVX1 U66457 ( .A(n62420), .Y(n62417) );
  XNOR2X1 U66458 ( .A(n41253), .B(n62417), .Y(n62401) );
  XNOR2X1 U66459 ( .A(n62401), .B(n39344), .Y(n62402) );
  XNOR2X1 U66460 ( .A(n37388), .B(n62402), .Y(n62403) );
  INVX1 U66461 ( .A(n62403), .Y(n63010) );
  NOR2X1 U66462 ( .A(n63008), .B(n63010), .Y(n62408) );
  NAND2X1 U66463 ( .A(n62405), .B(n62403), .Y(n63007) );
  NAND2X1 U66464 ( .A(n62405), .B(n62404), .Y(n62406) );
  NAND2X1 U66465 ( .A(n63007), .B(n62406), .Y(n62407) );
  XNOR2X1 U66466 ( .A(n39344), .B(n62409), .Y(n62410) );
  XNOR2X1 U66467 ( .A(n62410), .B(n62417), .Y(n62415) );
  NOR2X1 U66468 ( .A(n39275), .B(n41506), .Y(n62413) );
  NAND2X1 U66469 ( .A(n62413), .B(n62412), .Y(n62414) );
  NAND2X1 U66470 ( .A(n62415), .B(n62414), .Y(n62997) );
  NAND2X1 U66471 ( .A(n62998), .B(n62997), .Y(n63322) );
  NOR2X1 U66472 ( .A(n38638), .B(n62416), .Y(n62419) );
  NOR2X1 U66473 ( .A(n62417), .B(n62416), .Y(n62418) );
  NOR2X1 U66474 ( .A(n62418), .B(n62419), .Y(n62422) );
  NAND2X1 U66475 ( .A(n62420), .B(n38655), .Y(n62421) );
  NAND2X1 U66476 ( .A(n62422), .B(n62421), .Y(n62870) );
  NAND2X1 U66477 ( .A(n43962), .B(n43796), .Y(n62874) );
  NAND2X1 U66478 ( .A(n43860), .B(n43776), .Y(n63305) );
  NAND2X1 U66479 ( .A(n43850), .B(n43479), .Y(n63290) );
  NAND2X1 U66480 ( .A(n62426), .B(n62425), .Y(n62429) );
  INVX1 U66481 ( .A(n62427), .Y(n62430) );
  NOR2X1 U66482 ( .A(n40024), .B(n62431), .Y(n62487) );
  INVX1 U66483 ( .A(n62433), .Y(n62435) );
  NAND2X1 U66484 ( .A(n62435), .B(n62434), .Y(n62436) );
  NAND2X1 U66485 ( .A(n62437), .B(n62436), .Y(n62962) );
  NAND2X1 U66486 ( .A(n39943), .B(n43496), .Y(n63253) );
  INVX1 U66487 ( .A(n62440), .Y(n62438) );
  NAND2X1 U66488 ( .A(n62438), .B(n62439), .Y(n62943) );
  INVX1 U66489 ( .A(n62439), .Y(n62441) );
  NAND2X1 U66490 ( .A(n62943), .B(n62945), .Y(n62938) );
  NAND2X1 U66491 ( .A(n61191), .B(n42153), .Y(n63183) );
  NAND2X1 U66492 ( .A(n63830), .B(n63183), .Y(n62451) );
  INVX1 U66493 ( .A(n64087), .Y(n72336) );
  NAND2X1 U66494 ( .A(n43603), .B(n62903), .Y(n62444) );
  NOR2X1 U66495 ( .A(n43454), .B(n62444), .Y(n62446) );
  NOR2X1 U66496 ( .A(n64087), .B(n62909), .Y(n62445) );
  NOR2X1 U66497 ( .A(n62446), .B(n62445), .Y(n62450) );
  NAND2X1 U66498 ( .A(n62907), .B(n62905), .Y(n62447) );
  NOR2X1 U66499 ( .A(n64087), .B(n62447), .Y(n62448) );
  NAND2X1 U66500 ( .A(n62448), .B(n62453), .Y(n62449) );
  NAND2X1 U66501 ( .A(n62450), .B(n62449), .Y(n63208) );
  NAND2X1 U66502 ( .A(n63208), .B(n63183), .Y(n63193) );
  XNOR2X1 U66503 ( .A(n62451), .B(n63193), .Y(n63556) );
  NOR2X1 U66504 ( .A(n63823), .B(n63822), .Y(n62452) );
  INVX1 U66505 ( .A(n62453), .Y(n62454) );
  NOR2X1 U66506 ( .A(n62454), .B(n42799), .Y(n62456) );
  NOR2X1 U66507 ( .A(n62456), .B(n62455), .Y(n62457) );
  NOR2X1 U66508 ( .A(n62458), .B(n62457), .Y(n62459) );
  NAND2X1 U66509 ( .A(n63827), .B(n62459), .Y(n62464) );
  INVX1 U66510 ( .A(n62460), .Y(n62461) );
  NOR2X1 U66511 ( .A(n62461), .B(n63190), .Y(n62462) );
  NOR2X1 U66512 ( .A(n38235), .B(n62462), .Y(n62463) );
  XNOR2X1 U66513 ( .A(n41770), .B(n38691), .Y(n62467) );
  INVX1 U66514 ( .A(n62465), .Y(n62466) );
  NAND2X1 U66515 ( .A(n39641), .B(n63555), .Y(n62939) );
  XNOR2X1 U66516 ( .A(n62467), .B(n39621), .Y(n62468) );
  XNOR2X1 U66517 ( .A(n63253), .B(n37373), .Y(n62477) );
  NOR2X1 U66518 ( .A(n40086), .B(n62469), .Y(n62472) );
  INVX1 U66519 ( .A(n62473), .Y(n62470) );
  NOR2X1 U66520 ( .A(n62470), .B(n62469), .Y(n62471) );
  NOR2X1 U66521 ( .A(n62472), .B(n62471), .Y(n62476) );
  NAND2X1 U66522 ( .A(n62474), .B(n62473), .Y(n62475) );
  NAND2X1 U66523 ( .A(n62476), .B(n62475), .Y(n62951) );
  INVX1 U66524 ( .A(n62951), .Y(n62950) );
  XNOR2X1 U66525 ( .A(n62477), .B(n62950), .Y(n62963) );
  NAND2X1 U66526 ( .A(n43493), .B(n43842), .Y(n62958) );
  XNOR2X1 U66527 ( .A(n62963), .B(n62958), .Y(n62478) );
  XNOR2X1 U66528 ( .A(n62962), .B(n62478), .Y(n62977) );
  NAND2X1 U66529 ( .A(n44035), .B(n43482), .Y(n63274) );
  INVX1 U66530 ( .A(n63274), .Y(n63279) );
  NAND2X1 U66531 ( .A(n38382), .B(n38310), .Y(n62978) );
  INVX1 U66532 ( .A(n62978), .Y(n62968) );
  XNOR2X1 U66533 ( .A(n63279), .B(n62968), .Y(n62484) );
  INVX1 U66534 ( .A(n62479), .Y(n62482) );
  NAND2X1 U66535 ( .A(n62482), .B(n62481), .Y(n62973) );
  NAND2X1 U66536 ( .A(n62973), .B(n62972), .Y(n62483) );
  NOR2X1 U66537 ( .A(n39723), .B(n62483), .Y(n62964) );
  XNOR2X1 U66538 ( .A(n62484), .B(n62964), .Y(n62485) );
  XNOR2X1 U66539 ( .A(n62977), .B(n62485), .Y(n62486) );
  XNOR2X1 U66540 ( .A(n62487), .B(n62486), .Y(n62885) );
  INVX1 U66541 ( .A(n62885), .Y(n63291) );
  INVX1 U66542 ( .A(n62488), .Y(n62489) );
  NAND2X1 U66543 ( .A(n62491), .B(n62490), .Y(n62883) );
  INVX1 U66544 ( .A(n63306), .Y(n62881) );
  NAND2X1 U66545 ( .A(n62493), .B(n62494), .Y(n62877) );
  INVX1 U66546 ( .A(n62877), .Y(n62497) );
  INVX1 U66547 ( .A(n62492), .Y(n62495) );
  NAND2X1 U66548 ( .A(n62495), .B(n62493), .Y(n62878) );
  NAND2X1 U66549 ( .A(n62495), .B(n62494), .Y(n62879) );
  NAND2X1 U66550 ( .A(n62878), .B(n62879), .Y(n62496) );
  NOR2X1 U66551 ( .A(n62497), .B(n62496), .Y(n62498) );
  XNOR2X1 U66552 ( .A(n62874), .B(n38257), .Y(n62506) );
  NOR2X1 U66553 ( .A(n40082), .B(n62499), .Y(n62502) );
  NOR2X1 U66554 ( .A(n62500), .B(n62499), .Y(n62501) );
  NOR2X1 U66555 ( .A(n62502), .B(n62501), .Y(n62505) );
  NAND2X1 U66556 ( .A(n39709), .B(n62503), .Y(n62504) );
  NAND2X1 U66557 ( .A(n62505), .B(n62504), .Y(n62873) );
  XNOR2X1 U66558 ( .A(n62506), .B(n38397), .Y(n62871) );
  NAND2X1 U66559 ( .A(n43953), .B(n42714), .Y(n63156) );
  XNOR2X1 U66560 ( .A(n62871), .B(n63156), .Y(n62507) );
  XNOR2X1 U66561 ( .A(n62870), .B(n62507), .Y(n63324) );
  NAND2X1 U66562 ( .A(n42661), .B(n43871), .Y(n63320) );
  XNOR2X1 U66563 ( .A(n63324), .B(n63320), .Y(n62508) );
  XNOR2X1 U66564 ( .A(n63322), .B(n62508), .Y(n63015) );
  INVX1 U66565 ( .A(n63015), .Y(n63013) );
  XNOR2X1 U66566 ( .A(n62509), .B(n63013), .Y(n62869) );
  INVX1 U66567 ( .A(n62869), .Y(n63347) );
  XNOR2X1 U66568 ( .A(n62510), .B(n63347), .Y(n63020) );
  INVX1 U66569 ( .A(n63020), .Y(n63356) );
  INVX1 U66570 ( .A(n62864), .Y(n62867) );
  NAND2X1 U66571 ( .A(n43724), .B(n43904), .Y(n62863) );
  NOR2X1 U66572 ( .A(n62514), .B(n62511), .Y(n62512) );
  INVX1 U66573 ( .A(n62514), .Y(n62516) );
  XNOR2X1 U66574 ( .A(n62863), .B(n39765), .Y(n62517) );
  XNOR2X1 U66575 ( .A(n62867), .B(n62517), .Y(n63141) );
  NAND2X1 U66576 ( .A(n43910), .B(n43788), .Y(n63140) );
  INVX1 U66577 ( .A(n63140), .Y(n62860) );
  XNOR2X1 U66578 ( .A(n63141), .B(n62860), .Y(n62518) );
  XNOR2X1 U66579 ( .A(n40452), .B(n62518), .Y(n62855) );
  INVX1 U66580 ( .A(n62855), .Y(n62858) );
  NAND2X1 U66581 ( .A(n62520), .B(n62519), .Y(n62521) );
  NAND2X1 U66582 ( .A(n62521), .B(n62850), .Y(n62851) );
  INVX1 U66583 ( .A(n62851), .Y(n62523) );
  INVX1 U66584 ( .A(n62521), .Y(n62849) );
  NAND2X1 U66585 ( .A(n38479), .B(n62850), .Y(n62524) );
  XNOR2X1 U66586 ( .A(n62859), .B(n41966), .Y(n62525) );
  XNOR2X1 U66587 ( .A(n62858), .B(n62525), .Y(n62847) );
  INVX1 U66588 ( .A(n62847), .Y(n62842) );
  NAND2X1 U66589 ( .A(n43927), .B(n40471), .Y(n62846) );
  NAND2X1 U66590 ( .A(n62526), .B(n39417), .Y(n62532) );
  INVX1 U66591 ( .A(n62527), .Y(n62530) );
  NAND2X1 U66592 ( .A(n62530), .B(n62529), .Y(n62531) );
  AND2X1 U66593 ( .A(n62532), .B(n62531), .Y(n62843) );
  XNOR2X1 U66594 ( .A(n62846), .B(n62843), .Y(n62533) );
  XNOR2X1 U66595 ( .A(n62842), .B(n62533), .Y(n62839) );
  INVX1 U66596 ( .A(n62839), .Y(n62541) );
  NAND2X1 U66597 ( .A(n40461), .B(n43935), .Y(n62838) );
  INVX1 U66598 ( .A(n62537), .Y(n62539) );
  XNOR2X1 U66599 ( .A(n62838), .B(n41268), .Y(n62540) );
  XNOR2X1 U66600 ( .A(n62541), .B(n62540), .Y(n63371) );
  INVX1 U66601 ( .A(n63371), .Y(n63028) );
  NAND2X1 U66602 ( .A(n43820), .B(n43974), .Y(n63121) );
  INVX1 U66603 ( .A(n63121), .Y(n63041) );
  NOR2X1 U66604 ( .A(n63041), .B(n63034), .Y(n62543) );
  NAND2X1 U66605 ( .A(n43947), .B(n63121), .Y(n62542) );
  NAND2X1 U66606 ( .A(n62542), .B(n43821), .Y(n62547) );
  NOR2X1 U66607 ( .A(n62543), .B(n62547), .Y(n62544) );
  NOR2X1 U66608 ( .A(n62544), .B(n40279), .Y(n62554) );
  NAND2X1 U66609 ( .A(n63041), .B(n63034), .Y(n62545) );
  NAND2X1 U66610 ( .A(n63041), .B(n43944), .Y(n62548) );
  NAND2X1 U66611 ( .A(n62545), .B(n62548), .Y(n62546) );
  NAND2X1 U66612 ( .A(n62546), .B(n40280), .Y(n62552) );
  OR2X1 U66613 ( .A(n38598), .B(n62547), .Y(n62550) );
  NAND2X1 U66614 ( .A(n62548), .B(n38598), .Y(n62549) );
  NAND2X1 U66615 ( .A(n62550), .B(n62549), .Y(n62551) );
  NAND2X1 U66616 ( .A(n62552), .B(n62551), .Y(n62553) );
  NOR2X1 U66617 ( .A(n62554), .B(n62553), .Y(n62555) );
  XOR2X1 U66618 ( .A(n63036), .B(n62555), .Y(n62832) );
  INVX1 U66619 ( .A(n62832), .Y(n62831) );
  XNOR2X1 U66620 ( .A(n38164), .B(n62831), .Y(n62556) );
  XNOR2X1 U66621 ( .A(n42028), .B(n62556), .Y(n62828) );
  NAND2X1 U66622 ( .A(n43735), .B(n43993), .Y(n62829) );
  XNOR2X1 U66623 ( .A(n62828), .B(n62829), .Y(n62557) );
  INVX1 U66624 ( .A(n62559), .Y(n62558) );
  NAND2X1 U66625 ( .A(n62558), .B(n36513), .Y(n63047) );
  NAND2X1 U66626 ( .A(n63047), .B(n63048), .Y(n63046) );
  XNOR2X1 U66627 ( .A(n63046), .B(n42062), .Y(n62560) );
  XNOR2X1 U66628 ( .A(n36782), .B(n62560), .Y(n62823) );
  INVX1 U66629 ( .A(n62823), .Y(n62825) );
  XNOR2X1 U66630 ( .A(n62824), .B(n62825), .Y(n62561) );
  XNOR2X1 U66631 ( .A(n42075), .B(n62561), .Y(n63055) );
  INVX1 U66632 ( .A(n63055), .Y(n63053) );
  XNOR2X1 U66633 ( .A(n63054), .B(n63053), .Y(n62562) );
  XNOR2X1 U66634 ( .A(n42093), .B(n62562), .Y(n62818) );
  NAND2X1 U66635 ( .A(n62564), .B(n62563), .Y(n62567) );
  INVX1 U66636 ( .A(n62564), .Y(n62565) );
  NAND2X1 U66637 ( .A(n62567), .B(n62566), .Y(n62817) );
  INVX1 U66638 ( .A(n62817), .Y(n62819) );
  XNOR2X1 U66639 ( .A(n62818), .B(n62819), .Y(n62568) );
  XNOR2X1 U66640 ( .A(n42101), .B(n62568), .Y(n63061) );
  INVX1 U66641 ( .A(n63061), .Y(n63059) );
  XNOR2X1 U66642 ( .A(n63060), .B(n63059), .Y(n62569) );
  XNOR2X1 U66643 ( .A(n42117), .B(n62569), .Y(n62812) );
  INVX1 U66644 ( .A(n62571), .Y(n62572) );
  NAND2X1 U66645 ( .A(n62573), .B(n62572), .Y(n62574) );
  XNOR2X1 U66646 ( .A(n62812), .B(n39302), .Y(n62575) );
  XNOR2X1 U66647 ( .A(n42126), .B(n62575), .Y(n62805) );
  NAND2X1 U66648 ( .A(n43612), .B(n43752), .Y(n72698) );
  XNOR2X1 U66649 ( .A(n62805), .B(n43692), .Y(n62576) );
  XNOR2X1 U66650 ( .A(n62808), .B(n62576), .Y(n63068) );
  INVX1 U66651 ( .A(n63068), .Y(n63067) );
  XNOR2X1 U66652 ( .A(n43709), .B(n63067), .Y(n62800) );
  XNOR2X1 U66653 ( .A(n62577), .B(n38906), .Y(n62578) );
  XNOR2X1 U66654 ( .A(n42128), .B(n62578), .Y(n62579) );
  NAND2X1 U66655 ( .A(n43706), .B(n62579), .Y(n62799) );
  INVX1 U66656 ( .A(n62579), .Y(n72729) );
  NAND2X1 U66657 ( .A(n72729), .B(n72708), .Y(n62797) );
  XNOR2X1 U66658 ( .A(n62580), .B(n37924), .Y(n62581) );
  XNOR2X1 U66659 ( .A(n42124), .B(n62581), .Y(n62795) );
  XNOR2X1 U66660 ( .A(n62582), .B(n38419), .Y(n62583) );
  XNOR2X1 U66661 ( .A(n42118), .B(n62583), .Y(n72112) );
  INVX1 U66662 ( .A(n72112), .Y(n62789) );
  XNOR2X1 U66663 ( .A(n62584), .B(n38754), .Y(n62585) );
  XNOR2X1 U66664 ( .A(n42114), .B(n62585), .Y(n71718) );
  INVX1 U66665 ( .A(n71718), .Y(n62786) );
  XNOR2X1 U66666 ( .A(n62587), .B(n62586), .Y(n62588) );
  XNOR2X1 U66667 ( .A(n42108), .B(n62588), .Y(n71408) );
  XNOR2X1 U66668 ( .A(n62589), .B(n38027), .Y(n62590) );
  XNOR2X1 U66669 ( .A(n42102), .B(n62590), .Y(n62778) );
  XNOR2X1 U66670 ( .A(n62591), .B(n38037), .Y(n62592) );
  XNOR2X1 U66671 ( .A(n42096), .B(n62592), .Y(n70798) );
  INVX1 U66672 ( .A(n70798), .Y(n62775) );
  XNOR2X1 U66673 ( .A(n62594), .B(n62593), .Y(n62595) );
  XNOR2X1 U66674 ( .A(n42087), .B(n62595), .Y(n62771) );
  XNOR2X1 U66675 ( .A(n62596), .B(n36367), .Y(n62597) );
  XNOR2X1 U66676 ( .A(n42077), .B(n62597), .Y(n70195) );
  INVX1 U66677 ( .A(n70195), .Y(n62765) );
  XNOR2X1 U66678 ( .A(n62598), .B(n36364), .Y(n62599) );
  XNOR2X1 U66679 ( .A(n42066), .B(n62599), .Y(n69907) );
  INVX1 U66680 ( .A(n69907), .Y(n62760) );
  XNOR2X1 U66681 ( .A(n62600), .B(n36378), .Y(n62601) );
  XNOR2X1 U66682 ( .A(n42055), .B(n62601), .Y(n69566) );
  INVX1 U66683 ( .A(n69566), .Y(n62756) );
  XNOR2X1 U66684 ( .A(n62603), .B(n62602), .Y(n62604) );
  XNOR2X1 U66685 ( .A(n42041), .B(n62604), .Y(n62752) );
  XNOR2X1 U66686 ( .A(n62606), .B(n62605), .Y(n62607) );
  XNOR2X1 U66687 ( .A(n42029), .B(n62607), .Y(n68850) );
  INVX1 U66688 ( .A(n68850), .Y(n62746) );
  XNOR2X1 U66689 ( .A(n62608), .B(n38071), .Y(n62609) );
  XNOR2X1 U66690 ( .A(n42017), .B(n62609), .Y(n68533) );
  INVX1 U66691 ( .A(n68533), .Y(n62741) );
  XNOR2X1 U66692 ( .A(n62610), .B(n38070), .Y(n62611) );
  XNOR2X1 U66693 ( .A(n42009), .B(n62611), .Y(n62737) );
  XNOR2X1 U66694 ( .A(n62613), .B(n62612), .Y(n62614) );
  XNOR2X1 U66695 ( .A(n41996), .B(n62614), .Y(n67906) );
  INVX1 U66696 ( .A(n67906), .Y(n62732) );
  XNOR2X1 U66697 ( .A(n62616), .B(n62615), .Y(n62617) );
  XNOR2X1 U66698 ( .A(n41985), .B(n62617), .Y(n62728) );
  XNOR2X1 U66699 ( .A(n62619), .B(n62618), .Y(n62620) );
  XNOR2X1 U66700 ( .A(n41975), .B(n62620), .Y(n67240) );
  INVX1 U66701 ( .A(n67240), .Y(n62722) );
  XNOR2X1 U66702 ( .A(n62622), .B(n62621), .Y(n62623) );
  XNOR2X1 U66703 ( .A(n41964), .B(n62623), .Y(n62718) );
  XNOR2X1 U66704 ( .A(n62625), .B(n62624), .Y(n62626) );
  XNOR2X1 U66705 ( .A(n41955), .B(n62626), .Y(n66558) );
  INVX1 U66706 ( .A(n66558), .Y(n62712) );
  XNOR2X1 U66707 ( .A(n62628), .B(n62627), .Y(n62629) );
  XNOR2X1 U66708 ( .A(n41946), .B(n62629), .Y(n62708) );
  XNOR2X1 U66709 ( .A(n62631), .B(n62630), .Y(n62632) );
  XNOR2X1 U66710 ( .A(n41934), .B(n62632), .Y(n65940) );
  INVX1 U66711 ( .A(n65940), .Y(n62703) );
  XNOR2X1 U66712 ( .A(n62634), .B(n62633), .Y(n62635) );
  XNOR2X1 U66713 ( .A(n41925), .B(n62635), .Y(n62701) );
  XNOR2X1 U66714 ( .A(n62637), .B(n62636), .Y(n62638) );
  XNOR2X1 U66715 ( .A(n41915), .B(n62638), .Y(n65214) );
  INVX1 U66716 ( .A(n65214), .Y(n62695) );
  XNOR2X1 U66717 ( .A(n62640), .B(n62639), .Y(n62641) );
  XNOR2X1 U66718 ( .A(n41904), .B(n62641), .Y(n62691) );
  XNOR2X1 U66719 ( .A(n62643), .B(n62642), .Y(n62644) );
  XNOR2X1 U66720 ( .A(n41892), .B(n62644), .Y(n64569) );
  INVX1 U66721 ( .A(n64569), .Y(n62685) );
  XNOR2X1 U66722 ( .A(n62645), .B(n36385), .Y(n62646) );
  XNOR2X1 U66723 ( .A(n41883), .B(n62646), .Y(n62681) );
  XNOR2X1 U66724 ( .A(n62647), .B(n36389), .Y(n62648) );
  XNOR2X1 U66725 ( .A(n41872), .B(n62648), .Y(n63958) );
  INVX1 U66726 ( .A(n63958), .Y(n62675) );
  XNOR2X1 U66727 ( .A(n62649), .B(n38034), .Y(n62650) );
  XNOR2X1 U66728 ( .A(n41860), .B(n62650), .Y(n62671) );
  XNOR2X1 U66729 ( .A(n62652), .B(n62651), .Y(n62653) );
  XNOR2X1 U66730 ( .A(n41846), .B(n62653), .Y(n63398) );
  INVX1 U66731 ( .A(n63398), .Y(n62665) );
  NOR2X1 U66732 ( .A(n62458), .B(n62655), .Y(n62654) );
  NAND2X1 U66733 ( .A(n62654), .B(n43731), .Y(n62660) );
  INVX1 U66734 ( .A(n62660), .Y(n63073) );
  NAND2X1 U66735 ( .A(n62656), .B(n62655), .Y(n62658) );
  NAND2X1 U66736 ( .A(n62658), .B(n62657), .Y(n62661) );
  INVX1 U66737 ( .A(n62661), .Y(n63074) );
  NAND2X1 U66738 ( .A(n63073), .B(n63074), .Y(n62664) );
  NAND2X1 U66739 ( .A(n62661), .B(n62660), .Y(n62662) );
  NAND2X1 U66740 ( .A(n41866), .B(n62662), .Y(n62663) );
  NAND2X1 U66741 ( .A(n62664), .B(n62663), .Y(n62666) );
  NAND2X1 U66742 ( .A(n62665), .B(n62666), .Y(n62669) );
  INVX1 U66743 ( .A(n62666), .Y(n63397) );
  NAND2X1 U66744 ( .A(n63397), .B(n63398), .Y(n62667) );
  NAND2X1 U66745 ( .A(n41876), .B(n62667), .Y(n62668) );
  NAND2X1 U66746 ( .A(n62669), .B(n62668), .Y(n62670) );
  NAND2X1 U66747 ( .A(n62671), .B(n62670), .Y(n62674) );
  INVX1 U66748 ( .A(n62670), .Y(n63692) );
  INVX1 U66749 ( .A(n62671), .Y(n63691) );
  NAND2X1 U66750 ( .A(n63692), .B(n63691), .Y(n62672) );
  NAND2X1 U66751 ( .A(n41887), .B(n62672), .Y(n62673) );
  NAND2X1 U66752 ( .A(n62674), .B(n62673), .Y(n62676) );
  NAND2X1 U66753 ( .A(n62675), .B(n62676), .Y(n62679) );
  INVX1 U66754 ( .A(n62676), .Y(n63957) );
  NAND2X1 U66755 ( .A(n63957), .B(n63958), .Y(n62677) );
  NAND2X1 U66756 ( .A(n41898), .B(n62677), .Y(n62678) );
  NAND2X1 U66757 ( .A(n62679), .B(n62678), .Y(n62680) );
  NAND2X1 U66758 ( .A(n62681), .B(n62680), .Y(n62684) );
  INVX1 U66759 ( .A(n62680), .Y(n64283) );
  INVX1 U66760 ( .A(n62681), .Y(n64282) );
  NAND2X1 U66761 ( .A(n64283), .B(n64282), .Y(n62682) );
  NAND2X1 U66762 ( .A(n41908), .B(n62682), .Y(n62683) );
  NAND2X1 U66763 ( .A(n62684), .B(n62683), .Y(n62686) );
  NAND2X1 U66764 ( .A(n62685), .B(n62686), .Y(n62689) );
  INVX1 U66765 ( .A(n62686), .Y(n64568) );
  NAND2X1 U66766 ( .A(n64568), .B(n64569), .Y(n62687) );
  NAND2X1 U66767 ( .A(n41918), .B(n62687), .Y(n62688) );
  NAND2X1 U66768 ( .A(n62689), .B(n62688), .Y(n62690) );
  NAND2X1 U66769 ( .A(n62691), .B(n62690), .Y(n62694) );
  INVX1 U66770 ( .A(n62690), .Y(n64898) );
  INVX1 U66771 ( .A(n62691), .Y(n64897) );
  NAND2X1 U66772 ( .A(n64898), .B(n64897), .Y(n62692) );
  NAND2X1 U66773 ( .A(n41928), .B(n62692), .Y(n62693) );
  NAND2X1 U66774 ( .A(n62694), .B(n62693), .Y(n62696) );
  NAND2X1 U66775 ( .A(n62695), .B(n62696), .Y(n62699) );
  INVX1 U66776 ( .A(n62696), .Y(n65213) );
  NAND2X1 U66777 ( .A(n65213), .B(n65214), .Y(n62697) );
  NAND2X1 U66778 ( .A(n41940), .B(n62697), .Y(n62698) );
  NAND2X1 U66779 ( .A(n62699), .B(n62698), .Y(n62700) );
  INVX1 U66780 ( .A(n62700), .Y(n65576) );
  INVX1 U66781 ( .A(n62701), .Y(n65575) );
  NAND2X1 U66782 ( .A(n65576), .B(n65575), .Y(n62702) );
  NAND2X1 U66783 ( .A(n62703), .B(n65941), .Y(n62706) );
  NAND2X1 U66784 ( .A(n36358), .B(n65940), .Y(n62704) );
  NAND2X1 U66785 ( .A(n41959), .B(n62704), .Y(n62705) );
  NAND2X1 U66786 ( .A(n62706), .B(n62705), .Y(n62707) );
  NAND2X1 U66787 ( .A(n62708), .B(n62707), .Y(n62711) );
  INVX1 U66788 ( .A(n62707), .Y(n66246) );
  INVX1 U66789 ( .A(n62708), .Y(n66245) );
  NAND2X1 U66790 ( .A(n66246), .B(n66245), .Y(n62709) );
  NAND2X1 U66791 ( .A(n41969), .B(n62709), .Y(n62710) );
  NAND2X1 U66792 ( .A(n62711), .B(n62710), .Y(n62713) );
  NAND2X1 U66793 ( .A(n62712), .B(n62713), .Y(n62716) );
  INVX1 U66794 ( .A(n62713), .Y(n66557) );
  NAND2X1 U66795 ( .A(n66557), .B(n66558), .Y(n62714) );
  NAND2X1 U66796 ( .A(n41979), .B(n62714), .Y(n62715) );
  NAND2X1 U66797 ( .A(n62716), .B(n62715), .Y(n62717) );
  NAND2X1 U66798 ( .A(n62718), .B(n62717), .Y(n62721) );
  INVX1 U66799 ( .A(n62717), .Y(n66909) );
  INVX1 U66800 ( .A(n62718), .Y(n66908) );
  NAND2X1 U66801 ( .A(n66909), .B(n66908), .Y(n62719) );
  NAND2X1 U66802 ( .A(n41988), .B(n62719), .Y(n62720) );
  NAND2X1 U66803 ( .A(n62721), .B(n62720), .Y(n62723) );
  NAND2X1 U66804 ( .A(n62722), .B(n62723), .Y(n62726) );
  INVX1 U66805 ( .A(n62723), .Y(n67239) );
  NAND2X1 U66806 ( .A(n67239), .B(n67240), .Y(n62724) );
  NAND2X1 U66807 ( .A(n42001), .B(n62724), .Y(n62725) );
  NAND2X1 U66808 ( .A(n62726), .B(n62725), .Y(n62727) );
  NAND2X1 U66809 ( .A(n62728), .B(n62727), .Y(n62731) );
  INVX1 U66810 ( .A(n62727), .Y(n67601) );
  INVX1 U66811 ( .A(n62728), .Y(n67600) );
  NAND2X1 U66812 ( .A(n67601), .B(n67600), .Y(n62729) );
  NAND2X1 U66813 ( .A(n42012), .B(n62729), .Y(n62730) );
  NAND2X1 U66814 ( .A(n62731), .B(n62730), .Y(n67907) );
  NAND2X1 U66815 ( .A(n62732), .B(n67907), .Y(n62735) );
  NAND2X1 U66816 ( .A(n37903), .B(n67906), .Y(n62733) );
  NAND2X1 U66817 ( .A(n42022), .B(n62733), .Y(n62734) );
  NAND2X1 U66818 ( .A(n62735), .B(n62734), .Y(n62736) );
  NAND2X1 U66819 ( .A(n62737), .B(n62736), .Y(n62740) );
  INVX1 U66820 ( .A(n62736), .Y(n68225) );
  INVX1 U66821 ( .A(n62737), .Y(n68224) );
  NAND2X1 U66822 ( .A(n68225), .B(n68224), .Y(n62738) );
  NAND2X1 U66823 ( .A(n42036), .B(n62738), .Y(n62739) );
  NAND2X1 U66824 ( .A(n62740), .B(n62739), .Y(n62742) );
  NAND2X1 U66825 ( .A(n62741), .B(n62742), .Y(n62745) );
  INVX1 U66826 ( .A(n62742), .Y(n68532) );
  NAND2X1 U66827 ( .A(n68532), .B(n68533), .Y(n62743) );
  NAND2X1 U66828 ( .A(n42049), .B(n62743), .Y(n62744) );
  NAND2X1 U66829 ( .A(n62745), .B(n62744), .Y(n62747) );
  NAND2X1 U66830 ( .A(n62746), .B(n62747), .Y(n62750) );
  INVX1 U66831 ( .A(n62747), .Y(n68849) );
  NAND2X1 U66832 ( .A(n68849), .B(n68850), .Y(n62748) );
  NAND2X1 U66833 ( .A(n42059), .B(n62748), .Y(n62749) );
  NAND2X1 U66834 ( .A(n62750), .B(n62749), .Y(n62751) );
  NAND2X1 U66835 ( .A(n62752), .B(n62751), .Y(n62755) );
  INVX1 U66836 ( .A(n62751), .Y(n69235) );
  INVX1 U66837 ( .A(n62752), .Y(n69234) );
  NAND2X1 U66838 ( .A(n69235), .B(n69234), .Y(n62753) );
  NAND2X1 U66839 ( .A(n42070), .B(n62753), .Y(n62754) );
  NAND2X1 U66840 ( .A(n62755), .B(n62754), .Y(n69567) );
  NAND2X1 U66841 ( .A(n62756), .B(n69567), .Y(n62759) );
  NAND2X1 U66842 ( .A(n37972), .B(n69566), .Y(n62757) );
  NAND2X1 U66843 ( .A(n42079), .B(n62757), .Y(n62758) );
  NAND2X1 U66844 ( .A(n62759), .B(n62758), .Y(n62761) );
  NAND2X1 U66845 ( .A(n62760), .B(n62761), .Y(n62764) );
  INVX1 U66846 ( .A(n62761), .Y(n69906) );
  NAND2X1 U66847 ( .A(n69906), .B(n69907), .Y(n62762) );
  NAND2X1 U66848 ( .A(n42089), .B(n62762), .Y(n62763) );
  NAND2X1 U66849 ( .A(n62764), .B(n62763), .Y(n62766) );
  NAND2X1 U66850 ( .A(n62765), .B(n62766), .Y(n62769) );
  INVX1 U66851 ( .A(n62766), .Y(n70194) );
  NAND2X1 U66852 ( .A(n70194), .B(n70195), .Y(n62767) );
  NAND2X1 U66853 ( .A(n42097), .B(n62767), .Y(n62768) );
  NAND2X1 U66854 ( .A(n62769), .B(n62768), .Y(n62770) );
  NAND2X1 U66855 ( .A(n62771), .B(n62770), .Y(n62774) );
  INVX1 U66856 ( .A(n62770), .Y(n70496) );
  INVX1 U66857 ( .A(n62771), .Y(n70495) );
  NAND2X1 U66858 ( .A(n70496), .B(n70495), .Y(n62772) );
  NAND2X1 U66859 ( .A(n42103), .B(n62772), .Y(n62773) );
  NAND2X1 U66860 ( .A(n62774), .B(n62773), .Y(n70799) );
  NAND2X1 U66861 ( .A(n38066), .B(n70798), .Y(n62776) );
  INVX1 U66862 ( .A(n62778), .Y(n71121) );
  NAND2X1 U66863 ( .A(n36350), .B(n71121), .Y(n62779) );
  NAND2X1 U66864 ( .A(n71408), .B(n62780), .Y(n62785) );
  NAND2X1 U66865 ( .A(n43729), .B(n44018), .Y(n71410) );
  INVX1 U66866 ( .A(n71410), .Y(n62783) );
  INVX1 U66867 ( .A(n71408), .Y(n62781) );
  NAND2X1 U66868 ( .A(n36353), .B(n62781), .Y(n62782) );
  NAND2X1 U66869 ( .A(n62783), .B(n62782), .Y(n62784) );
  NAND2X1 U66870 ( .A(n62785), .B(n62784), .Y(n62787) );
  INVX1 U66871 ( .A(n62787), .Y(n71717) );
  NAND2X1 U66872 ( .A(n71717), .B(n71718), .Y(n62788) );
  NAND2X1 U66873 ( .A(n62789), .B(n72113), .Y(n62793) );
  INVX1 U66874 ( .A(n72113), .Y(n62790) );
  NAND2X1 U66875 ( .A(n62790), .B(n72112), .Y(n62791) );
  NAND2X1 U66876 ( .A(n42129), .B(n62791), .Y(n62792) );
  NAND2X1 U66877 ( .A(n62793), .B(n62792), .Y(n62794) );
  INVX1 U66878 ( .A(n62794), .Y(n72128) );
  INVX1 U66879 ( .A(n62795), .Y(n72127) );
  NAND2X1 U66880 ( .A(n72128), .B(n72127), .Y(n62796) );
  NAND2X1 U66881 ( .A(n62797), .B(n72730), .Y(n62798) );
  XNOR2X1 U66882 ( .A(n62800), .B(n41497), .Y(n62804) );
  NAND2X1 U66883 ( .A(n43729), .B(n42720), .Y(n62802) );
  NOR2X1 U66884 ( .A(n39625), .B(n43754), .Y(n62801) );
  XNOR2X1 U66885 ( .A(n62802), .B(n62801), .Y(n62803) );
  INVX1 U66886 ( .A(n72732), .Y(n72728) );
  MX2X1 U66887 ( .A(n62804), .B(n62803), .S0(n43718), .Y(u_muldiv_result_r[1])
         );
  NAND2X1 U66888 ( .A(n44631), .B(u_muldiv_mult_result_q[1]), .Y(n14134) );
  NAND2X1 U66889 ( .A(n62805), .B(n43699), .Y(n62810) );
  INVX1 U66890 ( .A(n62805), .Y(n62806) );
  NAND2X1 U66891 ( .A(n43703), .B(n62806), .Y(n62807) );
  NAND2X1 U66892 ( .A(n62808), .B(n62807), .Y(n62809) );
  NAND2X1 U66893 ( .A(n62812), .B(n62811), .Y(n62816) );
  INVX1 U66894 ( .A(n62812), .Y(n62813) );
  NAND2X1 U66895 ( .A(n42126), .B(n62814), .Y(n62815) );
  NAND2X1 U66896 ( .A(n62818), .B(n62817), .Y(n62822) );
  NAND2X1 U66897 ( .A(n42101), .B(n62820), .Y(n62821) );
  NAND2X1 U66898 ( .A(n62822), .B(n62821), .Y(n63388) );
  NAND2X1 U66899 ( .A(n62828), .B(n62827), .Y(n63445) );
  OR2X1 U66900 ( .A(n62830), .B(n62829), .Y(n63444) );
  NAND2X1 U66901 ( .A(n43735), .B(n44001), .Y(n63112) );
  NAND2X1 U66902 ( .A(n62831), .B(n38164), .Y(n62835) );
  NAND2X1 U66903 ( .A(n40028), .B(n62832), .Y(n62833) );
  NAND2X1 U66904 ( .A(n42028), .B(n62833), .Y(n62834) );
  NAND2X1 U66905 ( .A(n62835), .B(n62834), .Y(n63117) );
  NAND2X1 U66906 ( .A(n43758), .B(n43993), .Y(n63115) );
  NOR2X1 U66907 ( .A(n62839), .B(n41268), .Y(n62836) );
  NOR2X1 U66908 ( .A(n62837), .B(n62836), .Y(n62841) );
  OR2X1 U66909 ( .A(n62839), .B(n62838), .Y(n62840) );
  NOR2X1 U66910 ( .A(n62843), .B(n62846), .Y(n62845) );
  NOR2X1 U66911 ( .A(n62843), .B(n62842), .Y(n62844) );
  INVX1 U66912 ( .A(n62846), .Y(n62848) );
  NOR2X1 U66913 ( .A(n43914), .B(n62849), .Y(n62854) );
  NAND2X1 U66914 ( .A(n62850), .B(n43911), .Y(n62852) );
  NAND2X1 U66915 ( .A(n62852), .B(n62851), .Y(n62853) );
  NOR2X1 U66916 ( .A(n62854), .B(n62853), .Y(n62856) );
  NAND2X1 U66917 ( .A(n62856), .B(n62855), .Y(n62857) );
  NAND2X1 U66918 ( .A(n41966), .B(n62857), .Y(n63134) );
  NAND2X1 U66919 ( .A(n62859), .B(n62858), .Y(n63135) );
  NAND2X1 U66920 ( .A(n63134), .B(n63135), .Y(n63025) );
  NAND2X1 U66921 ( .A(n43919), .B(n43788), .Y(n63144) );
  NOR2X1 U66922 ( .A(n62863), .B(n39827), .Y(n62866) );
  NOR2X1 U66923 ( .A(n62864), .B(n62863), .Y(n62865) );
  INVX1 U66924 ( .A(n63629), .Y(n63149) );
  INVX1 U66925 ( .A(n63345), .Y(n63348) );
  NAND2X1 U66926 ( .A(n63340), .B(n63341), .Y(n63358) );
  NAND2X1 U66927 ( .A(n62871), .B(n62870), .Y(n63159) );
  NAND2X1 U66928 ( .A(n63157), .B(n63158), .Y(n62872) );
  NAND2X1 U66929 ( .A(n63159), .B(n62872), .Y(n62996) );
  INVX1 U66930 ( .A(n62874), .Y(n63168) );
  NAND2X1 U66931 ( .A(n63168), .B(n63167), .Y(n62876) );
  NAND2X1 U66932 ( .A(n63169), .B(n62876), .Y(n63152) );
  NAND2X1 U66933 ( .A(n63306), .B(n62880), .Y(n63308) );
  INVX1 U66934 ( .A(n63305), .Y(n63307) );
  NAND2X1 U66935 ( .A(n39296), .B(n62881), .Y(n62882) );
  NOR2X1 U66936 ( .A(n41061), .B(n41085), .Y(n62884) );
  NAND2X1 U66937 ( .A(n40960), .B(n62885), .Y(n62889) );
  NAND2X1 U66938 ( .A(n43860), .B(n43478), .Y(n63295) );
  NAND2X1 U66939 ( .A(n62886), .B(n63291), .Y(n63287) );
  NAND2X1 U66940 ( .A(n63295), .B(n63287), .Y(n62887) );
  NOR2X1 U66941 ( .A(n62888), .B(n62887), .Y(n62893) );
  OR2X1 U66942 ( .A(n63295), .B(n63287), .Y(n62891) );
  NAND2X1 U66943 ( .A(n62891), .B(n62890), .Y(n62892) );
  NOR2X1 U66944 ( .A(n62892), .B(n62893), .Y(n63301) );
  NAND2X1 U66945 ( .A(n39941), .B(n43502), .Y(n63235) );
  NOR2X1 U66946 ( .A(n40627), .B(n38235), .Y(n62894) );
  NAND2X1 U66947 ( .A(n63556), .B(n63555), .Y(n63563) );
  NAND2X1 U66948 ( .A(n62894), .B(n63563), .Y(n63816) );
  INVX1 U66949 ( .A(n62895), .Y(n62901) );
  NAND2X1 U66950 ( .A(n38799), .B(n38804), .Y(n62898) );
  NOR2X1 U66951 ( .A(n36772), .B(n62898), .Y(n62899) );
  NOR2X1 U66952 ( .A(n62899), .B(n42799), .Y(n62900) );
  NOR2X1 U66953 ( .A(n62901), .B(n62900), .Y(n62914) );
  INVX1 U66954 ( .A(n62902), .Y(n62912) );
  NOR2X1 U66955 ( .A(n62904), .B(n62903), .Y(n62906) );
  NOR2X1 U66956 ( .A(n62906), .B(n62905), .Y(n62908) );
  NAND2X1 U66957 ( .A(n62908), .B(n62907), .Y(n62910) );
  NAND2X1 U66958 ( .A(n62910), .B(n62909), .Y(n62911) );
  NOR2X1 U66959 ( .A(n62912), .B(n62911), .Y(n62913) );
  NOR2X1 U66960 ( .A(n42236), .B(n64087), .Y(n62921) );
  NOR2X1 U66961 ( .A(n62915), .B(n43450), .Y(n62918) );
  NOR2X1 U66962 ( .A(n62916), .B(n42800), .Y(n62917) );
  OR2X1 U66963 ( .A(n62918), .B(n62917), .Y(n62919) );
  NOR2X1 U66964 ( .A(n63190), .B(n62919), .Y(n63182) );
  NOR2X1 U66965 ( .A(n63182), .B(n64087), .Y(n62920) );
  XNOR2X1 U66966 ( .A(n62921), .B(n62920), .Y(n63562) );
  NOR2X1 U66967 ( .A(n43611), .B(n63562), .Y(n62922) );
  XNOR2X1 U66968 ( .A(n63199), .B(n62922), .Y(n63231) );
  INVX1 U66969 ( .A(n63221), .Y(n63224) );
  NAND2X1 U66970 ( .A(n62940), .B(n62939), .Y(n62926) );
  NAND2X1 U66971 ( .A(n38691), .B(n62926), .Y(n62924) );
  NAND2X1 U66972 ( .A(n62924), .B(n63226), .Y(n62925) );
  NOR2X1 U66973 ( .A(n63224), .B(n62925), .Y(n62936) );
  NAND2X1 U66974 ( .A(n38514), .B(n62926), .Y(n62927) );
  NAND2X1 U66975 ( .A(n38691), .B(n38514), .Y(n62930) );
  NAND2X1 U66976 ( .A(n62927), .B(n62930), .Y(n62928) );
  NAND2X1 U66977 ( .A(n62928), .B(n63224), .Y(n62934) );
  NAND2X1 U66978 ( .A(n63226), .B(n62929), .Y(n63229) );
  NAND2X1 U66979 ( .A(n39621), .B(n63229), .Y(n62932) );
  NAND2X1 U66980 ( .A(n62930), .B(n62941), .Y(n62931) );
  NAND2X1 U66981 ( .A(n62932), .B(n62931), .Y(n62933) );
  NAND2X1 U66982 ( .A(n62934), .B(n62933), .Y(n62935) );
  NOR2X1 U66983 ( .A(n62936), .B(n62935), .Y(n62937) );
  XNOR2X1 U66984 ( .A(n63235), .B(n63241), .Y(n62949) );
  NAND2X1 U66985 ( .A(n62940), .B(n62939), .Y(n62941) );
  XNOR2X1 U66986 ( .A(n62941), .B(n38691), .Y(n62942) );
  XNOR2X1 U66987 ( .A(n63224), .B(n62942), .Y(n62948) );
  INVX1 U66988 ( .A(n62943), .Y(n62944) );
  NOR2X1 U66989 ( .A(n62944), .B(n41770), .Y(n62946) );
  NAND2X1 U66990 ( .A(n62946), .B(n62945), .Y(n62947) );
  NAND2X1 U66991 ( .A(n62948), .B(n62947), .Y(n63239) );
  NAND2X1 U66992 ( .A(n63237), .B(n63239), .Y(n63236) );
  INVX1 U66993 ( .A(n63249), .Y(n63243) );
  INVX1 U66994 ( .A(n63245), .Y(n63254) );
  NAND2X1 U66995 ( .A(n43840), .B(n43497), .Y(n63244) );
  NOR2X1 U66996 ( .A(n62953), .B(n62952), .Y(n62956) );
  INVX1 U66997 ( .A(n63244), .Y(n63250) );
  NOR2X1 U66998 ( .A(n63253), .B(n63244), .Y(n62954) );
  NOR2X1 U66999 ( .A(n62955), .B(n62956), .Y(n62957) );
  XNOR2X1 U67000 ( .A(n63243), .B(n62957), .Y(n63178) );
  NOR2X1 U67001 ( .A(n40094), .B(n62958), .Y(n62961) );
  INVX1 U67002 ( .A(n62963), .Y(n62959) );
  NOR2X1 U67003 ( .A(n62959), .B(n62958), .Y(n62960) );
  NAND2X1 U67004 ( .A(n43493), .B(n38382), .Y(n63175) );
  NOR2X1 U67005 ( .A(n40015), .B(n62977), .Y(n62966) );
  NOR2X1 U67006 ( .A(n40015), .B(n62978), .Y(n62965) );
  NOR2X1 U67007 ( .A(n62966), .B(n62965), .Y(n62970) );
  INVX1 U67008 ( .A(n62977), .Y(n62967) );
  NAND2X1 U67009 ( .A(n62968), .B(n62967), .Y(n62969) );
  NAND2X1 U67010 ( .A(n62970), .B(n62969), .Y(n63269) );
  NAND2X1 U67011 ( .A(n44035), .B(n38311), .Y(n63264) );
  INVX1 U67012 ( .A(n63283), .Y(n63293) );
  XNOR2X1 U67013 ( .A(n37407), .B(n63293), .Y(n62991) );
  NOR2X1 U67014 ( .A(n40024), .B(n62971), .Y(n63275) );
  INVX1 U67015 ( .A(n62972), .Y(n62974) );
  NOR2X1 U67016 ( .A(n62974), .B(n38465), .Y(n62975) );
  NAND2X1 U67017 ( .A(n62976), .B(n62975), .Y(n62980) );
  XNOR2X1 U67018 ( .A(n62978), .B(n62977), .Y(n62979) );
  XNOR2X1 U67019 ( .A(n62980), .B(n62979), .Y(n63278) );
  INVX1 U67020 ( .A(n63278), .Y(n62981) );
  NOR2X1 U67021 ( .A(n39771), .B(n63274), .Y(n62986) );
  NAND2X1 U67022 ( .A(n43851), .B(n38313), .Y(n63280) );
  NOR2X1 U67023 ( .A(n38432), .B(n40014), .Y(n62983) );
  NAND2X1 U67024 ( .A(n62983), .B(n62982), .Y(n62984) );
  NAND2X1 U67025 ( .A(n63278), .B(n62984), .Y(n63273) );
  NAND2X1 U67026 ( .A(n63280), .B(n63273), .Y(n62985) );
  NOR2X1 U67027 ( .A(n62986), .B(n62985), .Y(n62990) );
  OR2X1 U67028 ( .A(n63280), .B(n63273), .Y(n62987) );
  NAND2X1 U67029 ( .A(n62988), .B(n62987), .Y(n62989) );
  NOR2X1 U67030 ( .A(n62990), .B(n62989), .Y(n63294) );
  XNOR2X1 U67031 ( .A(n62991), .B(n63294), .Y(n62992) );
  XNOR2X1 U67032 ( .A(n39910), .B(n41394), .Y(n63172) );
  NAND2X1 U67033 ( .A(n43870), .B(n42714), .Y(n63161) );
  NAND2X1 U67034 ( .A(n43952), .B(n43796), .Y(n63166) );
  XNOR2X1 U67035 ( .A(n63161), .B(n63166), .Y(n62993) );
  XNOR2X1 U67036 ( .A(n63172), .B(n62993), .Y(n62994) );
  XNOR2X1 U67037 ( .A(n63152), .B(n62994), .Y(n62995) );
  XOR2X1 U67038 ( .A(n62996), .B(n62995), .Y(n63327) );
  NAND2X1 U67039 ( .A(n38981), .B(n39423), .Y(n63318) );
  NAND2X1 U67040 ( .A(n38902), .B(n63322), .Y(n63319) );
  NAND2X1 U67041 ( .A(n42661), .B(n43880), .Y(n63000) );
  NOR2X1 U67042 ( .A(n39724), .B(n62999), .Y(n63005) );
  NAND2X1 U67043 ( .A(n40480), .B(n38896), .Y(n63003) );
  NAND2X1 U67044 ( .A(n63001), .B(n38896), .Y(n63002) );
  NAND2X1 U67045 ( .A(n63003), .B(n63002), .Y(n63004) );
  NOR2X1 U67046 ( .A(n63005), .B(n63004), .Y(n63006) );
  XNOR2X1 U67047 ( .A(n63327), .B(n63006), .Y(n63338) );
  INVX1 U67048 ( .A(n63338), .Y(n63335) );
  NAND2X1 U67049 ( .A(n63008), .B(n63007), .Y(n63012) );
  NAND2X1 U67050 ( .A(n63010), .B(n63009), .Y(n63011) );
  INVX1 U67051 ( .A(n63014), .Y(n63016) );
  NAND2X1 U67052 ( .A(n63016), .B(n63015), .Y(n63331) );
  XNOR2X1 U67053 ( .A(n63335), .B(n41120), .Y(n63361) );
  NAND2X1 U67054 ( .A(n43798), .B(n43890), .Y(n63329) );
  INVX1 U67055 ( .A(n63329), .Y(n63337) );
  XNOR2X1 U67056 ( .A(n63337), .B(n42182), .Y(n63359) );
  INVX1 U67057 ( .A(n63611), .Y(n63364) );
  XNOR2X1 U67058 ( .A(n63359), .B(n63364), .Y(n63017) );
  XNOR2X1 U67059 ( .A(n63358), .B(n63018), .Y(n63146) );
  XNOR2X1 U67060 ( .A(n41922), .B(n63146), .Y(n63021) );
  INVX1 U67061 ( .A(n63612), .Y(n63147) );
  XNOR2X1 U67062 ( .A(n63021), .B(n63147), .Y(n63022) );
  XNOR2X1 U67063 ( .A(n63144), .B(n36697), .Y(n63023) );
  XNOR2X1 U67064 ( .A(n41259), .B(n63023), .Y(n63139) );
  NAND2X1 U67065 ( .A(n43926), .B(n40484), .Y(n63136) );
  XNOR2X1 U67066 ( .A(n63139), .B(n63136), .Y(n63024) );
  XNOR2X1 U67067 ( .A(n63025), .B(n63024), .Y(n63131) );
  XNOR2X1 U67068 ( .A(n63131), .B(n41983), .Y(n63026) );
  XNOR2X1 U67069 ( .A(n63130), .B(n41994), .Y(n63027) );
  INVX1 U67070 ( .A(n63455), .Y(n63380) );
  NAND2X1 U67071 ( .A(n63371), .B(n63029), .Y(n63374) );
  NAND2X1 U67072 ( .A(n63030), .B(n63374), .Y(n63378) );
  NAND2X1 U67073 ( .A(n43809), .B(n43974), .Y(n63377) );
  INVX1 U67074 ( .A(n63377), .Y(n63381) );
  XNOR2X1 U67075 ( .A(n63378), .B(n63381), .Y(n63031) );
  XNOR2X1 U67076 ( .A(n63380), .B(n63031), .Y(n63128) );
  NAND2X1 U67077 ( .A(n43820), .B(n43984), .Y(n63119) );
  NOR2X1 U67078 ( .A(n63036), .B(n63121), .Y(n63038) );
  NAND2X1 U67079 ( .A(n40279), .B(n38598), .Y(n63040) );
  NAND2X1 U67080 ( .A(n63040), .B(n63039), .Y(n63037) );
  NOR2X1 U67081 ( .A(n63038), .B(n41326), .Y(n63043) );
  NAND2X1 U67082 ( .A(n63039), .B(n63040), .Y(n63120) );
  NAND2X1 U67083 ( .A(n63041), .B(n39478), .Y(n63042) );
  NAND2X1 U67084 ( .A(n63043), .B(n63042), .Y(n63127) );
  XNOR2X1 U67085 ( .A(n63115), .B(n37382), .Y(n63044) );
  XNOR2X1 U67086 ( .A(n36454), .B(n63044), .Y(n63447) );
  INVX1 U67087 ( .A(n63447), .Y(n63113) );
  XNOR2X1 U67088 ( .A(n63112), .B(n63113), .Y(n63045) );
  XNOR2X1 U67089 ( .A(n39987), .B(n63045), .Y(n63111) );
  INVX1 U67090 ( .A(n63111), .Y(n63109) );
  NAND2X1 U67091 ( .A(n63048), .B(n63047), .Y(n63049) );
  OR2X1 U67092 ( .A(n36782), .B(n63049), .Y(n63050) );
  XNOR2X1 U67093 ( .A(n63110), .B(n42073), .Y(n63051) );
  XNOR2X1 U67094 ( .A(n63109), .B(n63051), .Y(n63104) );
  INVX1 U67095 ( .A(n63104), .Y(n63106) );
  XNOR2X1 U67096 ( .A(n63105), .B(n63106), .Y(n63052) );
  XNOR2X1 U67097 ( .A(n42085), .B(n63052), .Y(n63101) );
  INVX1 U67098 ( .A(n63099), .Y(n63102) );
  XNOR2X1 U67099 ( .A(n63101), .B(n63102), .Y(n63057) );
  XNOR2X1 U67100 ( .A(n42100), .B(n63057), .Y(n63387) );
  INVX1 U67101 ( .A(n63387), .Y(n63389) );
  XNOR2X1 U67102 ( .A(n63388), .B(n63389), .Y(n63058) );
  XNOR2X1 U67103 ( .A(n42107), .B(n63058), .Y(n63095) );
  INVX1 U67104 ( .A(n63060), .Y(n63062) );
  NAND2X1 U67105 ( .A(n63062), .B(n63061), .Y(n63063) );
  XNOR2X1 U67106 ( .A(n63095), .B(n38119), .Y(n63064) );
  XNOR2X1 U67107 ( .A(n42120), .B(n63064), .Y(n63090) );
  NAND2X1 U67108 ( .A(n43612), .B(n43816), .Y(n71734) );
  XNOR2X1 U67109 ( .A(n63090), .B(n43508), .Y(n63065) );
  XNOR2X1 U67110 ( .A(n41674), .B(n63065), .Y(n63085) );
  XNOR2X1 U67111 ( .A(n63085), .B(n43692), .Y(n63066) );
  XNOR2X1 U67112 ( .A(n41487), .B(n63066), .Y(n63078) );
  INVX1 U67113 ( .A(n63078), .Y(n63079) );
  XNOR2X1 U67114 ( .A(n43709), .B(n63079), .Y(n63072) );
  NAND2X1 U67115 ( .A(n63067), .B(n43712), .Y(n63071) );
  NAND2X1 U67116 ( .A(n43706), .B(n63068), .Y(n63069) );
  NAND2X1 U67117 ( .A(n41497), .B(n63069), .Y(n63070) );
  NAND2X1 U67118 ( .A(n63071), .B(n63070), .Y(n63080) );
  XNOR2X1 U67119 ( .A(n63072), .B(n36356), .Y(n63077) );
  XNOR2X1 U67120 ( .A(n41866), .B(n63073), .Y(n63075) );
  XNOR2X1 U67121 ( .A(n63075), .B(n63074), .Y(n63076) );
  MX2X1 U67122 ( .A(n63077), .B(n63076), .S0(n43720), .Y(u_muldiv_result_r[2])
         );
  NOR2X1 U67123 ( .A(n1889), .B(n37333), .Y(n14130) );
  NAND2X1 U67124 ( .A(n63078), .B(n43714), .Y(n63083) );
  NAND2X1 U67125 ( .A(n43706), .B(n63079), .Y(n63081) );
  NAND2X1 U67126 ( .A(n63081), .B(n63080), .Y(n63082) );
  INVX1 U67127 ( .A(n63085), .Y(n63084) );
  NAND2X1 U67128 ( .A(n41466), .B(n63084), .Y(n63088) );
  NAND2X1 U67129 ( .A(n63085), .B(n43701), .Y(n63086) );
  NAND2X1 U67130 ( .A(n41487), .B(n63086), .Y(n63087) );
  AND2X1 U67131 ( .A(n63088), .B(n63087), .Y(n63410) );
  INVX1 U67132 ( .A(n63090), .Y(n63089) );
  NAND2X1 U67133 ( .A(n63089), .B(n43513), .Y(n63093) );
  NAND2X1 U67134 ( .A(n43506), .B(n63090), .Y(n63091) );
  NAND2X1 U67135 ( .A(n41674), .B(n63091), .Y(n63092) );
  AND2X1 U67136 ( .A(n63093), .B(n63092), .Y(n63416) );
  INVX1 U67137 ( .A(n63095), .Y(n63094) );
  NAND2X1 U67138 ( .A(n63094), .B(n38065), .Y(n63098) );
  NAND2X1 U67139 ( .A(n38119), .B(n63095), .Y(n63096) );
  NAND2X1 U67140 ( .A(n42120), .B(n63096), .Y(n63097) );
  NAND2X1 U67141 ( .A(n63098), .B(n63097), .Y(n63421) );
  INVX1 U67142 ( .A(n63101), .Y(n63100) );
  INVX1 U67143 ( .A(n63105), .Y(n63107) );
  NAND2X1 U67144 ( .A(n63107), .B(n63106), .Y(n63108) );
  NAND2X1 U67145 ( .A(n63109), .B(n63110), .Y(n63431) );
  NAND2X1 U67146 ( .A(n63431), .B(n63432), .Y(n63430) );
  NAND2X1 U67147 ( .A(n63114), .B(n63443), .Y(n63441) );
  INVX1 U67148 ( .A(n63115), .Y(n63116) );
  NAND2X1 U67149 ( .A(n63116), .B(n63672), .Y(n63118) );
  NAND2X1 U67150 ( .A(n63118), .B(n63673), .Y(n63671) );
  INVX1 U67151 ( .A(n63119), .Y(n63126) );
  NOR2X1 U67152 ( .A(n38295), .B(n63120), .Y(n63122) );
  NOR2X1 U67153 ( .A(n63122), .B(n63121), .Y(n63123) );
  NOR2X1 U67154 ( .A(n41326), .B(n63123), .Y(n63125) );
  INVX1 U67155 ( .A(n63128), .Y(n63124) );
  NAND2X1 U67156 ( .A(n63125), .B(n63124), .Y(n63669) );
  NAND2X1 U67157 ( .A(n63126), .B(n63669), .Y(n63129) );
  NAND2X1 U67158 ( .A(n63129), .B(n63670), .Y(n63667) );
  NAND2X1 U67159 ( .A(n41994), .B(n63130), .Y(n63903) );
  INVX1 U67160 ( .A(n63659), .Y(n63656) );
  NAND2X1 U67161 ( .A(n40461), .B(n43974), .Y(n63657) );
  INVX1 U67162 ( .A(n63131), .Y(n63133) );
  NAND2X1 U67163 ( .A(n63135), .B(n63134), .Y(n63467) );
  NOR2X1 U67164 ( .A(n39881), .B(n63136), .Y(n63138) );
  INVX1 U67165 ( .A(n63139), .Y(n63464) );
  NOR2X1 U67166 ( .A(n63464), .B(n63136), .Y(n63137) );
  NAND2X1 U67167 ( .A(n63642), .B(n63144), .Y(n63143) );
  OR2X1 U67168 ( .A(n63642), .B(n63144), .Y(n63145) );
  INVX1 U67169 ( .A(n63649), .Y(n63369) );
  INVX1 U67170 ( .A(n63626), .Y(n63148) );
  NOR2X1 U67171 ( .A(n63149), .B(n63148), .Y(n63151) );
  NAND2X1 U67172 ( .A(n41922), .B(n63626), .Y(n63627) );
  NAND2X1 U67173 ( .A(n42661), .B(n43890), .Y(n63485) );
  INVX1 U67174 ( .A(n63166), .Y(n63174) );
  XNOR2X1 U67175 ( .A(n63174), .B(n39768), .Y(n63153) );
  XNOR2X1 U67176 ( .A(n63153), .B(n41394), .Y(n63154) );
  INVX1 U67177 ( .A(n63162), .Y(n63155) );
  INVX1 U67178 ( .A(n63156), .Y(n63158) );
  NAND2X1 U67179 ( .A(n63158), .B(n63157), .Y(n63160) );
  INVX1 U67180 ( .A(n63161), .Y(n63163) );
  NAND2X1 U67181 ( .A(n63163), .B(n63162), .Y(n63164) );
  NAND2X1 U67182 ( .A(n63165), .B(n63164), .Y(n63493) );
  NAND2X1 U67183 ( .A(n63172), .B(n63166), .Y(n63171) );
  NAND2X1 U67184 ( .A(n62876), .B(n63169), .Y(n63170) );
  INVX1 U67185 ( .A(n63172), .Y(n63173) );
  NAND2X1 U67186 ( .A(n43871), .B(n43796), .Y(n63593) );
  NAND2X1 U67187 ( .A(n43861), .B(n43484), .Y(n63514) );
  NOR2X1 U67188 ( .A(n63177), .B(n63176), .Y(n63180) );
  NAND2X1 U67189 ( .A(n63178), .B(n40241), .Y(n63179) );
  NAND2X1 U67190 ( .A(n63180), .B(n63179), .Y(n63521) );
  NAND2X1 U67191 ( .A(n43492), .B(n44037), .Y(n63524) );
  NAND2X1 U67192 ( .A(n43603), .B(n63209), .Y(n63181) );
  NOR2X1 U67193 ( .A(n43611), .B(n63181), .Y(n63187) );
  XNOR2X1 U67194 ( .A(n42236), .B(n63182), .Y(n63185) );
  NAND2X1 U67195 ( .A(n43603), .B(n63183), .Y(n63184) );
  NOR2X1 U67196 ( .A(n63185), .B(n63184), .Y(n63186) );
  XNOR2X1 U67197 ( .A(n63187), .B(n63186), .Y(n63565) );
  NAND2X1 U67198 ( .A(n39937), .B(n39960), .Y(n63548) );
  INVX1 U67199 ( .A(n63548), .Y(n63547) );
  NOR2X1 U67200 ( .A(n42799), .B(n64087), .Y(n63189) );
  NAND2X1 U67201 ( .A(n63189), .B(n63188), .Y(n63192) );
  NAND2X1 U67202 ( .A(n43603), .B(n63190), .Y(n63191) );
  NAND2X1 U67203 ( .A(n63192), .B(n63191), .Y(n63195) );
  NOR2X1 U67204 ( .A(n63196), .B(n63193), .Y(n63198) );
  NAND2X1 U67205 ( .A(n63195), .B(n43609), .Y(n63196) );
  NOR2X1 U67206 ( .A(n36719), .B(n63196), .Y(n63197) );
  NOR2X1 U67207 ( .A(n63198), .B(n63197), .Y(n63571) );
  XNOR2X1 U67208 ( .A(n63547), .B(n63571), .Y(n63219) );
  NOR2X1 U67209 ( .A(n63200), .B(n42800), .Y(n63202) );
  NOR2X1 U67210 ( .A(n42379), .B(n42799), .Y(n63201) );
  NOR2X1 U67211 ( .A(n63202), .B(n63201), .Y(n63203) );
  NAND2X1 U67212 ( .A(n63203), .B(n42515), .Y(n63205) );
  NAND2X1 U67213 ( .A(n63205), .B(n39653), .Y(n63552) );
  NAND2X1 U67214 ( .A(n38305), .B(n63552), .Y(n63204) );
  NOR2X1 U67215 ( .A(n63204), .B(n38500), .Y(n63215) );
  INVX1 U67216 ( .A(n63205), .Y(n63569) );
  NOR2X1 U67217 ( .A(n63569), .B(n38592), .Y(n63207) );
  NOR2X1 U67218 ( .A(n43476), .B(n63205), .Y(n63206) );
  NOR2X1 U67219 ( .A(n63207), .B(n63206), .Y(n63213) );
  NOR2X1 U67220 ( .A(n63208), .B(n63830), .Y(n63210) );
  NAND2X1 U67221 ( .A(n63210), .B(n38644), .Y(n63211) );
  NAND2X1 U67222 ( .A(n63211), .B(n43608), .Y(n63212) );
  NOR2X1 U67223 ( .A(n63213), .B(n63212), .Y(n63214) );
  NOR2X1 U67224 ( .A(n63215), .B(n63214), .Y(n63218) );
  NOR2X1 U67225 ( .A(n63552), .B(n38610), .Y(n63216) );
  NAND2X1 U67226 ( .A(n63216), .B(n63816), .Y(n63217) );
  XNOR2X1 U67227 ( .A(n63219), .B(n41801), .Y(n63220) );
  XNOR2X1 U67228 ( .A(n63565), .B(n63220), .Y(n63234) );
  NAND2X1 U67229 ( .A(n39621), .B(n63221), .Y(n63230) );
  NAND2X1 U67230 ( .A(n63230), .B(n43472), .Y(n63223) );
  NOR2X1 U67231 ( .A(n63226), .B(n63223), .Y(n63228) );
  NAND2X1 U67232 ( .A(n63224), .B(n62941), .Y(n63225) );
  NOR2X1 U67233 ( .A(n63226), .B(n63225), .Y(n63227) );
  XNOR2X1 U67234 ( .A(n63816), .B(n63231), .Y(n63232) );
  NAND2X1 U67235 ( .A(n43840), .B(n43502), .Y(n63543) );
  INVX1 U67236 ( .A(n63235), .Y(n63238) );
  NOR2X1 U67237 ( .A(n63238), .B(n38205), .Y(n63240) );
  NAND2X1 U67238 ( .A(n63240), .B(n63239), .Y(n63242) );
  INVX1 U67239 ( .A(n63253), .Y(n63246) );
  NAND2X1 U67240 ( .A(n63246), .B(n63245), .Y(n63248) );
  NAND2X1 U67241 ( .A(n63248), .B(n63247), .Y(n63532) );
  NAND2X1 U67242 ( .A(n63250), .B(n63249), .Y(n63534) );
  NAND2X1 U67243 ( .A(n38380), .B(n43496), .Y(n63530) );
  NAND2X1 U67244 ( .A(n63534), .B(n63530), .Y(n63251) );
  NOR2X1 U67245 ( .A(n63252), .B(n63251), .Y(n63262) );
  OR2X1 U67246 ( .A(n63530), .B(n63534), .Y(n63260) );
  NOR2X1 U67247 ( .A(n63254), .B(n63253), .Y(n63255) );
  INVX1 U67248 ( .A(n63530), .Y(n63529) );
  NAND2X1 U67249 ( .A(n63255), .B(n63529), .Y(n63257) );
  NAND2X1 U67250 ( .A(n63529), .B(n40237), .Y(n63256) );
  NAND2X1 U67251 ( .A(n63257), .B(n63256), .Y(n63258) );
  NAND2X1 U67252 ( .A(n63258), .B(n63533), .Y(n63259) );
  NAND2X1 U67253 ( .A(n63260), .B(n63259), .Y(n63261) );
  NOR2X1 U67254 ( .A(n63262), .B(n63261), .Y(n63263) );
  XOR2X1 U67255 ( .A(n63531), .B(n63263), .Y(n63525) );
  NAND2X1 U67256 ( .A(n43851), .B(n43487), .Y(n63579) );
  NOR2X1 U67257 ( .A(n63268), .B(n63264), .Y(n63267) );
  INVX1 U67258 ( .A(n63269), .Y(n63265) );
  NOR2X1 U67259 ( .A(n63265), .B(n63264), .Y(n63266) );
  NOR2X1 U67260 ( .A(n63267), .B(n63266), .Y(n63272) );
  INVX1 U67261 ( .A(n63268), .Y(n63270) );
  NAND2X1 U67262 ( .A(n63270), .B(n63269), .Y(n63271) );
  NAND2X1 U67263 ( .A(n63272), .B(n63271), .Y(n63581) );
  INVX1 U67264 ( .A(n63273), .Y(n63277) );
  NOR2X1 U67265 ( .A(n63275), .B(n63274), .Y(n63276) );
  NOR2X1 U67266 ( .A(n38425), .B(n63280), .Y(n63282) );
  NOR2X1 U67267 ( .A(n63293), .B(n63280), .Y(n63281) );
  NOR2X1 U67268 ( .A(n63282), .B(n63281), .Y(n63286) );
  NAND2X1 U67269 ( .A(n63284), .B(n63283), .Y(n63285) );
  NAND2X1 U67270 ( .A(n63286), .B(n63285), .Y(n63516) );
  NAND2X1 U67271 ( .A(n43962), .B(n43478), .Y(n63509) );
  INVX1 U67272 ( .A(n63287), .Y(n63289) );
  NOR2X1 U67273 ( .A(n40960), .B(n63290), .Y(n63288) );
  INVX1 U67274 ( .A(n63290), .Y(n63292) );
  NOR2X1 U67275 ( .A(n63295), .B(n38976), .Y(n63297) );
  XNOR2X1 U67276 ( .A(n63294), .B(n63293), .Y(n63298) );
  INVX1 U67277 ( .A(n63298), .Y(n63300) );
  NOR2X1 U67278 ( .A(n63300), .B(n63295), .Y(n63296) );
  XOR2X1 U67279 ( .A(n63509), .B(n63511), .Y(n63299) );
  XNOR2X1 U67280 ( .A(n63301), .B(n63300), .Y(n63302) );
  NOR2X1 U67281 ( .A(n39910), .B(n38660), .Y(n63304) );
  NAND2X1 U67282 ( .A(n37407), .B(n63302), .Y(n63772) );
  NAND2X1 U67283 ( .A(n43952), .B(n43775), .Y(n63773) );
  NAND2X1 U67284 ( .A(n63772), .B(n63773), .Y(n63303) );
  NOR2X1 U67285 ( .A(n63304), .B(n63303), .Y(n63316) );
  INVX1 U67286 ( .A(n63773), .Y(n63502) );
  NOR2X1 U67287 ( .A(n39296), .B(n63305), .Y(n63311) );
  NAND2X1 U67288 ( .A(n63307), .B(n63306), .Y(n63309) );
  NAND2X1 U67289 ( .A(n63309), .B(n63308), .Y(n63310) );
  NOR2X1 U67290 ( .A(n63311), .B(n63310), .Y(n63312) );
  NAND2X1 U67291 ( .A(n63314), .B(n63313), .Y(n63315) );
  NOR2X1 U67292 ( .A(n63316), .B(n63315), .Y(n63317) );
  XNOR2X1 U67293 ( .A(n63507), .B(n63317), .Y(n63590) );
  NAND2X1 U67294 ( .A(n43879), .B(n42712), .Y(n63497) );
  XNOR2X1 U67295 ( .A(n63485), .B(n63491), .Y(n63328) );
  NOR2X1 U67296 ( .A(n63324), .B(n63320), .Y(n63321) );
  INVX1 U67297 ( .A(n63322), .Y(n63323) );
  NOR2X1 U67298 ( .A(n63324), .B(n63323), .Y(n63325) );
  NAND2X1 U67299 ( .A(n63327), .B(n63326), .Y(n63489) );
  NAND2X1 U67300 ( .A(n63487), .B(n63489), .Y(n63486) );
  NAND2X1 U67301 ( .A(n63338), .B(n63329), .Y(n63334) );
  NAND2X1 U67302 ( .A(n41325), .B(n63330), .Y(n63332) );
  NAND2X1 U67303 ( .A(n63332), .B(n63331), .Y(n63333) );
  NAND2X1 U67304 ( .A(n43798), .B(n43898), .Y(n63599) );
  NAND2X1 U67305 ( .A(n40259), .B(n43904), .Y(n63477) );
  XNOR2X1 U67306 ( .A(n63603), .B(n63336), .Y(n63633) );
  XNOR2X1 U67307 ( .A(n63338), .B(n63337), .Y(n63339) );
  XNOR2X1 U67308 ( .A(n41120), .B(n63339), .Y(n63344) );
  NOR2X1 U67309 ( .A(n40605), .B(n42182), .Y(n63342) );
  NAND2X1 U67310 ( .A(n63342), .B(n63341), .Y(n63343) );
  NOR2X1 U67311 ( .A(n39563), .B(n63345), .Y(n63346) );
  NOR2X1 U67312 ( .A(n40605), .B(n63346), .Y(n63350) );
  NAND2X1 U67313 ( .A(n63348), .B(n63347), .Y(n63349) );
  NAND2X1 U67314 ( .A(n63350), .B(n63349), .Y(n63351) );
  INVX1 U67315 ( .A(n63481), .Y(n63632) );
  XNOR2X1 U67316 ( .A(n63633), .B(n63632), .Y(n63609) );
  INVX1 U67317 ( .A(n63609), .Y(n63607) );
  NAND2X1 U67318 ( .A(n43918), .B(n43724), .Y(n63637) );
  XNOR2X1 U67319 ( .A(n63637), .B(n37412), .Y(n63352) );
  XNOR2X1 U67320 ( .A(n63607), .B(n63352), .Y(n63365) );
  NOR2X1 U67321 ( .A(n63353), .B(n63355), .Y(n63354) );
  NOR2X1 U67322 ( .A(n63356), .B(n63355), .Y(n63357) );
  INVX1 U67323 ( .A(n63359), .Y(n63360) );
  XNOR2X1 U67324 ( .A(n63361), .B(n63360), .Y(n63362) );
  INVX1 U67325 ( .A(n63614), .Y(n63363) );
  INVX1 U67326 ( .A(n63608), .Y(n63636) );
  XNOR2X1 U67327 ( .A(n63365), .B(n63636), .Y(n63366) );
  NAND2X1 U67328 ( .A(n40483), .B(n43935), .Y(n63463) );
  NAND2X1 U67329 ( .A(n43926), .B(n43788), .Y(n63646) );
  XNOR2X1 U67330 ( .A(n63463), .B(n63646), .Y(n63367) );
  XOR2X1 U67331 ( .A(n63650), .B(n63367), .Y(n63368) );
  INVX1 U67332 ( .A(n63905), .Y(n63658) );
  XNOR2X1 U67333 ( .A(n63657), .B(n63658), .Y(n63370) );
  XNOR2X1 U67334 ( .A(n63656), .B(n63370), .Y(n63919) );
  INVX1 U67335 ( .A(n63919), .Y(n63452) );
  NOR2X1 U67336 ( .A(n63028), .B(n63372), .Y(n63376) );
  OR2X1 U67337 ( .A(n38851), .B(n63372), .Y(n63373) );
  NAND2X1 U67338 ( .A(n63374), .B(n63373), .Y(n63375) );
  NOR2X1 U67339 ( .A(n63376), .B(n63375), .Y(n63456) );
  NOR2X1 U67340 ( .A(n63456), .B(n63377), .Y(n63379) );
  NAND2X1 U67341 ( .A(n43809), .B(n43984), .Y(n63920) );
  INVX1 U67342 ( .A(n63920), .Y(n63460) );
  XNOR2X1 U67343 ( .A(n63453), .B(n63460), .Y(n63382) );
  XNOR2X1 U67344 ( .A(n63452), .B(n63382), .Y(n63668) );
  NAND2X1 U67345 ( .A(n43758), .B(n44001), .Y(n63438) );
  NAND2X1 U67346 ( .A(n43735), .B(n44009), .Y(n63442) );
  XNOR2X1 U67347 ( .A(n63438), .B(n63442), .Y(n63383) );
  XOR2X1 U67348 ( .A(n63675), .B(n63383), .Y(n63384) );
  XNOR2X1 U67349 ( .A(n63428), .B(n42094), .Y(n63385) );
  XNOR2X1 U67350 ( .A(n38852), .B(n63385), .Y(n63423) );
  INVX1 U67351 ( .A(n63423), .Y(n63425) );
  XNOR2X1 U67352 ( .A(n63424), .B(n63425), .Y(n63386) );
  XNOR2X1 U67353 ( .A(n42106), .B(n63386), .Y(n63683) );
  INVX1 U67354 ( .A(n63388), .Y(n63390) );
  NAND2X1 U67355 ( .A(n63390), .B(n63389), .Y(n63391) );
  INVX1 U67356 ( .A(n63681), .Y(n63684) );
  XNOR2X1 U67357 ( .A(n63683), .B(n63684), .Y(n63392) );
  XNOR2X1 U67358 ( .A(n42113), .B(n63392), .Y(n63419) );
  NAND2X1 U67359 ( .A(n43612), .B(n43805), .Y(n72675) );
  XNOR2X1 U67360 ( .A(n63419), .B(n43679), .Y(n63393) );
  XNOR2X1 U67361 ( .A(n63414), .B(n43508), .Y(n63394) );
  XNOR2X1 U67362 ( .A(n63416), .B(n63394), .Y(n63407) );
  XNOR2X1 U67363 ( .A(n63407), .B(n43693), .Y(n63395) );
  XNOR2X1 U67364 ( .A(n63410), .B(n63395), .Y(n63402) );
  XNOR2X1 U67365 ( .A(n63402), .B(n43708), .Y(n63396) );
  XNOR2X1 U67366 ( .A(n41494), .B(n63396), .Y(n63401) );
  XNOR2X1 U67367 ( .A(n63398), .B(n63397), .Y(n63399) );
  XNOR2X1 U67368 ( .A(n41876), .B(n63399), .Y(n63400) );
  MX2X1 U67369 ( .A(n63401), .B(n63400), .S0(n43720), .Y(u_muldiv_result_r[3])
         );
  NAND2X1 U67370 ( .A(u_muldiv_mult_result_q[3]), .B(n44631), .Y(n14111) );
  NAND2X1 U67371 ( .A(n43706), .B(n63402), .Y(n63406) );
  INVX1 U67372 ( .A(n63402), .Y(n63403) );
  NAND2X1 U67373 ( .A(n63403), .B(n43713), .Y(n63404) );
  NAND2X1 U67374 ( .A(n41494), .B(n63404), .Y(n63405) );
  NAND2X1 U67375 ( .A(n63406), .B(n63405), .Y(n63952) );
  NAND2X1 U67376 ( .A(n63407), .B(n43700), .Y(n63412) );
  INVX1 U67377 ( .A(n63407), .Y(n63408) );
  NAND2X1 U67378 ( .A(n43694), .B(n63408), .Y(n63409) );
  NAND2X1 U67379 ( .A(n63410), .B(n63409), .Y(n63411) );
  INVX1 U67380 ( .A(n63414), .Y(n63413) );
  NAND2X1 U67381 ( .A(n43506), .B(n63413), .Y(n63418) );
  NAND2X1 U67382 ( .A(n63414), .B(n43513), .Y(n63415) );
  NAND2X1 U67383 ( .A(n63416), .B(n63415), .Y(n63417) );
  AND2X1 U67384 ( .A(n63418), .B(n63417), .Y(n63940) );
  INVX1 U67385 ( .A(n63419), .Y(n63420) );
  NAND2X1 U67386 ( .A(n63420), .B(n43688), .Y(n63422) );
  NAND2X1 U67387 ( .A(n38665), .B(n63425), .Y(n63426) );
  INVX1 U67388 ( .A(n63702), .Y(n63705) );
  NAND2X1 U67389 ( .A(n43791), .B(n44049), .Y(n63709) );
  INVX1 U67390 ( .A(n63428), .Y(n63427) );
  NAND2X1 U67391 ( .A(n38852), .B(n63428), .Y(n63429) );
  NAND2X1 U67392 ( .A(n63434), .B(n63430), .Y(n63437) );
  NAND2X1 U67393 ( .A(n63432), .B(n63431), .Y(n63433) );
  OR2X1 U67394 ( .A(n63434), .B(n63433), .Y(n63435) );
  NAND2X1 U67395 ( .A(n42078), .B(n63435), .Y(n63436) );
  NAND2X1 U67396 ( .A(n63437), .B(n63436), .Y(n63715) );
  NAND2X1 U67397 ( .A(n43779), .B(n44026), .Y(n63713) );
  INVX1 U67398 ( .A(n63438), .Y(n63676) );
  XNOR2X1 U67399 ( .A(n63675), .B(n63676), .Y(n63439) );
  INVX1 U67400 ( .A(n63450), .Y(n63440) );
  NAND2X1 U67401 ( .A(n63441), .B(n63440), .Y(n63718) );
  NAND2X1 U67402 ( .A(n63445), .B(n63444), .Y(n63446) );
  NOR2X1 U67403 ( .A(n63447), .B(n63446), .Y(n63448) );
  NOR2X1 U67404 ( .A(n44005), .B(n63448), .Y(n63449) );
  NOR2X1 U67405 ( .A(n39986), .B(n63449), .Y(n63451) );
  NAND2X1 U67406 ( .A(n63718), .B(n63719), .Y(n63721) );
  NAND2X1 U67407 ( .A(n43735), .B(n44018), .Y(n63717) );
  NOR2X1 U67408 ( .A(n63452), .B(n63920), .Y(n63454) );
  NAND2X1 U67409 ( .A(n63456), .B(n63455), .Y(n63457) );
  NAND2X1 U67410 ( .A(n63457), .B(n43974), .Y(n63459) );
  NAND2X1 U67411 ( .A(n63459), .B(n63458), .Y(n63918) );
  NAND2X1 U67412 ( .A(n43809), .B(n43993), .Y(n63996) );
  NAND2X1 U67413 ( .A(n40461), .B(n43984), .Y(n63901) );
  NAND2X1 U67414 ( .A(n63462), .B(n63461), .Y(n63897) );
  NAND2X1 U67415 ( .A(n63897), .B(n63898), .Y(n63896) );
  INVX1 U67416 ( .A(n63463), .Y(n63472) );
  NOR2X1 U67417 ( .A(n39881), .B(n63464), .Y(n63466) );
  NOR2X1 U67418 ( .A(n43930), .B(n63464), .Y(n63465) );
  NOR2X1 U67419 ( .A(n63465), .B(n63466), .Y(n63469) );
  NAND2X1 U67420 ( .A(n63467), .B(n43929), .Y(n63468) );
  NAND2X1 U67421 ( .A(n63469), .B(n63468), .Y(n63470) );
  XNOR2X1 U67422 ( .A(n63646), .B(n63650), .Y(n63471) );
  XOR2X1 U67423 ( .A(n63649), .B(n63471), .Y(n63473) );
  NOR2X1 U67424 ( .A(n41353), .B(n41457), .Y(n63475) );
  NAND2X1 U67425 ( .A(n63474), .B(n63473), .Y(n63741) );
  NAND2X1 U67426 ( .A(n63475), .B(n63741), .Y(n63739) );
  XNOR2X1 U67427 ( .A(n39636), .B(n41998), .Y(n63654) );
  XNOR2X1 U67428 ( .A(n42842), .B(n63476), .Y(n63480) );
  NOR2X1 U67429 ( .A(n63480), .B(n63477), .Y(n63478) );
  NOR2X1 U67430 ( .A(n63479), .B(n63478), .Y(n63484) );
  INVX1 U67431 ( .A(n63480), .Y(n63482) );
  NAND2X1 U67432 ( .A(n63482), .B(n63481), .Y(n63483) );
  NAND2X1 U67433 ( .A(n63484), .B(n63483), .Y(n63876) );
  NAND2X1 U67434 ( .A(n43798), .B(n43904), .Y(n63752) );
  INVX1 U67435 ( .A(n63485), .Y(n63488) );
  NAND2X1 U67436 ( .A(n63488), .B(n63486), .Y(n64208) );
  NOR2X1 U67437 ( .A(n63488), .B(n39347), .Y(n63490) );
  NAND2X1 U67438 ( .A(n63490), .B(n63489), .Y(n63492) );
  NAND2X1 U67439 ( .A(n63492), .B(n63491), .Y(n64207) );
  NAND2X1 U67440 ( .A(n64208), .B(n64207), .Y(n63760) );
  INVX1 U67441 ( .A(n63760), .Y(n63758) );
  NOR2X1 U67442 ( .A(n40064), .B(n63497), .Y(n63496) );
  INVX1 U67443 ( .A(n63498), .Y(n63494) );
  NOR2X1 U67444 ( .A(n40064), .B(n63494), .Y(n63495) );
  NOR2X1 U67445 ( .A(n63496), .B(n63495), .Y(n63501) );
  INVX1 U67446 ( .A(n63497), .Y(n63499) );
  NAND2X1 U67447 ( .A(n63499), .B(n63498), .Y(n63500) );
  NAND2X1 U67448 ( .A(n63501), .B(n63500), .Y(n63765) );
  NAND2X1 U67449 ( .A(n63774), .B(n39705), .Y(n63503) );
  NAND2X1 U67450 ( .A(n63503), .B(n63772), .Y(n63506) );
  INVX1 U67451 ( .A(n63506), .Y(n63504) );
  NOR2X1 U67452 ( .A(n63504), .B(n63773), .Y(n63505) );
  NOR2X1 U67453 ( .A(n41391), .B(n63505), .Y(n63508) );
  NAND2X1 U67454 ( .A(n63507), .B(n63506), .Y(n63770) );
  NAND2X1 U67455 ( .A(n63508), .B(n63770), .Y(n63866) );
  INVX1 U67456 ( .A(n63509), .Y(n63510) );
  NOR2X1 U67457 ( .A(n41198), .B(n41202), .Y(n63513) );
  NAND2X1 U67458 ( .A(n63512), .B(n63511), .Y(n63792) );
  NAND2X1 U67459 ( .A(n63513), .B(n63792), .Y(n63865) );
  INVX1 U67460 ( .A(n63514), .Y(n63517) );
  NOR2X1 U67461 ( .A(n41190), .B(n41189), .Y(n63518) );
  NAND2X1 U67462 ( .A(n63517), .B(n63516), .Y(n63797) );
  NAND2X1 U67463 ( .A(n63518), .B(n63797), .Y(n63804) );
  INVX1 U67464 ( .A(n63804), .Y(n63782) );
  NAND2X1 U67465 ( .A(n43870), .B(n43775), .Y(n63788) );
  XNOR2X1 U67466 ( .A(n63788), .B(n41689), .Y(n63520) );
  NAND2X1 U67467 ( .A(n43860), .B(n38310), .Y(n64159) );
  INVX1 U67468 ( .A(n64159), .Y(n64168) );
  XNOR2X1 U67469 ( .A(n64168), .B(n41688), .Y(n63790) );
  INVX1 U67470 ( .A(n63790), .Y(n63519) );
  XNOR2X1 U67471 ( .A(n63520), .B(n63519), .Y(n63584) );
  NAND2X1 U67472 ( .A(n43492), .B(n43851), .Y(n64148) );
  NOR2X1 U67473 ( .A(n38565), .B(n63525), .Y(n63522) );
  NOR2X1 U67474 ( .A(n63523), .B(n63522), .Y(n63527) );
  OR2X1 U67475 ( .A(n63525), .B(n63524), .Y(n63526) );
  XNOR2X1 U67476 ( .A(n64148), .B(n40469), .Y(n63578) );
  INVX1 U67477 ( .A(n63531), .Y(n63528) );
  NAND2X1 U67478 ( .A(n63529), .B(n63528), .Y(n63539) );
  NAND2X1 U67479 ( .A(n63531), .B(n63530), .Y(n63537) );
  NAND2X1 U67480 ( .A(n63533), .B(n63532), .Y(n63535) );
  NAND2X1 U67481 ( .A(n63535), .B(n63534), .Y(n63536) );
  NAND2X1 U67482 ( .A(n63537), .B(n63536), .Y(n63538) );
  NAND2X1 U67483 ( .A(n63539), .B(n63538), .Y(n63848) );
  NAND2X1 U67484 ( .A(n44035), .B(n43496), .Y(n63846) );
  INVX1 U67485 ( .A(n63846), .Y(n63845) );
  XNOR2X1 U67486 ( .A(n63848), .B(n63845), .Y(n63577) );
  INVX1 U67487 ( .A(n63544), .Y(n63540) );
  NAND2X1 U67488 ( .A(n63540), .B(n63543), .Y(n63542) );
  NAND2X1 U67489 ( .A(n63542), .B(n63541), .Y(n63807) );
  INVX1 U67490 ( .A(n63543), .Y(n63545) );
  NAND2X1 U67491 ( .A(n63545), .B(n63544), .Y(n63808) );
  NAND2X1 U67492 ( .A(n63808), .B(n63807), .Y(n63576) );
  INVX1 U67493 ( .A(n63565), .Y(n63557) );
  XNOR2X1 U67494 ( .A(n63571), .B(n63557), .Y(n64102) );
  INVX1 U67495 ( .A(n63549), .Y(n63546) );
  NAND2X1 U67496 ( .A(n63547), .B(n63546), .Y(n64069) );
  NAND2X1 U67497 ( .A(n63549), .B(n63548), .Y(n63813) );
  NAND2X1 U67498 ( .A(n64069), .B(n64070), .Y(n63811) );
  NAND2X1 U67499 ( .A(n43840), .B(n39961), .Y(n64109) );
  INVX1 U67500 ( .A(n64109), .Y(n64112) );
  NAND2X1 U67501 ( .A(n63835), .B(n63550), .Y(n63551) );
  NAND2X1 U67502 ( .A(n39082), .B(n63552), .Y(n63554) );
  NAND2X1 U67503 ( .A(n42162), .B(n38610), .Y(n63553) );
  NAND2X1 U67504 ( .A(n63554), .B(n63553), .Y(n63561) );
  NAND2X1 U67505 ( .A(n42162), .B(n63563), .Y(n63559) );
  NAND2X1 U67506 ( .A(n42162), .B(n63557), .Y(n63558) );
  NAND2X1 U67507 ( .A(n63559), .B(n63558), .Y(n63560) );
  NOR2X1 U67508 ( .A(n63561), .B(n63560), .Y(n63568) );
  NAND2X1 U67509 ( .A(n39082), .B(n63562), .Y(n63564) );
  NOR2X1 U67510 ( .A(n63564), .B(n63563), .Y(n63566) );
  NAND2X1 U67511 ( .A(n63566), .B(n63565), .Y(n63567) );
  XNOR2X1 U67512 ( .A(n64112), .B(n42161), .Y(n63573) );
  NOR2X1 U67513 ( .A(n43611), .B(n63569), .Y(n63570) );
  NAND2X1 U67514 ( .A(n63570), .B(n43603), .Y(n63828) );
  INVX1 U67515 ( .A(n63828), .Y(n64101) );
  NAND2X1 U67516 ( .A(n63571), .B(n38500), .Y(n63572) );
  XNOR2X1 U67517 ( .A(n63573), .B(n63818), .Y(n63574) );
  NAND2X1 U67518 ( .A(n38383), .B(n43502), .Y(n64121) );
  XNOR2X1 U67519 ( .A(n63809), .B(n64121), .Y(n63575) );
  XNOR2X1 U67520 ( .A(n63576), .B(n63575), .Y(n63847) );
  INVX1 U67521 ( .A(n63847), .Y(n63844) );
  XNOR2X1 U67522 ( .A(n63578), .B(n36777), .Y(n64165) );
  INVX1 U67523 ( .A(n63579), .Y(n63580) );
  NOR2X1 U67524 ( .A(n40992), .B(n40988), .Y(n63583) );
  NAND2X1 U67525 ( .A(n63582), .B(n63581), .Y(n63851) );
  XNOR2X1 U67526 ( .A(n63584), .B(n40946), .Y(n63585) );
  XNOR2X1 U67527 ( .A(n63782), .B(n63585), .Y(n63864) );
  NAND2X1 U67528 ( .A(n43879), .B(n43796), .Y(n64190) );
  INVX1 U67529 ( .A(n64190), .Y(n63586) );
  XNOR2X1 U67530 ( .A(n63864), .B(n63586), .Y(n63587) );
  XNOR2X1 U67531 ( .A(n63865), .B(n63587), .Y(n63588) );
  NAND2X1 U67532 ( .A(n43889), .B(n42712), .Y(n63764) );
  NOR2X1 U67533 ( .A(n63590), .B(n63593), .Y(n63592) );
  INVX1 U67534 ( .A(n63594), .Y(n63589) );
  NOR2X1 U67535 ( .A(n63590), .B(n63589), .Y(n63591) );
  INVX1 U67536 ( .A(n63593), .Y(n63595) );
  XNOR2X1 U67537 ( .A(n63764), .B(n64192), .Y(n63596) );
  NAND2X1 U67538 ( .A(n42651), .B(n43898), .Y(n63757) );
  INVX1 U67539 ( .A(n63757), .Y(n64204) );
  XNOR2X1 U67540 ( .A(n64205), .B(n64204), .Y(n63597) );
  XNOR2X1 U67541 ( .A(n63758), .B(n63597), .Y(n63755) );
  INVX1 U67542 ( .A(n63755), .Y(n63751) );
  XNOR2X1 U67543 ( .A(n63752), .B(n63751), .Y(n63606) );
  INVX1 U67544 ( .A(n63603), .Y(n63598) );
  NOR2X1 U67545 ( .A(n63598), .B(n63599), .Y(n63601) );
  NOR2X1 U67546 ( .A(n63601), .B(n63600), .Y(n63605) );
  NAND2X1 U67547 ( .A(n63604), .B(n63605), .Y(n63756) );
  XNOR2X1 U67548 ( .A(n63606), .B(n36739), .Y(n63875) );
  NAND2X1 U67549 ( .A(n37412), .B(n63609), .Y(n63886) );
  NAND2X1 U67550 ( .A(n43918), .B(n42641), .Y(n63882) );
  NAND2X1 U67551 ( .A(n63886), .B(n63882), .Y(n63610) );
  NOR2X1 U67552 ( .A(n39793), .B(n63610), .Y(n63624) );
  OR2X1 U67553 ( .A(n63882), .B(n63886), .Y(n63622) );
  NOR2X1 U67554 ( .A(n63611), .B(n63882), .Y(n63613) );
  NAND2X1 U67555 ( .A(n63613), .B(n63612), .Y(n63618) );
  NOR2X1 U67556 ( .A(n63614), .B(n63882), .Y(n63616) );
  NAND2X1 U67557 ( .A(n63616), .B(n63615), .Y(n63617) );
  NAND2X1 U67558 ( .A(n63618), .B(n63617), .Y(n63620) );
  NAND2X1 U67559 ( .A(n63620), .B(n63619), .Y(n63621) );
  NAND2X1 U67560 ( .A(n63622), .B(n63621), .Y(n63623) );
  NOR2X1 U67561 ( .A(n63623), .B(n63624), .Y(n63625) );
  XOR2X1 U67562 ( .A(n63888), .B(n63625), .Y(n64030) );
  NOR2X1 U67563 ( .A(n41922), .B(n63626), .Y(n63631) );
  INVX1 U67564 ( .A(n63627), .Y(n63628) );
  NOR2X1 U67565 ( .A(n39008), .B(n63628), .Y(n63630) );
  XNOR2X1 U67566 ( .A(n63632), .B(n37412), .Y(n63634) );
  XNOR2X1 U67567 ( .A(n63634), .B(n63633), .Y(n63635) );
  XNOR2X1 U67568 ( .A(n63636), .B(n63635), .Y(n63638) );
  OR2X1 U67569 ( .A(n63638), .B(n63637), .Y(n63639) );
  NAND2X1 U67570 ( .A(n63640), .B(n63639), .Y(n63749) );
  NAND2X1 U67571 ( .A(n43927), .B(n43724), .Y(n63746) );
  XNOR2X1 U67572 ( .A(n63749), .B(n63746), .Y(n63641) );
  XOR2X1 U67573 ( .A(n64030), .B(n63641), .Y(n63743) );
  XNOR2X1 U67574 ( .A(n41967), .B(n37318), .Y(n63653) );
  NOR2X1 U67575 ( .A(n43923), .B(n63642), .Y(n63645) );
  NOR2X1 U67576 ( .A(n36697), .B(n43921), .Y(n63643) );
  NOR2X1 U67577 ( .A(n63643), .B(n41259), .Y(n63644) );
  NAND2X1 U67578 ( .A(n63650), .B(n63649), .Y(n63651) );
  INVX1 U67579 ( .A(n40533), .Y(n63652) );
  XNOR2X1 U67580 ( .A(n63654), .B(n41644), .Y(n63655) );
  XNOR2X1 U67581 ( .A(n36487), .B(n63655), .Y(n63913) );
  NOR2X1 U67582 ( .A(n63656), .B(n63657), .Y(n63662) );
  INVX1 U67583 ( .A(n63657), .Y(n63907) );
  NAND2X1 U67584 ( .A(n63907), .B(n63658), .Y(n63660) );
  NAND2X1 U67585 ( .A(n63659), .B(n63658), .Y(n63910) );
  NAND2X1 U67586 ( .A(n63660), .B(n63910), .Y(n63661) );
  NOR2X1 U67587 ( .A(n63662), .B(n63661), .Y(n63663) );
  XNOR2X1 U67588 ( .A(n63664), .B(n63663), .Y(n64001) );
  INVX1 U67589 ( .A(n64001), .Y(n63916) );
  XNOR2X1 U67590 ( .A(n63996), .B(n63916), .Y(n63665) );
  NAND2X1 U67591 ( .A(n43820), .B(n44001), .Y(n63736) );
  INVX1 U67592 ( .A(n63668), .Y(n63666) );
  NAND2X1 U67593 ( .A(n63667), .B(n63666), .Y(n63733) );
  NAND2X1 U67594 ( .A(n63733), .B(n63732), .Y(n63731) );
  NAND2X1 U67595 ( .A(n43758), .B(n44009), .Y(n63724) );
  NAND2X1 U67596 ( .A(n63675), .B(n63671), .Y(n63725) );
  NAND2X1 U67597 ( .A(n63725), .B(n63726), .Y(n63730) );
  XNOR2X1 U67598 ( .A(n63717), .B(n63722), .Y(n63677) );
  INVX1 U67599 ( .A(n63980), .Y(n63716) );
  XNOR2X1 U67600 ( .A(n63713), .B(n63716), .Y(n63678) );
  XNOR2X1 U67601 ( .A(n39162), .B(n63678), .Y(n63712) );
  XNOR2X1 U67602 ( .A(n63711), .B(n63712), .Y(n63679) );
  XNOR2X1 U67603 ( .A(n63704), .B(n42111), .Y(n63680) );
  XNOR2X1 U67604 ( .A(n63705), .B(n63680), .Y(n63930) );
  INVX1 U67605 ( .A(n63930), .Y(n63931) );
  INVX1 U67606 ( .A(n63683), .Y(n63682) );
  NAND2X1 U67607 ( .A(n63682), .B(n63681), .Y(n63686) );
  NAND2X1 U67608 ( .A(n63686), .B(n63685), .Y(n63932) );
  NAND2X1 U67609 ( .A(n43612), .B(n43766), .Y(n72139) );
  XNOR2X1 U67610 ( .A(n63932), .B(n43524), .Y(n63687) );
  XNOR2X1 U67611 ( .A(n63931), .B(n63687), .Y(n63697) );
  XNOR2X1 U67612 ( .A(n63938), .B(n43508), .Y(n63688) );
  XNOR2X1 U67613 ( .A(n63940), .B(n63688), .Y(n63945) );
  XNOR2X1 U67614 ( .A(n63945), .B(n43694), .Y(n63689) );
  XNOR2X1 U67615 ( .A(n41484), .B(n63689), .Y(n63951) );
  XNOR2X1 U67616 ( .A(n63951), .B(n43708), .Y(n63690) );
  XNOR2X1 U67617 ( .A(n37904), .B(n63690), .Y(n63695) );
  XNOR2X1 U67618 ( .A(n63692), .B(n63691), .Y(n63693) );
  XNOR2X1 U67619 ( .A(n63693), .B(n41887), .Y(n63694) );
  MX2X1 U67620 ( .A(n63695), .B(n63694), .S0(n43720), .Y(u_muldiv_result_r[4])
         );
  NAND2X1 U67621 ( .A(u_muldiv_mult_result_q[4]), .B(n44633), .Y(n14103) );
  INVX1 U67622 ( .A(n63697), .Y(n63696) );
  NAND2X1 U67623 ( .A(n43676), .B(n63696), .Y(n63701) );
  NAND2X1 U67624 ( .A(n63697), .B(n43686), .Y(n63699) );
  NAND2X1 U67625 ( .A(n63699), .B(n63698), .Y(n63700) );
  NAND2X1 U67626 ( .A(n63701), .B(n63700), .Y(n63971) );
  INVX1 U67627 ( .A(n63704), .Y(n63703) );
  NAND2X1 U67628 ( .A(n63703), .B(n63702), .Y(n63708) );
  NAND2X1 U67629 ( .A(n42111), .B(n63706), .Y(n63707) );
  AND2X1 U67630 ( .A(n63708), .B(n63707), .Y(n64265) );
  NOR2X1 U67631 ( .A(n63712), .B(n63711), .Y(n63710) );
  OR2X1 U67632 ( .A(n63710), .B(n63709), .Y(n64254) );
  NAND2X1 U67633 ( .A(n63712), .B(n63711), .Y(n64257) );
  NAND2X1 U67634 ( .A(n64254), .B(n64257), .Y(n63928) );
  NAND2X1 U67635 ( .A(n43791), .B(n44056), .Y(n64253) );
  INVX1 U67636 ( .A(n63713), .Y(n63981) );
  NAND2X1 U67637 ( .A(n39162), .B(n63980), .Y(n63714) );
  INVX1 U67638 ( .A(n63717), .Y(n63720) );
  NAND2X1 U67639 ( .A(n63720), .B(n63987), .Y(n63723) );
  XNOR2X1 U67640 ( .A(n37360), .B(n42088), .Y(n63926) );
  INVX1 U67641 ( .A(n63724), .Y(n63727) );
  INVX1 U67642 ( .A(n63728), .Y(n63729) );
  NOR2X1 U67643 ( .A(n63734), .B(n63736), .Y(n63735) );
  INVX1 U67644 ( .A(n63736), .Y(n63737) );
  NAND2X1 U67645 ( .A(n43820), .B(n44009), .Y(n63989) );
  XNOR2X1 U67646 ( .A(n40533), .B(n41967), .Y(n63738) );
  XNOR2X1 U67647 ( .A(n63743), .B(n63738), .Y(n63740) );
  NAND2X1 U67648 ( .A(n63740), .B(n63739), .Y(n64020) );
  NAND2X1 U67649 ( .A(n39185), .B(n37318), .Y(n63742) );
  NAND2X1 U67650 ( .A(n64020), .B(n63742), .Y(n63895) );
  NOR2X1 U67651 ( .A(n41575), .B(n41537), .Y(n63745) );
  NAND2X1 U67652 ( .A(n40533), .B(n63743), .Y(n64016) );
  NAND2X1 U67653 ( .A(n63745), .B(n64016), .Y(n64029) );
  INVX1 U67654 ( .A(n64029), .Y(n63893) );
  NAND2X1 U67655 ( .A(n43724), .B(n43934), .Y(n64038) );
  NOR2X1 U67656 ( .A(n40217), .B(n63746), .Y(n63747) );
  NOR2X1 U67657 ( .A(n63748), .B(n63747), .Y(n63750) );
  NAND2X1 U67658 ( .A(n64030), .B(n63749), .Y(n64031) );
  NOR2X1 U67659 ( .A(n63751), .B(n63752), .Y(n63754) );
  NOR2X1 U67660 ( .A(n36739), .B(n63752), .Y(n63753) );
  INVX1 U67661 ( .A(n64205), .Y(n63761) );
  NOR2X1 U67662 ( .A(n63758), .B(n63757), .Y(n63759) );
  NAND2X1 U67663 ( .A(n42652), .B(n43904), .Y(n64209) );
  XNOR2X1 U67664 ( .A(n64209), .B(n41709), .Y(n63769) );
  NAND2X1 U67665 ( .A(n41343), .B(n63763), .Y(n63768) );
  NAND2X1 U67666 ( .A(n63766), .B(n63765), .Y(n63767) );
  NAND2X1 U67667 ( .A(n63768), .B(n63767), .Y(n64051) );
  XNOR2X1 U67668 ( .A(n63769), .B(n36726), .Y(n63870) );
  NAND2X1 U67669 ( .A(n43889), .B(n43796), .Y(n64188) );
  INVX1 U67670 ( .A(n63770), .Y(n63771) );
  NOR2X1 U67671 ( .A(n41391), .B(n63771), .Y(n63780) );
  NOR2X1 U67672 ( .A(n63773), .B(n63772), .Y(n63778) );
  NOR2X1 U67673 ( .A(n39768), .B(n63773), .Y(n63775) );
  NAND2X1 U67674 ( .A(n63775), .B(n63774), .Y(n63776) );
  NAND2X1 U67675 ( .A(n63776), .B(n63788), .Y(n63777) );
  NOR2X1 U67676 ( .A(n63778), .B(n63777), .Y(n63779) );
  NAND2X1 U67677 ( .A(n63780), .B(n63779), .Y(n63787) );
  INVX1 U67678 ( .A(n63865), .Y(n63785) );
  XNOR2X1 U67679 ( .A(n63790), .B(n41689), .Y(n63781) );
  XNOR2X1 U67680 ( .A(n40946), .B(n63781), .Y(n63783) );
  XNOR2X1 U67681 ( .A(n63783), .B(n63782), .Y(n63784) );
  XNOR2X1 U67682 ( .A(n63785), .B(n63784), .Y(n63786) );
  NAND2X1 U67683 ( .A(n63787), .B(n63786), .Y(n64179) );
  INVX1 U67684 ( .A(n63788), .Y(n63789) );
  NAND2X1 U67685 ( .A(n63789), .B(n63866), .Y(n64180) );
  NAND2X1 U67686 ( .A(n64179), .B(n64180), .Y(n64372) );
  XNOR2X1 U67687 ( .A(n63790), .B(n40948), .Y(n63791) );
  NOR2X1 U67688 ( .A(n41198), .B(n41202), .Y(n63793) );
  NAND2X1 U67689 ( .A(n63793), .B(n63792), .Y(n63795) );
  NOR2X1 U67690 ( .A(n41456), .B(n40991), .Y(n63796) );
  NAND2X1 U67691 ( .A(n41689), .B(n63795), .Y(n64055) );
  NAND2X1 U67692 ( .A(n63796), .B(n64055), .Y(n64181) );
  NOR2X1 U67693 ( .A(n41189), .B(n41688), .Y(n63800) );
  INVX1 U67694 ( .A(n63797), .Y(n63798) );
  NOR2X1 U67695 ( .A(n41190), .B(n63798), .Y(n63799) );
  NAND2X1 U67696 ( .A(n63800), .B(n63799), .Y(n63803) );
  XNOR2X1 U67697 ( .A(n64159), .B(n38619), .Y(n63801) );
  XNOR2X1 U67698 ( .A(n40948), .B(n63801), .Y(n63802) );
  NAND2X1 U67699 ( .A(n63803), .B(n63802), .Y(n63806) );
  NAND2X1 U67700 ( .A(n41688), .B(n63804), .Y(n63805) );
  NAND2X1 U67701 ( .A(n63806), .B(n63805), .Y(n64177) );
  INVX1 U67702 ( .A(n64148), .Y(n64149) );
  INVX1 U67703 ( .A(n64121), .Y(n64426) );
  NAND2X1 U67704 ( .A(n63808), .B(n63807), .Y(n63810) );
  INVX1 U67705 ( .A(n63809), .Y(n64120) );
  NAND2X1 U67706 ( .A(n64419), .B(n64427), .Y(n63843) );
  XNOR2X1 U67707 ( .A(n63818), .B(n42161), .Y(n64110) );
  INVX1 U67708 ( .A(n64110), .Y(n64072) );
  NAND2X1 U67709 ( .A(n63813), .B(n63812), .Y(n64070) );
  NAND2X1 U67710 ( .A(n64070), .B(n64069), .Y(n64111) );
  INVX1 U67711 ( .A(n64111), .Y(n63814) );
  NAND2X1 U67712 ( .A(n63814), .B(n64110), .Y(n63815) );
  INVX1 U67713 ( .A(n65067), .Y(n64133) );
  NAND2X1 U67714 ( .A(n38500), .B(n63816), .Y(n63817) );
  NOR2X1 U67715 ( .A(n42166), .B(n64102), .Y(n63819) );
  NAND2X1 U67716 ( .A(n63819), .B(n63818), .Y(n64065) );
  NAND2X1 U67717 ( .A(n39082), .B(n64065), .Y(n64129) );
  NAND2X1 U67718 ( .A(n43850), .B(n43497), .Y(n64140) );
  INVX1 U67719 ( .A(n64140), .Y(n63820) );
  NAND2X1 U67720 ( .A(n44035), .B(n43502), .Y(n64431) );
  INVX1 U67721 ( .A(n64431), .Y(n64126) );
  XNOR2X1 U67722 ( .A(n63820), .B(n64126), .Y(n63840) );
  NAND2X1 U67723 ( .A(n36781), .B(n63821), .Y(n63822) );
  NOR2X1 U67724 ( .A(n62452), .B(n64087), .Y(n63827) );
  NAND2X1 U67725 ( .A(n63827), .B(n63826), .Y(n63829) );
  NAND2X1 U67726 ( .A(n63829), .B(n63828), .Y(n64089) );
  INVX1 U67727 ( .A(n64089), .Y(n63832) );
  INVX1 U67728 ( .A(n63196), .Y(n63831) );
  NAND2X1 U67729 ( .A(n63831), .B(n63830), .Y(n64090) );
  NAND2X1 U67730 ( .A(n38297), .B(n38500), .Y(n64079) );
  NOR2X1 U67731 ( .A(n63834), .B(n63833), .Y(n63838) );
  NAND2X1 U67732 ( .A(n63835), .B(n42799), .Y(n63836) );
  NAND2X1 U67733 ( .A(n43603), .B(n63836), .Y(n63837) );
  NOR2X1 U67734 ( .A(n63838), .B(n63837), .Y(n63839) );
  NAND2X1 U67735 ( .A(n43840), .B(n43608), .Y(n64064) );
  NAND2X1 U67736 ( .A(n38379), .B(n43518), .Y(n64413) );
  XNOR2X1 U67737 ( .A(n63840), .B(n64130), .Y(n63841) );
  XNOR2X1 U67738 ( .A(n64129), .B(n63841), .Y(n63842) );
  XNOR2X1 U67739 ( .A(n64133), .B(n63842), .Y(n64060) );
  NAND2X1 U67740 ( .A(n43492), .B(n43861), .Y(n64062) );
  NAND2X1 U67741 ( .A(n63845), .B(n63844), .Y(n64136) );
  NAND2X1 U67742 ( .A(n63847), .B(n63846), .Y(n63849) );
  NAND2X1 U67743 ( .A(n63849), .B(n63848), .Y(n64137) );
  NAND2X1 U67744 ( .A(n64136), .B(n64137), .Y(n64146) );
  NAND2X1 U67745 ( .A(n43962), .B(n43486), .Y(n64380) );
  XNOR2X1 U67746 ( .A(n64146), .B(n64380), .Y(n63850) );
  NAND2X1 U67747 ( .A(n63583), .B(n63851), .Y(n64167) );
  INVX1 U67748 ( .A(n64167), .Y(n64166) );
  NAND2X1 U67749 ( .A(n64159), .B(n64165), .Y(n63856) );
  INVX1 U67750 ( .A(n63856), .Y(n63852) );
  NOR2X1 U67751 ( .A(n64166), .B(n63852), .Y(n63854) );
  NAND2X1 U67752 ( .A(n43952), .B(n43482), .Y(n64175) );
  NAND2X1 U67753 ( .A(n38880), .B(n64175), .Y(n63853) );
  NOR2X1 U67754 ( .A(n63854), .B(n63853), .Y(n63861) );
  NOR2X1 U67755 ( .A(n64159), .B(n64165), .Y(n63855) );
  INVX1 U67756 ( .A(n64175), .Y(n64174) );
  NAND2X1 U67757 ( .A(n63855), .B(n64174), .Y(n63859) );
  NOR2X1 U67758 ( .A(n64166), .B(n64175), .Y(n63857) );
  NAND2X1 U67759 ( .A(n63857), .B(n63856), .Y(n63858) );
  NAND2X1 U67760 ( .A(n63859), .B(n63858), .Y(n63860) );
  XNOR2X1 U67761 ( .A(n39483), .B(n64184), .Y(n64057) );
  INVX1 U67762 ( .A(n64057), .Y(n64054) );
  NAND2X1 U67763 ( .A(n43879), .B(n43775), .Y(n64375) );
  NAND2X1 U67764 ( .A(n43871), .B(n43478), .Y(n64182) );
  XNOR2X1 U67765 ( .A(n64375), .B(n64182), .Y(n63862) );
  XNOR2X1 U67766 ( .A(n64372), .B(n63863), .Y(n64197) );
  XNOR2X1 U67767 ( .A(n64188), .B(n64197), .Y(n63869) );
  NOR2X1 U67768 ( .A(n38524), .B(n64190), .Y(n63867) );
  INVX1 U67769 ( .A(n64191), .Y(n63868) );
  INVX1 U67770 ( .A(n64052), .Y(n64202) );
  NAND2X1 U67771 ( .A(n43798), .B(n43911), .Y(n64046) );
  INVX1 U67772 ( .A(n64046), .Y(n64050) );
  XNOR2X1 U67773 ( .A(n64045), .B(n64050), .Y(n63871) );
  XNOR2X1 U67774 ( .A(n39656), .B(n63871), .Y(n64226) );
  NAND2X1 U67775 ( .A(n43918), .B(n40259), .Y(n64041) );
  INVX1 U67776 ( .A(n64041), .Y(n64225) );
  XNOR2X1 U67777 ( .A(n41513), .B(n64225), .Y(n63880) );
  NOR2X1 U67778 ( .A(n63875), .B(n63872), .Y(n63873) );
  NOR2X1 U67779 ( .A(n63874), .B(n63873), .Y(n63879) );
  INVX1 U67780 ( .A(n63875), .Y(n63877) );
  NAND2X1 U67781 ( .A(n63877), .B(n40218), .Y(n63878) );
  XNOR2X1 U67782 ( .A(n63880), .B(n39758), .Y(n63881) );
  XNOR2X1 U67783 ( .A(n64226), .B(n63881), .Y(n63890) );
  INVX1 U67784 ( .A(n63882), .Y(n63885) );
  NAND2X1 U67785 ( .A(n63886), .B(n63883), .Y(n63884) );
  NAND2X1 U67786 ( .A(n63885), .B(n63884), .Y(n64222) );
  NOR2X1 U67787 ( .A(n39793), .B(n63885), .Y(n63887) );
  NAND2X1 U67788 ( .A(n63887), .B(n63886), .Y(n63889) );
  NAND2X1 U67789 ( .A(n63889), .B(n63888), .Y(n64223) );
  NAND2X1 U67790 ( .A(n64222), .B(n64223), .Y(n64221) );
  NAND2X1 U67791 ( .A(n43788), .B(n43943), .Y(n64018) );
  NAND2X1 U67792 ( .A(n40486), .B(n43973), .Y(n64024) );
  XNOR2X1 U67793 ( .A(n64018), .B(n64024), .Y(n63891) );
  XOR2X1 U67794 ( .A(n64028), .B(n63891), .Y(n63892) );
  XNOR2X1 U67795 ( .A(n63893), .B(n63892), .Y(n63894) );
  XNOR2X1 U67796 ( .A(n63895), .B(n63894), .Y(n64327) );
  NAND2X1 U67797 ( .A(n40475), .B(n43984), .Y(n64008) );
  XNOR2X1 U67798 ( .A(n39636), .B(n41644), .Y(n64009) );
  INVX1 U67799 ( .A(n64009), .Y(n64010) );
  INVX1 U67800 ( .A(n64009), .Y(n63900) );
  NAND2X1 U67801 ( .A(n63898), .B(n63897), .Y(n63899) );
  INVX1 U67802 ( .A(n63901), .Y(n63909) );
  NAND2X1 U67803 ( .A(n63903), .B(n63902), .Y(n63904) );
  NOR2X1 U67804 ( .A(n39757), .B(n63904), .Y(n63906) );
  NAND2X1 U67805 ( .A(n63910), .B(n63911), .Y(n63908) );
  OR2X1 U67806 ( .A(n63913), .B(n63908), .Y(n64235) );
  NAND2X1 U67807 ( .A(n63909), .B(n64235), .Y(n63914) );
  NAND2X1 U67808 ( .A(n63911), .B(n63910), .Y(n63912) );
  NAND2X1 U67809 ( .A(n63913), .B(n63912), .Y(n64236) );
  NAND2X1 U67810 ( .A(n64236), .B(n63914), .Y(n64239) );
  XNOR2X1 U67811 ( .A(n64239), .B(n42020), .Y(n63915) );
  XNOR2X1 U67812 ( .A(n64240), .B(n63915), .Y(n64311) );
  INVX1 U67813 ( .A(n64311), .Y(n63999) );
  XNOR2X1 U67814 ( .A(n63989), .B(n63999), .Y(n63925) );
  NAND2X1 U67815 ( .A(n43809), .B(n44001), .Y(n64645) );
  NAND2X1 U67816 ( .A(n63917), .B(n63916), .Y(n64644) );
  NOR2X1 U67817 ( .A(n63995), .B(n63996), .Y(n63921) );
  NOR2X1 U67818 ( .A(n40438), .B(n63921), .Y(n63923) );
  OR2X1 U67819 ( .A(n64001), .B(n63996), .Y(n63922) );
  NAND2X1 U67820 ( .A(n63923), .B(n63922), .Y(n64312) );
  XNOR2X1 U67821 ( .A(n40198), .B(n64645), .Y(n63924) );
  NAND2X1 U67822 ( .A(n43759), .B(n44018), .Y(n64296) );
  XNOR2X1 U67823 ( .A(n63926), .B(n41640), .Y(n63927) );
  NAND2X1 U67824 ( .A(n43612), .B(n38611), .Y(n72620) );
  XNOR2X1 U67825 ( .A(n64263), .B(n43654), .Y(n63929) );
  XNOR2X1 U67826 ( .A(n64265), .B(n63929), .Y(n63973) );
  INVX1 U67827 ( .A(n63973), .Y(n63975) );
  NAND2X1 U67828 ( .A(n43521), .B(n63930), .Y(n63935) );
  NAND2X1 U67829 ( .A(n63931), .B(n43527), .Y(n63933) );
  NAND2X1 U67830 ( .A(n63933), .B(n63932), .Y(n63934) );
  NAND2X1 U67831 ( .A(n63935), .B(n63934), .Y(n63974) );
  XNOR2X1 U67832 ( .A(n63974), .B(n43524), .Y(n63936) );
  XNOR2X1 U67833 ( .A(n63975), .B(n63936), .Y(n63969) );
  INVX1 U67834 ( .A(n64274), .Y(n64271) );
  INVX1 U67835 ( .A(n63938), .Y(n63937) );
  NAND2X1 U67836 ( .A(n63937), .B(n43514), .Y(n63942) );
  NAND2X1 U67837 ( .A(n43506), .B(n63938), .Y(n63939) );
  NAND2X1 U67838 ( .A(n63940), .B(n63939), .Y(n63941) );
  NAND2X1 U67839 ( .A(n63942), .B(n63941), .Y(n64272) );
  XNOR2X1 U67840 ( .A(n64272), .B(n43509), .Y(n63943) );
  XNOR2X1 U67841 ( .A(n64271), .B(n63943), .Y(n63962) );
  INVX1 U67842 ( .A(n63962), .Y(n63964) );
  INVX1 U67843 ( .A(n63945), .Y(n63944) );
  NAND2X1 U67844 ( .A(n43691), .B(n63944), .Y(n63948) );
  NAND2X1 U67845 ( .A(n63945), .B(n43701), .Y(n63946) );
  NAND2X1 U67846 ( .A(n41484), .B(n63946), .Y(n63947) );
  NAND2X1 U67847 ( .A(n63948), .B(n63947), .Y(n63963) );
  XNOR2X1 U67848 ( .A(n63963), .B(n43694), .Y(n63949) );
  XNOR2X1 U67849 ( .A(n63964), .B(n63949), .Y(n64276) );
  INVX1 U67850 ( .A(n64276), .Y(n64277) );
  XNOR2X1 U67851 ( .A(n43709), .B(n64277), .Y(n63956) );
  INVX1 U67852 ( .A(n63951), .Y(n63950) );
  NAND2X1 U67853 ( .A(n43707), .B(n63950), .Y(n63955) );
  NAND2X1 U67854 ( .A(n63951), .B(n43713), .Y(n63953) );
  NAND2X1 U67855 ( .A(n63953), .B(n63952), .Y(n63954) );
  NAND2X1 U67856 ( .A(n63955), .B(n63954), .Y(n64278) );
  XNOR2X1 U67857 ( .A(n63956), .B(n36357), .Y(n63961) );
  XNOR2X1 U67858 ( .A(n63958), .B(n63957), .Y(n63959) );
  XNOR2X1 U67859 ( .A(n41898), .B(n63959), .Y(n63960) );
  MX2X1 U67860 ( .A(n63961), .B(n63960), .S0(n43720), .Y(u_muldiv_result_r[5])
         );
  NAND2X1 U67861 ( .A(u_muldiv_mult_result_q[5]), .B(n44633), .Y(n14092) );
  NAND2X1 U67862 ( .A(n63962), .B(n43700), .Y(n63968) );
  INVX1 U67863 ( .A(n63963), .Y(n63966) );
  NAND2X1 U67864 ( .A(n43691), .B(n63964), .Y(n63965) );
  NAND2X1 U67865 ( .A(n63966), .B(n63965), .Y(n63967) );
  NAND2X1 U67866 ( .A(n63968), .B(n63967), .Y(n64555) );
  INVX1 U67867 ( .A(n63969), .Y(n63970) );
  NAND2X1 U67868 ( .A(n63970), .B(n43686), .Y(n63972) );
  NAND2X1 U67869 ( .A(n63973), .B(n43532), .Y(n63977) );
  NAND2X1 U67870 ( .A(n43521), .B(n63975), .Y(n63976) );
  XNOR2X1 U67871 ( .A(n37360), .B(n41640), .Y(n63979) );
  NAND2X1 U67872 ( .A(n63978), .B(n63979), .Y(n64520) );
  NOR2X1 U67873 ( .A(n37381), .B(n63979), .Y(n63983) );
  NAND2X1 U67874 ( .A(n63981), .B(n63714), .Y(n63982) );
  NAND2X1 U67875 ( .A(n63983), .B(n63982), .Y(n63984) );
  NAND2X1 U67876 ( .A(n42088), .B(n63984), .Y(n64521) );
  NAND2X1 U67877 ( .A(n64520), .B(n64521), .Y(n64525) );
  NAND2X1 U67878 ( .A(n43779), .B(n44056), .Y(n64519) );
  NAND2X1 U67879 ( .A(n63990), .B(n63988), .Y(n64507) );
  NOR2X1 U67880 ( .A(n41308), .B(n63990), .Y(n63994) );
  NAND2X1 U67881 ( .A(n44001), .B(n63992), .Y(n63993) );
  NAND2X1 U67882 ( .A(n64507), .B(n64508), .Y(n64510) );
  NAND2X1 U67883 ( .A(n43821), .B(n44018), .Y(n64506) );
  NOR2X1 U67884 ( .A(n41265), .B(n64000), .Y(n63995) );
  NOR2X1 U67885 ( .A(n41360), .B(n63996), .Y(n63997) );
  NOR2X1 U67886 ( .A(n40438), .B(n63997), .Y(n63998) );
  NOR2X1 U67887 ( .A(n63999), .B(n63998), .Y(n64007) );
  INVX1 U67888 ( .A(n64645), .Y(n64642) );
  NAND2X1 U67889 ( .A(n64642), .B(n64311), .Y(n64648) );
  NOR2X1 U67890 ( .A(n41265), .B(n64000), .Y(n64002) );
  NAND2X1 U67891 ( .A(n64002), .B(n64001), .Y(n64003) );
  NAND2X1 U67892 ( .A(n64003), .B(n43993), .Y(n64004) );
  NAND2X1 U67893 ( .A(n64004), .B(n64644), .Y(n64005) );
  NAND2X1 U67894 ( .A(n64642), .B(n64005), .Y(n64310) );
  NAND2X1 U67895 ( .A(n64648), .B(n64310), .Y(n64006) );
  NOR2X1 U67896 ( .A(n64007), .B(n64006), .Y(n64244) );
  NOR2X1 U67897 ( .A(n43977), .B(n64009), .Y(n64013) );
  NOR2X1 U67898 ( .A(n64010), .B(n43975), .Y(n64011) );
  NOR2X1 U67899 ( .A(n36487), .B(n64011), .Y(n64012) );
  NOR2X1 U67900 ( .A(n64013), .B(n64012), .Y(n64015) );
  INVX1 U67901 ( .A(n64327), .Y(n64014) );
  NAND2X1 U67902 ( .A(n64330), .B(n64329), .Y(n64317) );
  NOR2X1 U67903 ( .A(n41575), .B(n41537), .Y(n64017) );
  NAND2X1 U67904 ( .A(n64016), .B(n64017), .Y(n64026) );
  INVX1 U67905 ( .A(n64018), .Y(n64027) );
  XNOR2X1 U67906 ( .A(n64028), .B(n64027), .Y(n64019) );
  NAND2X1 U67907 ( .A(n64025), .B(n64024), .Y(n64023) );
  NAND2X1 U67908 ( .A(n64020), .B(n64021), .Y(n64022) );
  NAND2X1 U67909 ( .A(n64023), .B(n64022), .Y(n64859) );
  INVX1 U67910 ( .A(n64333), .Y(n64858) );
  NOR2X1 U67911 ( .A(n39913), .B(n64858), .Y(n64233) );
  XNOR2X1 U67912 ( .A(n39988), .B(n42004), .Y(n64231) );
  NOR2X1 U67913 ( .A(n43930), .B(n40217), .Y(n64034) );
  NAND2X1 U67914 ( .A(n64030), .B(n43929), .Y(n64032) );
  NAND2X1 U67915 ( .A(n64032), .B(n64031), .Y(n64033) );
  NOR2X1 U67916 ( .A(n64034), .B(n64033), .Y(n64035) );
  NOR2X1 U67917 ( .A(n64035), .B(n64038), .Y(n64037) );
  NOR2X1 U67918 ( .A(n64039), .B(n41566), .Y(n64036) );
  OR2X1 U67919 ( .A(n64039), .B(n64038), .Y(n64040) );
  NAND2X1 U67920 ( .A(n42632), .B(n43934), .Y(n64344) );
  NOR2X1 U67921 ( .A(n39758), .B(n64226), .Y(n64043) );
  NOR2X1 U67922 ( .A(n64226), .B(n64041), .Y(n64042) );
  NAND2X1 U67923 ( .A(n43927), .B(n43772), .Y(n64486) );
  INVX1 U67924 ( .A(n64045), .Y(n64047) );
  NOR2X1 U67925 ( .A(n64047), .B(n64046), .Y(n64049) );
  NOR2X1 U67926 ( .A(n64047), .B(n39656), .Y(n64048) );
  NAND2X1 U67927 ( .A(n42653), .B(n43911), .Y(n64361) );
  NOR2X1 U67928 ( .A(n41111), .B(n41372), .Y(n64053) );
  NAND2X1 U67929 ( .A(n41709), .B(n64052), .Y(n64366) );
  NAND2X1 U67930 ( .A(n64053), .B(n64366), .Y(n65122) );
  NOR2X1 U67931 ( .A(n41456), .B(n40991), .Y(n64056) );
  NAND2X1 U67932 ( .A(n64056), .B(n64055), .Y(n64059) );
  NAND2X1 U67933 ( .A(n64182), .B(n64057), .Y(n64058) );
  NAND2X1 U67934 ( .A(n64059), .B(n64058), .Y(n64466) );
  NAND2X1 U67935 ( .A(n64464), .B(n64466), .Y(n64463) );
  NAND2X1 U67936 ( .A(n43879), .B(n43478), .Y(n64462) );
  NAND2X1 U67937 ( .A(n43870), .B(n38312), .Y(n64455) );
  OR2X1 U67938 ( .A(n64063), .B(n64062), .Y(n64730) );
  NAND2X1 U67939 ( .A(n64729), .B(n64730), .Y(n64445) );
  NAND2X1 U67940 ( .A(n43492), .B(n43963), .Y(n64446) );
  INVX1 U67941 ( .A(n64064), .Y(n64106) );
  INVX1 U67942 ( .A(n64065), .Y(n64067) );
  NOR2X1 U67943 ( .A(n64067), .B(n64066), .Y(n64068) );
  XNOR2X1 U67944 ( .A(n41805), .B(n64068), .Y(n64415) );
  NAND2X1 U67945 ( .A(n64415), .B(n65067), .Y(n64078) );
  INVX1 U67946 ( .A(n64413), .Y(n64402) );
  NAND2X1 U67947 ( .A(n64070), .B(n64069), .Y(n64071) );
  NOR2X1 U67948 ( .A(n64072), .B(n64071), .Y(n64073) );
  NOR2X1 U67949 ( .A(n64073), .B(n64109), .Y(n64074) );
  NOR2X1 U67950 ( .A(n38293), .B(n64074), .Y(n64076) );
  INVX1 U67951 ( .A(n64415), .Y(n64075) );
  NAND2X1 U67952 ( .A(n64076), .B(n64075), .Y(n65047) );
  NAND2X1 U67953 ( .A(n64402), .B(n65047), .Y(n64077) );
  NAND2X1 U67954 ( .A(n64078), .B(n64077), .Y(n64795) );
  INVX1 U67955 ( .A(n64795), .Y(n64424) );
  OR2X1 U67956 ( .A(n64081), .B(n64080), .Y(n64085) );
  NAND2X1 U67957 ( .A(n64083), .B(n42798), .Y(n64084) );
  NAND2X1 U67958 ( .A(n64085), .B(n64084), .Y(n64086) );
  NOR2X1 U67959 ( .A(n64087), .B(n64086), .Y(n64088) );
  NAND2X1 U67960 ( .A(n64088), .B(n43608), .Y(n64773) );
  INVX1 U67961 ( .A(n64773), .Y(n64406) );
  XNOR2X1 U67962 ( .A(n42237), .B(n64406), .Y(n64094) );
  NAND2X1 U67963 ( .A(n41803), .B(n64094), .Y(n64098) );
  NOR2X1 U67964 ( .A(n38610), .B(n64089), .Y(n64091) );
  NAND2X1 U67965 ( .A(n64091), .B(n64090), .Y(n64093) );
  NOR2X1 U67966 ( .A(n64094), .B(n64093), .Y(n64092) );
  NOR2X1 U67967 ( .A(n64092), .B(n41803), .Y(n64096) );
  NAND2X1 U67968 ( .A(n64094), .B(n64093), .Y(n64095) );
  NAND2X1 U67969 ( .A(n64096), .B(n64095), .Y(n64097) );
  NAND2X1 U67970 ( .A(n44035), .B(n43518), .Y(n64403) );
  INVX1 U67971 ( .A(n64403), .Y(n64798) );
  NAND2X1 U67972 ( .A(n38378), .B(n43607), .Y(n64400) );
  INVX1 U67973 ( .A(n64400), .Y(n64405) );
  XNOR2X1 U67974 ( .A(n64798), .B(n64405), .Y(n64099) );
  NAND2X1 U67975 ( .A(n43850), .B(n43502), .Y(n64760) );
  INVX1 U67976 ( .A(n64760), .Y(n64755) );
  XNOR2X1 U67977 ( .A(n64099), .B(n64755), .Y(n64100) );
  XNOR2X1 U67978 ( .A(n41802), .B(n64100), .Y(n64107) );
  NOR2X1 U67979 ( .A(n64101), .B(n42166), .Y(n64104) );
  NOR2X1 U67980 ( .A(n64102), .B(n64777), .Y(n64103) );
  NAND2X1 U67981 ( .A(n64104), .B(n64103), .Y(n64105) );
  NAND2X1 U67982 ( .A(n64106), .B(n64105), .Y(n64778) );
  INVX1 U67983 ( .A(n64778), .Y(n64410) );
  XNOR2X1 U67984 ( .A(n64107), .B(n64410), .Y(n64108) );
  XNOR2X1 U67985 ( .A(n64424), .B(n64108), .Y(n64440) );
  NAND2X1 U67986 ( .A(n64427), .B(n64419), .Y(n64119) );
  XNOR2X1 U67987 ( .A(n64129), .B(n64130), .Y(n64118) );
  NOR2X1 U67988 ( .A(n64110), .B(n64109), .Y(n64116) );
  NAND2X1 U67989 ( .A(n64112), .B(n64111), .Y(n64114) );
  NAND2X1 U67990 ( .A(n64114), .B(n64113), .Y(n64115) );
  NOR2X1 U67991 ( .A(n64116), .B(n64115), .Y(n64117) );
  XNOR2X1 U67992 ( .A(n64118), .B(n64117), .Y(n64123) );
  INVX1 U67993 ( .A(n64123), .Y(n64430) );
  NAND2X1 U67994 ( .A(n64119), .B(n64430), .Y(n64761) );
  NAND2X1 U67995 ( .A(n39207), .B(n64120), .Y(n64425) );
  NOR2X1 U67996 ( .A(n38674), .B(n64121), .Y(n64122) );
  NOR2X1 U67997 ( .A(n38504), .B(n64122), .Y(n64124) );
  NAND2X1 U67998 ( .A(n64124), .B(n64123), .Y(n64125) );
  NAND2X1 U67999 ( .A(n64126), .B(n64125), .Y(n64127) );
  NAND2X1 U68000 ( .A(n64761), .B(n64127), .Y(n64439) );
  NAND2X1 U68001 ( .A(n43860), .B(n43497), .Y(n64738) );
  INVX1 U68002 ( .A(n64738), .Y(n64443) );
  XNOR2X1 U68003 ( .A(n64439), .B(n64443), .Y(n64128) );
  XNOR2X1 U68004 ( .A(n64440), .B(n64128), .Y(n64144) );
  INVX1 U68005 ( .A(n64129), .Y(n64132) );
  XNOR2X1 U68006 ( .A(n64431), .B(n64130), .Y(n64131) );
  XNOR2X1 U68007 ( .A(n64132), .B(n64131), .Y(n64134) );
  INVX1 U68008 ( .A(n64139), .Y(n64135) );
  NOR2X1 U68009 ( .A(n36656), .B(n64135), .Y(n64143) );
  NAND2X1 U68010 ( .A(n64137), .B(n64136), .Y(n64138) );
  NOR2X1 U68011 ( .A(n64139), .B(n64138), .Y(n64141) );
  NOR2X1 U68012 ( .A(n64141), .B(n64140), .Y(n64142) );
  OR2X1 U68013 ( .A(n64143), .B(n64142), .Y(n64441) );
  INVX1 U68014 ( .A(n64441), .Y(n64737) );
  XNOR2X1 U68015 ( .A(n64144), .B(n64737), .Y(n64732) );
  XNOR2X1 U68016 ( .A(n64446), .B(n64732), .Y(n64145) );
  XOR2X1 U68017 ( .A(n64445), .B(n64145), .Y(n64393) );
  NOR2X1 U68018 ( .A(n36777), .B(n64148), .Y(n64153) );
  NAND2X1 U68019 ( .A(n64151), .B(n64150), .Y(n64152) );
  NOR2X1 U68020 ( .A(n64153), .B(n64152), .Y(n64154) );
  XNOR2X1 U68021 ( .A(n64155), .B(n64154), .Y(n64383) );
  INVX1 U68022 ( .A(n64383), .Y(n64381) );
  NAND2X1 U68023 ( .A(n43952), .B(n38311), .Y(n64158) );
  NAND2X1 U68024 ( .A(n41176), .B(n64158), .Y(n64157) );
  INVX1 U68025 ( .A(n64380), .Y(n64384) );
  INVX1 U68026 ( .A(n64158), .Y(n64391) );
  NAND2X1 U68027 ( .A(n40990), .B(n64391), .Y(n64156) );
  NAND2X1 U68028 ( .A(n64157), .B(n64156), .Y(n64163) );
  NOR2X1 U68029 ( .A(n41176), .B(n64158), .Y(n64161) );
  NAND2X1 U68030 ( .A(n64159), .B(n64165), .Y(n64160) );
  NAND2X1 U68031 ( .A(n64160), .B(n64167), .Y(n64388) );
  NAND2X1 U68032 ( .A(n64388), .B(n38880), .Y(n64382) );
  NOR2X1 U68033 ( .A(n64163), .B(n64162), .Y(n64164) );
  XOR2X1 U68034 ( .A(n64164), .B(n64393), .Y(n64459) );
  NOR2X1 U68035 ( .A(n64166), .B(n64165), .Y(n64171) );
  NAND2X1 U68036 ( .A(n64168), .B(n64167), .Y(n64169) );
  NAND2X1 U68037 ( .A(n38881), .B(n64169), .Y(n64170) );
  NOR2X1 U68038 ( .A(n64171), .B(n64170), .Y(n64172) );
  XNOR2X1 U68039 ( .A(n64173), .B(n64172), .Y(n64176) );
  NAND2X1 U68040 ( .A(n64176), .B(n64175), .Y(n64178) );
  NAND2X1 U68041 ( .A(n64178), .B(n64177), .Y(n64457) );
  NAND2X1 U68042 ( .A(n64456), .B(n64457), .Y(n64460) );
  INVX1 U68043 ( .A(n64181), .Y(n64373) );
  XNOR2X1 U68044 ( .A(n64182), .B(n39483), .Y(n64183) );
  XNOR2X1 U68045 ( .A(n64373), .B(n41423), .Y(n64700) );
  INVX1 U68046 ( .A(n64375), .Y(n64185) );
  NAND2X1 U68047 ( .A(n43889), .B(n43775), .Y(n64702) );
  NAND2X1 U68048 ( .A(n43896), .B(n43796), .Y(n64471) );
  INVX1 U68049 ( .A(n64471), .Y(n64478) );
  XNOR2X1 U68050 ( .A(n64702), .B(n64478), .Y(n64186) );
  XNOR2X1 U68051 ( .A(n64472), .B(n64186), .Y(n64187) );
  XNOR2X1 U68052 ( .A(n64473), .B(n64187), .Y(n64369) );
  NAND2X1 U68053 ( .A(n43903), .B(n42711), .Y(n64825) );
  INVX1 U68054 ( .A(n64188), .Y(n64199) );
  NOR2X1 U68055 ( .A(n64191), .B(n64190), .Y(n64189) );
  NOR2X1 U68056 ( .A(n64199), .B(n64189), .Y(n64195) );
  NAND2X1 U68057 ( .A(n64191), .B(n64190), .Y(n64193) );
  NAND2X1 U68058 ( .A(n64193), .B(n64192), .Y(n64194) );
  NAND2X1 U68059 ( .A(n64195), .B(n64194), .Y(n64196) );
  NAND2X1 U68060 ( .A(n64197), .B(n64196), .Y(n64367) );
  NAND2X1 U68061 ( .A(n64199), .B(n64198), .Y(n64368) );
  NAND2X1 U68062 ( .A(n64367), .B(n64368), .Y(n64200) );
  XOR2X1 U68063 ( .A(n65122), .B(n64201), .Y(n64358) );
  XNOR2X1 U68064 ( .A(n64361), .B(n64358), .Y(n64219) );
  XNOR2X1 U68065 ( .A(n64202), .B(n41709), .Y(n64203) );
  XNOR2X1 U68066 ( .A(n64203), .B(n36726), .Y(n64216) );
  INVX1 U68067 ( .A(n64209), .Y(n64218) );
  NOR2X1 U68068 ( .A(n64204), .B(n64218), .Y(n64206) );
  NAND2X1 U68069 ( .A(n64206), .B(n64205), .Y(n64212) );
  NAND2X1 U68070 ( .A(n64210), .B(n64209), .Y(n64211) );
  NAND2X1 U68071 ( .A(n64212), .B(n64211), .Y(n64214) );
  NAND2X1 U68072 ( .A(n64214), .B(n64213), .Y(n64215) );
  XNOR2X1 U68073 ( .A(n64219), .B(n38784), .Y(n64354) );
  XOR2X1 U68074 ( .A(n64354), .B(n64351), .Y(n64220) );
  XNOR2X1 U68075 ( .A(n64356), .B(n64220), .Y(n64488) );
  NOR2X1 U68076 ( .A(n41513), .B(n36689), .Y(n64224) );
  NAND2X1 U68077 ( .A(n64224), .B(n64223), .Y(n64229) );
  XNOR2X1 U68078 ( .A(n64226), .B(n64225), .Y(n64227) );
  XNOR2X1 U68079 ( .A(n39758), .B(n64227), .Y(n64228) );
  NAND2X1 U68080 ( .A(n43788), .B(n43973), .Y(n64682) );
  NAND2X1 U68081 ( .A(n43724), .B(n43943), .Y(n64340) );
  INVX1 U68082 ( .A(n64340), .Y(n64495) );
  XNOR2X1 U68083 ( .A(n64682), .B(n64495), .Y(n64230) );
  XNOR2X1 U68084 ( .A(n64231), .B(n64332), .Y(n64232) );
  XNOR2X1 U68085 ( .A(n64233), .B(n64232), .Y(n64936) );
  NAND2X1 U68086 ( .A(n40462), .B(n44001), .Y(n64320) );
  NAND2X1 U68087 ( .A(n40476), .B(n43993), .Y(n64318) );
  INVX1 U68088 ( .A(n64318), .Y(n64326) );
  XNOR2X1 U68089 ( .A(n64320), .B(n64326), .Y(n64234) );
  XNOR2X1 U68090 ( .A(n64313), .B(n42040), .Y(n64242) );
  NAND2X1 U68091 ( .A(n64235), .B(n43984), .Y(n64237) );
  NAND2X1 U68092 ( .A(n64237), .B(n64236), .Y(n64238) );
  NOR2X1 U68093 ( .A(n41564), .B(n41606), .Y(n64241) );
  NAND2X1 U68094 ( .A(n64240), .B(n64239), .Y(n64319) );
  XNOR2X1 U68095 ( .A(n64242), .B(n41298), .Y(n64243) );
  XNOR2X1 U68096 ( .A(n64244), .B(n64243), .Y(n64511) );
  XNOR2X1 U68097 ( .A(n64506), .B(n64511), .Y(n64245) );
  NAND2X1 U68098 ( .A(n43735), .B(n44049), .Y(n64594) );
  NAND2X1 U68099 ( .A(n43759), .B(n44026), .Y(n64601) );
  INVX1 U68100 ( .A(n64601), .Y(n64605) );
  XNOR2X1 U68101 ( .A(n64594), .B(n64605), .Y(n64246) );
  XNOR2X1 U68102 ( .A(n36540), .B(n64246), .Y(n64249) );
  NAND2X1 U68103 ( .A(n64301), .B(n64299), .Y(n64306) );
  INVX1 U68104 ( .A(n64296), .Y(n64248) );
  NAND2X1 U68105 ( .A(n64248), .B(n64297), .Y(n64305) );
  NAND2X1 U68106 ( .A(n64306), .B(n64305), .Y(n64514) );
  INVX1 U68107 ( .A(n64514), .Y(n64604) );
  XNOR2X1 U68108 ( .A(n64249), .B(n64604), .Y(n64250) );
  XNOR2X1 U68109 ( .A(n41331), .B(n64250), .Y(n65185) );
  INVX1 U68110 ( .A(n65185), .Y(n64524) );
  XNOR2X1 U68111 ( .A(n64519), .B(n64524), .Y(n64251) );
  XNOR2X1 U68112 ( .A(n40025), .B(n64251), .Y(n64528) );
  NAND2X1 U68113 ( .A(n43612), .B(n43791), .Y(n72613) );
  XNOR2X1 U68114 ( .A(n64528), .B(n43643), .Y(n64261) );
  XNOR2X1 U68115 ( .A(n43524), .B(n43654), .Y(n72586) );
  NOR2X1 U68116 ( .A(n64252), .B(n64253), .Y(n64256) );
  NOR2X1 U68117 ( .A(n37937), .B(n64254), .Y(n64255) );
  INVX1 U68118 ( .A(n64257), .Y(n64259) );
  INVX1 U68119 ( .A(n64530), .Y(n64290) );
  XNOR2X1 U68120 ( .A(n72586), .B(n64290), .Y(n64260) );
  XNOR2X1 U68121 ( .A(n64261), .B(n64260), .Y(n64268) );
  INVX1 U68122 ( .A(n64263), .Y(n64262) );
  NAND2X1 U68123 ( .A(n64262), .B(n43659), .Y(n64267) );
  NAND2X1 U68124 ( .A(n43663), .B(n64263), .Y(n64264) );
  NAND2X1 U68125 ( .A(n64265), .B(n64264), .Y(n64266) );
  AND2X1 U68126 ( .A(n64266), .B(n64267), .Y(n64538) );
  XNOR2X1 U68127 ( .A(n64268), .B(n64538), .Y(n64269) );
  XNOR2X1 U68128 ( .A(n64582), .B(n43679), .Y(n64270) );
  XNOR2X1 U68129 ( .A(n37905), .B(n64270), .Y(n64287) );
  XNOR2X1 U68130 ( .A(n64287), .B(n43509), .Y(n64275) );
  NAND2X1 U68131 ( .A(n43507), .B(n64271), .Y(n64273) );
  XNOR2X1 U68132 ( .A(n64275), .B(n64289), .Y(n64554) );
  INVX1 U68133 ( .A(n64560), .Y(n64561) );
  XNOR2X1 U68134 ( .A(n43709), .B(n64561), .Y(n64281) );
  NAND2X1 U68135 ( .A(n64277), .B(n43711), .Y(n64279) );
  INVX1 U68136 ( .A(n64562), .Y(n64280) );
  XNOR2X1 U68137 ( .A(n64281), .B(n64280), .Y(n64286) );
  XNOR2X1 U68138 ( .A(n64283), .B(n64282), .Y(n64284) );
  XNOR2X1 U68139 ( .A(n64284), .B(n41908), .Y(n64285) );
  MX2X1 U68140 ( .A(n64286), .B(n64285), .S0(n43720), .Y(u_muldiv_result_r[6])
         );
  NAND2X1 U68141 ( .A(u_muldiv_mult_result_q[6]), .B(n44633), .Y(n14084) );
  NOR2X1 U68142 ( .A(n41229), .B(n41480), .Y(n64289) );
  NAND2X1 U68143 ( .A(n37906), .B(n40203), .Y(n64288) );
  INVX1 U68144 ( .A(n64528), .Y(n64529) );
  NOR2X1 U68145 ( .A(n43642), .B(n64290), .Y(n64291) );
  XNOR2X1 U68146 ( .A(n64529), .B(n64291), .Y(n64536) );
  NAND2X1 U68147 ( .A(n37928), .B(n64536), .Y(n64295) );
  INVX1 U68148 ( .A(n64536), .Y(n64292) );
  NAND2X1 U68149 ( .A(n64292), .B(n43660), .Y(n64293) );
  NAND2X1 U68150 ( .A(n64538), .B(n64293), .Y(n64294) );
  NOR2X1 U68151 ( .A(n64607), .B(n64601), .Y(n64304) );
  NOR2X1 U68152 ( .A(n64601), .B(n64296), .Y(n64298) );
  INVX1 U68153 ( .A(n64299), .Y(n64300) );
  NOR2X1 U68154 ( .A(n64300), .B(n64601), .Y(n64302) );
  NOR2X1 U68155 ( .A(n64304), .B(n64303), .Y(n64309) );
  NAND2X1 U68156 ( .A(n64305), .B(n64306), .Y(n64307) );
  NAND2X1 U68157 ( .A(n36540), .B(n64307), .Y(n64308) );
  NAND2X1 U68158 ( .A(n64309), .B(n64308), .Y(n64627) );
  INVX1 U68159 ( .A(n64648), .Y(n64315) );
  XNOR2X1 U68160 ( .A(n41298), .B(n64313), .Y(n64650) );
  INVX1 U68161 ( .A(n64650), .Y(n64641) );
  NOR2X1 U68162 ( .A(n38989), .B(n64315), .Y(n64316) );
  NAND2X1 U68163 ( .A(n64316), .B(n40200), .Y(n64640) );
  INVX1 U68164 ( .A(n64936), .Y(n64669) );
  INVX1 U68165 ( .A(n64320), .Y(n64663) );
  INVX1 U68166 ( .A(n64667), .Y(n64658) );
  XNOR2X1 U68167 ( .A(n64658), .B(n42047), .Y(n64504) );
  NOR2X1 U68168 ( .A(n36531), .B(n64669), .Y(n64324) );
  NAND2X1 U68169 ( .A(n64324), .B(n64329), .Y(n64325) );
  NAND2X1 U68170 ( .A(n64326), .B(n64325), .Y(n64331) );
  NAND2X1 U68171 ( .A(n64330), .B(n64329), .Y(n64934) );
  NAND2X1 U68172 ( .A(n64934), .B(n64669), .Y(n64670) );
  NAND2X1 U68173 ( .A(n64331), .B(n64670), .Y(n64677) );
  XNOR2X1 U68174 ( .A(n40078), .B(n64332), .Y(n64857) );
  NAND2X1 U68175 ( .A(n64857), .B(n64334), .Y(n64861) );
  NOR2X1 U68176 ( .A(n64858), .B(n64857), .Y(n64335) );
  NAND2X1 U68177 ( .A(n64335), .B(n64859), .Y(n64336) );
  NAND2X1 U68178 ( .A(n42004), .B(n64336), .Y(n64337) );
  NAND2X1 U68179 ( .A(n64861), .B(n64337), .Y(n65157) );
  INVX1 U68180 ( .A(n65157), .Y(n64676) );
  NAND2X1 U68181 ( .A(n40470), .B(n44001), .Y(n64673) );
  INVX1 U68182 ( .A(n64673), .Y(n64938) );
  XNOR2X1 U68183 ( .A(n64676), .B(n64938), .Y(n64502) );
  INVX1 U68184 ( .A(n64682), .Y(n64338) );
  INVX1 U68185 ( .A(n64497), .Y(n64339) );
  XNOR2X1 U68186 ( .A(n64340), .B(n64339), .Y(n64341) );
  NOR2X1 U68187 ( .A(n41552), .B(n64684), .Y(n64343) );
  INVX1 U68188 ( .A(n64683), .Y(n64685) );
  NAND2X1 U68189 ( .A(n64685), .B(n64686), .Y(n64342) );
  NAND2X1 U68190 ( .A(n64343), .B(n64342), .Y(n64863) );
  INVX1 U68191 ( .A(n64344), .Y(n64347) );
  NAND2X1 U68192 ( .A(n64347), .B(n64345), .Y(n64692) );
  INVX1 U68193 ( .A(n64692), .Y(n64349) );
  NAND2X1 U68194 ( .A(n64347), .B(n64346), .Y(n64691) );
  INVX1 U68195 ( .A(n64691), .Y(n64348) );
  NOR2X1 U68196 ( .A(n64349), .B(n64348), .Y(n64350) );
  NAND2X1 U68197 ( .A(n64690), .B(n64350), .Y(n64494) );
  NAND2X1 U68198 ( .A(n40260), .B(n43934), .Y(n64851) );
  NAND2X1 U68199 ( .A(n43928), .B(n43798), .Y(n64842) );
  NOR2X1 U68200 ( .A(n64354), .B(n64351), .Y(n64353) );
  INVX1 U68201 ( .A(n64354), .Y(n64355) );
  NAND2X1 U68202 ( .A(n64356), .B(n64355), .Y(n64357) );
  NOR2X1 U68203 ( .A(n64358), .B(n64361), .Y(n64360) );
  NOR2X1 U68204 ( .A(n39338), .B(n64358), .Y(n64359) );
  NOR2X1 U68205 ( .A(n64360), .B(n64359), .Y(n64365) );
  INVX1 U68206 ( .A(n64361), .Y(n64363) );
  NAND2X1 U68207 ( .A(n64363), .B(n64362), .Y(n64364) );
  NAND2X1 U68208 ( .A(n64365), .B(n64364), .Y(n64838) );
  INVX1 U68209 ( .A(n64825), .Y(n65124) );
  XNOR2X1 U68210 ( .A(n64369), .B(n41156), .Y(n64826) );
  INVX1 U68211 ( .A(n64826), .Y(n65123) );
  NOR2X1 U68212 ( .A(n41132), .B(n39101), .Y(n64371) );
  NAND2X1 U68213 ( .A(n65123), .B(n64370), .Y(n65130) );
  NAND2X1 U68214 ( .A(n64371), .B(n65130), .Y(n65311) );
  INVX1 U68215 ( .A(n64702), .Y(n64703) );
  NAND2X1 U68216 ( .A(n64703), .B(n64472), .Y(n64379) );
  NOR2X1 U68217 ( .A(n36658), .B(n41188), .Y(n64374) );
  NOR2X1 U68218 ( .A(n36768), .B(n64374), .Y(n64378) );
  NOR2X1 U68219 ( .A(n41188), .B(n64375), .Y(n64376) );
  NOR2X1 U68220 ( .A(n64703), .B(n64376), .Y(n64377) );
  NAND2X1 U68221 ( .A(n64379), .B(n64707), .Y(n64816) );
  NAND2X1 U68222 ( .A(n43903), .B(n43796), .Y(n64820) );
  INVX1 U68223 ( .A(n64820), .Y(n64818) );
  XNOR2X1 U68224 ( .A(n64816), .B(n64818), .Y(n64470) );
  NAND2X1 U68225 ( .A(n64387), .B(n64382), .Y(n64385) );
  NAND2X1 U68226 ( .A(n64384), .B(n64383), .Y(n64390) );
  NAND2X1 U68227 ( .A(n64385), .B(n64390), .Y(n64386) );
  NAND2X1 U68228 ( .A(n64391), .B(n64386), .Y(n65016) );
  NOR2X1 U68229 ( .A(n39836), .B(n38881), .Y(n64389) );
  NOR2X1 U68230 ( .A(n64391), .B(n40990), .Y(n64392) );
  NAND2X1 U68231 ( .A(n65016), .B(n65017), .Y(n65010) );
  NAND2X1 U68232 ( .A(n44035), .B(n43607), .Y(n64772) );
  NAND2X1 U68233 ( .A(n64405), .B(n43605), .Y(n64774) );
  INVX1 U68234 ( .A(n64774), .Y(n65077) );
  NOR2X1 U68235 ( .A(n42237), .B(n64394), .Y(n64396) );
  NOR2X1 U68236 ( .A(n38610), .B(n64406), .Y(n64395) );
  NAND2X1 U68237 ( .A(n64396), .B(n64395), .Y(n65078) );
  NOR2X1 U68238 ( .A(n64410), .B(n41802), .Y(n64397) );
  NOR2X1 U68239 ( .A(n64397), .B(n64400), .Y(n64398) );
  XNOR2X1 U68240 ( .A(n64399), .B(n64398), .Y(n65058) );
  NAND2X1 U68241 ( .A(n43850), .B(n39960), .Y(n64793) );
  INVX1 U68242 ( .A(n64793), .Y(n65059) );
  XNOR2X1 U68243 ( .A(n65058), .B(n65059), .Y(n64417) );
  XNOR2X1 U68244 ( .A(n64400), .B(n41802), .Y(n64401) );
  XNOR2X1 U68245 ( .A(n64410), .B(n64401), .Y(n64794) );
  INVX1 U68246 ( .A(n64794), .Y(n64416) );
  NAND2X1 U68247 ( .A(n64402), .B(n64416), .Y(n65048) );
  NOR2X1 U68248 ( .A(n36779), .B(n65048), .Y(n64412) );
  NOR2X1 U68249 ( .A(n64413), .B(n64403), .Y(n64404) );
  NAND2X1 U68250 ( .A(n64404), .B(n64415), .Y(n65065) );
  XNOR2X1 U68251 ( .A(n64406), .B(n64405), .Y(n64408) );
  NOR2X1 U68252 ( .A(n64777), .B(n41803), .Y(n64407) );
  XNOR2X1 U68253 ( .A(n64408), .B(n64407), .Y(n64409) );
  XNOR2X1 U68254 ( .A(n64410), .B(n64409), .Y(n64411) );
  NAND2X1 U68255 ( .A(n64798), .B(n64411), .Y(n65064) );
  NAND2X1 U68256 ( .A(n65065), .B(n65064), .Y(n64797) );
  NOR2X1 U68257 ( .A(n64412), .B(n64797), .Y(n64786) );
  NAND2X1 U68258 ( .A(n41805), .B(n64413), .Y(n64414) );
  NAND2X1 U68259 ( .A(n64786), .B(n39613), .Y(n64804) );
  INVX1 U68260 ( .A(n64804), .Y(n64771) );
  XNOR2X1 U68261 ( .A(n64417), .B(n64771), .Y(n64768) );
  NAND2X1 U68262 ( .A(n43962), .B(n43496), .Y(n65089) );
  NAND2X1 U68263 ( .A(n43859), .B(n43501), .Y(n64766) );
  INVX1 U68264 ( .A(n64766), .Y(n64770) );
  XNOR2X1 U68265 ( .A(n65089), .B(n64770), .Y(n64418) );
  XNOR2X1 U68266 ( .A(n64768), .B(n64418), .Y(n64438) );
  NOR2X1 U68267 ( .A(n64431), .B(n64760), .Y(n64422) );
  NOR2X1 U68268 ( .A(n38504), .B(n64430), .Y(n64420) );
  NAND2X1 U68269 ( .A(n64420), .B(n64419), .Y(n64421) );
  NAND2X1 U68270 ( .A(n64422), .B(n64421), .Y(n65043) );
  XNOR2X1 U68271 ( .A(n64794), .B(n64798), .Y(n64423) );
  XNOR2X1 U68272 ( .A(n64424), .B(n64423), .Y(n64433) );
  NAND2X1 U68273 ( .A(n64755), .B(n64433), .Y(n65040) );
  NAND2X1 U68274 ( .A(n65043), .B(n65040), .Y(n64436) );
  INVX1 U68275 ( .A(n64761), .Y(n64756) );
  INVX1 U68276 ( .A(n64433), .Y(n64758) );
  NAND2X1 U68277 ( .A(n64426), .B(n64425), .Y(n64428) );
  NAND2X1 U68278 ( .A(n64428), .B(n64427), .Y(n64429) );
  NOR2X1 U68279 ( .A(n64430), .B(n64429), .Y(n64432) );
  NOR2X1 U68280 ( .A(n64432), .B(n64431), .Y(n64434) );
  NAND2X1 U68281 ( .A(n64434), .B(n64433), .Y(n64754) );
  NAND2X1 U68282 ( .A(n64744), .B(n64754), .Y(n64435) );
  NOR2X1 U68283 ( .A(n64436), .B(n64435), .Y(n64437) );
  XNOR2X1 U68284 ( .A(n64438), .B(n64437), .Y(n64727) );
  XNOR2X1 U68285 ( .A(n64727), .B(n41508), .Y(n64444) );
  NAND2X1 U68286 ( .A(n64740), .B(n64441), .Y(n64751) );
  INVX1 U68287 ( .A(n64739), .Y(n64442) );
  NAND2X1 U68288 ( .A(n64443), .B(n64442), .Y(n64750) );
  XNOR2X1 U68289 ( .A(n64444), .B(n40996), .Y(n64721) );
  INVX1 U68290 ( .A(n64446), .Y(n64723) );
  NOR2X1 U68291 ( .A(n64448), .B(n40151), .Y(n64449) );
  NOR2X1 U68292 ( .A(n64732), .B(n64449), .Y(n64450) );
  NAND2X1 U68293 ( .A(n64450), .B(n64730), .Y(n64722) );
  NAND2X1 U68294 ( .A(n64723), .B(n64722), .Y(n64451) );
  NAND2X1 U68295 ( .A(n65025), .B(n64451), .Y(n64452) );
  XNOR2X1 U68296 ( .A(n64452), .B(n37408), .Y(n64453) );
  XNOR2X1 U68297 ( .A(n64721), .B(n64453), .Y(n64454) );
  NAND2X1 U68298 ( .A(n43879), .B(n38313), .Y(n64997) );
  INVX1 U68299 ( .A(n64455), .Y(n64461) );
  NOR2X1 U68300 ( .A(n64461), .B(n39854), .Y(n64458) );
  INVX1 U68301 ( .A(n64462), .Y(n64465) );
  NAND2X1 U68302 ( .A(n64465), .B(n64463), .Y(n65101) );
  NOR2X1 U68303 ( .A(n64465), .B(n38864), .Y(n64467) );
  NAND2X1 U68304 ( .A(n65101), .B(n65100), .Y(n65105) );
  NAND2X1 U68305 ( .A(n43889), .B(n43478), .Y(n64717) );
  NAND2X1 U68306 ( .A(n43896), .B(n43775), .Y(n64712) );
  XNOR2X1 U68307 ( .A(n64717), .B(n64712), .Y(n64468) );
  XOR2X1 U68308 ( .A(n65105), .B(n64468), .Y(n64469) );
  XNOR2X1 U68309 ( .A(n65106), .B(n64469), .Y(n64817) );
  XNOR2X1 U68310 ( .A(n64470), .B(n64817), .Y(n64824) );
  NOR2X1 U68311 ( .A(n41156), .B(n64471), .Y(n64476) );
  INVX1 U68312 ( .A(n64477), .Y(n64474) );
  NOR2X1 U68313 ( .A(n41156), .B(n64474), .Y(n64475) );
  NOR2X1 U68314 ( .A(n64476), .B(n64475), .Y(n64480) );
  NAND2X1 U68315 ( .A(n64478), .B(n64477), .Y(n64479) );
  NAND2X1 U68316 ( .A(n64480), .B(n64479), .Y(n64823) );
  NAND2X1 U68317 ( .A(n43909), .B(n42711), .Y(n65337) );
  INVX1 U68318 ( .A(n65337), .Y(n65312) );
  XNOR2X1 U68319 ( .A(n64823), .B(n65312), .Y(n64481) );
  XNOR2X1 U68320 ( .A(n64824), .B(n64481), .Y(n64482) );
  XNOR2X1 U68321 ( .A(n36709), .B(n64482), .Y(n64839) );
  NAND2X1 U68322 ( .A(n42654), .B(n43920), .Y(n64835) );
  XOR2X1 U68323 ( .A(n64839), .B(n64835), .Y(n64483) );
  XNOR2X1 U68324 ( .A(n64838), .B(n64483), .Y(n64843) );
  XNOR2X1 U68325 ( .A(n64484), .B(n64843), .Y(n64852) );
  INVX1 U68326 ( .A(n64852), .Y(n64847) );
  INVX1 U68327 ( .A(n64487), .Y(n64485) );
  NOR2X1 U68328 ( .A(n64485), .B(n64486), .Y(n64492) );
  NOR2X1 U68329 ( .A(n64488), .B(n64486), .Y(n64490) );
  OR2X1 U68330 ( .A(n64490), .B(n64489), .Y(n64491) );
  NOR2X1 U68331 ( .A(n64492), .B(n64491), .Y(n64848) );
  XNOR2X1 U68332 ( .A(n64848), .B(n64493), .Y(n64970) );
  NAND2X1 U68333 ( .A(n42643), .B(n43943), .Y(n64695) );
  XNOR2X1 U68334 ( .A(n64494), .B(n39014), .Y(n64954) );
  INVX1 U68335 ( .A(n64954), .Y(n64950) );
  NAND2X1 U68336 ( .A(n64495), .B(n64496), .Y(n64688) );
  NAND2X1 U68337 ( .A(n64497), .B(n64496), .Y(n64689) );
  NAND2X1 U68338 ( .A(n64688), .B(n64689), .Y(n64498) );
  NOR2X1 U68339 ( .A(n38697), .B(n64498), .Y(n64499) );
  XNOR2X1 U68340 ( .A(n64500), .B(n64499), .Y(n64864) );
  NAND2X1 U68341 ( .A(n40489), .B(n43993), .Y(n64856) );
  XNOR2X1 U68342 ( .A(n64856), .B(n41999), .Y(n64501) );
  INVX1 U68343 ( .A(n64668), .Y(n64657) );
  INVX1 U68344 ( .A(n64659), .Y(n64503) );
  NAND2X1 U68345 ( .A(n43758), .B(n44049), .Y(n64600) );
  NAND2X1 U68346 ( .A(n43820), .B(n44026), .Y(n64608) );
  INVX1 U68347 ( .A(n64608), .Y(n64633) );
  XNOR2X1 U68348 ( .A(n64600), .B(n64633), .Y(n64505) );
  XNOR2X1 U68349 ( .A(n36566), .B(n64505), .Y(n64512) );
  INVX1 U68350 ( .A(n64506), .Y(n64509) );
  NAND2X1 U68351 ( .A(n64509), .B(n64631), .Y(n64635) );
  NAND2X1 U68352 ( .A(n64511), .B(n64510), .Y(n64634) );
  NAND2X1 U68353 ( .A(n43735), .B(n44056), .Y(n64591) );
  INVX1 U68354 ( .A(n64591), .Y(n64597) );
  XNOR2X1 U68355 ( .A(n64595), .B(n64597), .Y(n64518) );
  XNOR2X1 U68356 ( .A(n64607), .B(n64601), .Y(n64513) );
  XOR2X1 U68357 ( .A(n64514), .B(n64513), .Y(n64589) );
  NOR2X1 U68358 ( .A(n38363), .B(n64594), .Y(n64516) );
  NOR2X1 U68359 ( .A(n41331), .B(n64589), .Y(n64515) );
  NOR2X1 U68360 ( .A(n64515), .B(n64516), .Y(n64517) );
  XNOR2X1 U68361 ( .A(n64518), .B(n64517), .Y(n64873) );
  NAND2X1 U68362 ( .A(n43612), .B(n43780), .Y(n72626) );
  XNOR2X1 U68363 ( .A(n64873), .B(n43666), .Y(n64526) );
  INVX1 U68364 ( .A(n64519), .Y(n65187) );
  NOR2X1 U68365 ( .A(n38576), .B(n64524), .Y(n64522) );
  NAND2X1 U68366 ( .A(n64522), .B(n64521), .Y(n64523) );
  XNOR2X1 U68367 ( .A(n64881), .B(n43643), .Y(n64527) );
  XNOR2X1 U68368 ( .A(n43655), .B(n64527), .Y(n64534) );
  NAND2X1 U68369 ( .A(n43644), .B(n64528), .Y(n64533) );
  NAND2X1 U68370 ( .A(n64529), .B(n43649), .Y(n64531) );
  NAND2X1 U68371 ( .A(n64531), .B(n64530), .Y(n64532) );
  XNOR2X1 U68372 ( .A(n64534), .B(n41365), .Y(n64535) );
  XNOR2X1 U68373 ( .A(n41154), .B(n64535), .Y(n64886) );
  INVX1 U68374 ( .A(n64886), .Y(n64885) );
  XNOR2X1 U68375 ( .A(n64536), .B(n43654), .Y(n64537) );
  XNOR2X1 U68376 ( .A(n64538), .B(n64537), .Y(n64540) );
  INVX1 U68377 ( .A(n64540), .Y(n64539) );
  NAND2X1 U68378 ( .A(n64539), .B(n43532), .Y(n64544) );
  NAND2X1 U68379 ( .A(n43521), .B(n64540), .Y(n64542) );
  NAND2X1 U68380 ( .A(n64542), .B(n64541), .Y(n64543) );
  NAND2X1 U68381 ( .A(n64544), .B(n64543), .Y(n64884) );
  XNOR2X1 U68382 ( .A(n64884), .B(n43524), .Y(n64545) );
  XNOR2X1 U68383 ( .A(n64885), .B(n64545), .Y(n64580) );
  INVX1 U68384 ( .A(n64580), .Y(n64581) );
  NOR2X1 U68385 ( .A(n64581), .B(n64547), .Y(n64550) );
  NOR2X1 U68386 ( .A(n43678), .B(n64582), .Y(n64546) );
  NAND2X1 U68387 ( .A(n64546), .B(n64583), .Y(n64551) );
  NAND2X1 U68388 ( .A(n64551), .B(n64547), .Y(n64548) );
  NOR2X1 U68389 ( .A(n64580), .B(n64548), .Y(n64549) );
  INVX1 U68390 ( .A(n64551), .Y(n64552) );
  INVX1 U68391 ( .A(n64891), .Y(n64890) );
  INVX1 U68392 ( .A(n64554), .Y(n64553) );
  NAND2X1 U68393 ( .A(n64553), .B(n43700), .Y(n64558) );
  NAND2X1 U68394 ( .A(n41454), .B(n64554), .Y(n64556) );
  NAND2X1 U68395 ( .A(n64556), .B(n64555), .Y(n64557) );
  NAND2X1 U68396 ( .A(n64558), .B(n64557), .Y(n64892) );
  XNOR2X1 U68397 ( .A(n64892), .B(n43693), .Y(n64559) );
  XNOR2X1 U68398 ( .A(n64890), .B(n64559), .Y(n64573) );
  INVX1 U68399 ( .A(n64573), .Y(n64574) );
  XNOR2X1 U68400 ( .A(n43709), .B(n64574), .Y(n64567) );
  NAND2X1 U68401 ( .A(n43706), .B(n64560), .Y(n64565) );
  NAND2X1 U68402 ( .A(n64561), .B(n43715), .Y(n64563) );
  NAND2X1 U68403 ( .A(n64563), .B(n64562), .Y(n64564) );
  NAND2X1 U68404 ( .A(n64565), .B(n64564), .Y(n64575) );
  INVX1 U68405 ( .A(n64575), .Y(n64566) );
  XNOR2X1 U68406 ( .A(n64567), .B(n64566), .Y(n64572) );
  XNOR2X1 U68407 ( .A(n64569), .B(n64568), .Y(n64570) );
  XNOR2X1 U68408 ( .A(n41918), .B(n64570), .Y(n64571) );
  MX2X1 U68409 ( .A(n64572), .B(n64571), .S0(n43720), .Y(u_muldiv_result_r[7])
         );
  NAND2X1 U68410 ( .A(u_muldiv_mult_result_q[7]), .B(n44633), .Y(n14073) );
  INVX1 U68411 ( .A(n37920), .Y(n64896) );
  NAND2X1 U68412 ( .A(n64577), .B(n40203), .Y(n64579) );
  NAND2X1 U68413 ( .A(n64578), .B(n64579), .Y(n65589) );
  NAND2X1 U68414 ( .A(n43676), .B(n64580), .Y(n65556) );
  NAND2X1 U68415 ( .A(n64581), .B(n43684), .Y(n64586) );
  NAND2X1 U68416 ( .A(n64582), .B(n43686), .Y(n64584) );
  NAND2X1 U68417 ( .A(n64586), .B(n64585), .Y(n65555) );
  NAND2X1 U68418 ( .A(n65556), .B(n65555), .Y(n64904) );
  NAND2X1 U68419 ( .A(n64597), .B(n64595), .Y(n64592) );
  NAND2X1 U68420 ( .A(n64593), .B(n64592), .Y(n65904) );
  INVX1 U68421 ( .A(n64594), .Y(n64596) );
  NAND2X1 U68422 ( .A(n64597), .B(n44049), .Y(n64598) );
  INVX1 U68423 ( .A(n65179), .Y(n65183) );
  XNOR2X1 U68424 ( .A(n43666), .B(n65183), .Y(n64872) );
  INVX1 U68425 ( .A(n64600), .Y(n64609) );
  NAND2X1 U68426 ( .A(n64607), .B(n64601), .Y(n64602) );
  NAND2X1 U68427 ( .A(n64609), .B(n64602), .Y(n64603) );
  NOR2X1 U68428 ( .A(n64604), .B(n64603), .Y(n64625) );
  NAND2X1 U68429 ( .A(n64605), .B(n64609), .Y(n64606) );
  NOR2X1 U68430 ( .A(n64607), .B(n64606), .Y(n64615) );
  NAND2X1 U68431 ( .A(n64609), .B(n64608), .Y(n64616) );
  NAND2X1 U68432 ( .A(n64636), .B(n64616), .Y(n64611) );
  NAND2X1 U68433 ( .A(n64609), .B(n64633), .Y(n64619) );
  NAND2X1 U68434 ( .A(n64619), .B(n36566), .Y(n64610) );
  NAND2X1 U68435 ( .A(n64611), .B(n64610), .Y(n64612) );
  NOR2X1 U68436 ( .A(n64613), .B(n64612), .Y(n64614) );
  NOR2X1 U68437 ( .A(n64615), .B(n64614), .Y(n64623) );
  INVX1 U68438 ( .A(n64616), .Y(n64617) );
  NOR2X1 U68439 ( .A(n64636), .B(n64617), .Y(n64618) );
  NOR2X1 U68440 ( .A(n38129), .B(n64618), .Y(n64621) );
  NAND2X1 U68441 ( .A(n64636), .B(n64619), .Y(n64620) );
  NAND2X1 U68442 ( .A(n64621), .B(n64620), .Y(n64622) );
  NAND2X1 U68443 ( .A(n64623), .B(n64622), .Y(n64624) );
  NOR2X1 U68444 ( .A(n64625), .B(n64624), .Y(n64630) );
  XNOR2X1 U68445 ( .A(n64633), .B(n36566), .Y(n64626) );
  XNOR2X1 U68446 ( .A(n64626), .B(n38129), .Y(n64628) );
  NAND2X1 U68447 ( .A(n64628), .B(n64627), .Y(n64629) );
  NAND2X1 U68448 ( .A(n64630), .B(n64629), .Y(n65177) );
  NAND2X1 U68449 ( .A(n43612), .B(n43738), .Y(n72591) );
  NAND2X1 U68450 ( .A(n64633), .B(n64632), .Y(n64925) );
  NAND2X1 U68451 ( .A(n64633), .B(n64636), .Y(n64924) );
  INVX1 U68452 ( .A(n64924), .Y(n64928) );
  NOR2X1 U68453 ( .A(n39848), .B(n64928), .Y(n64637) );
  NAND2X1 U68454 ( .A(n64637), .B(n64929), .Y(n65252) );
  NAND2X1 U68455 ( .A(n43820), .B(n44049), .Y(n64917) );
  INVX1 U68456 ( .A(n64917), .Y(n65261) );
  NAND2X1 U68457 ( .A(n43758), .B(n44056), .Y(n64919) );
  INVX1 U68458 ( .A(n64919), .Y(n64923) );
  XNOR2X1 U68459 ( .A(n65261), .B(n64923), .Y(n64870) );
  XNOR2X1 U68460 ( .A(n64659), .B(n64658), .Y(n64639) );
  NAND2X1 U68461 ( .A(n64639), .B(n64638), .Y(n65273) );
  NAND2X1 U68462 ( .A(n64642), .B(n43993), .Y(n64643) );
  NOR2X1 U68463 ( .A(n41360), .B(n64643), .Y(n64647) );
  NOR2X1 U68464 ( .A(n64645), .B(n64644), .Y(n64646) );
  NOR2X1 U68465 ( .A(n64647), .B(n64646), .Y(n64649) );
  NAND2X1 U68466 ( .A(n64649), .B(n64648), .Y(n64652) );
  NOR2X1 U68467 ( .A(n64652), .B(n64651), .Y(n64654) );
  NAND2X1 U68468 ( .A(n42047), .B(n42040), .Y(n64653) );
  NOR2X1 U68469 ( .A(n64654), .B(n64653), .Y(n64655) );
  NOR2X1 U68470 ( .A(n64656), .B(n64655), .Y(n64661) );
  XNOR2X1 U68471 ( .A(n64657), .B(n42044), .Y(n64659) );
  NAND2X1 U68472 ( .A(n42047), .B(n64639), .Y(n64660) );
  NAND2X1 U68473 ( .A(n64661), .B(n64660), .Y(n65271) );
  NOR2X1 U68474 ( .A(n37366), .B(n64668), .Y(n64665) );
  NAND2X1 U68475 ( .A(n41298), .B(n38680), .Y(n64662) );
  NAND2X1 U68476 ( .A(n64663), .B(n64662), .Y(n64664) );
  NAND2X1 U68477 ( .A(n64665), .B(n64664), .Y(n64666) );
  NAND2X1 U68478 ( .A(n42044), .B(n64666), .Y(n65523) );
  NAND2X1 U68479 ( .A(n43809), .B(n44026), .Y(n65270) );
  NOR2X1 U68480 ( .A(n43995), .B(n38669), .Y(n64672) );
  NAND2X1 U68481 ( .A(n64669), .B(n43992), .Y(n64933) );
  NAND2X1 U68482 ( .A(n64933), .B(n64670), .Y(n64671) );
  NOR2X1 U68483 ( .A(n64672), .B(n64671), .Y(n64674) );
  NAND2X1 U68484 ( .A(n41428), .B(n64677), .Y(n64942) );
  NOR2X1 U68485 ( .A(n43979), .B(n39988), .Y(n64679) );
  NOR2X1 U68486 ( .A(n43979), .B(n64683), .Y(n64678) );
  NOR2X1 U68487 ( .A(n64679), .B(n64678), .Y(n64681) );
  NAND2X1 U68488 ( .A(n64686), .B(n64685), .Y(n64680) );
  NOR2X1 U68489 ( .A(n64683), .B(n64682), .Y(n64684) );
  NAND2X1 U68490 ( .A(n40482), .B(n44001), .Y(n65163) );
  NAND2X1 U68491 ( .A(n40361), .B(n64953), .Y(n64960) );
  NOR2X1 U68492 ( .A(n64970), .B(n64695), .Y(n64694) );
  INVX1 U68493 ( .A(n64972), .Y(n64967) );
  NOR2X1 U68494 ( .A(n64970), .B(n64967), .Y(n64693) );
  NOR2X1 U68495 ( .A(n64694), .B(n64693), .Y(n64698) );
  INVX1 U68496 ( .A(n64695), .Y(n64696) );
  NAND2X1 U68497 ( .A(n64696), .B(n64972), .Y(n64697) );
  NAND2X1 U68498 ( .A(n64698), .B(n64697), .Y(n64978) );
  NAND2X1 U68499 ( .A(n42644), .B(n43973), .Y(n64966) );
  NAND2X1 U68500 ( .A(n43918), .B(n42711), .Y(n65336) );
  NAND2X1 U68501 ( .A(n43909), .B(n43795), .Y(n64983) );
  NAND2X1 U68502 ( .A(n64700), .B(n64699), .Y(n64701) );
  NOR2X1 U68503 ( .A(n64702), .B(n64701), .Y(n64706) );
  NAND2X1 U68504 ( .A(n36768), .B(n64703), .Y(n64704) );
  NAND2X1 U68505 ( .A(n64704), .B(n64712), .Y(n64705) );
  NOR2X1 U68506 ( .A(n64706), .B(n64705), .Y(n64708) );
  NAND2X1 U68507 ( .A(n64708), .B(n64707), .Y(n64711) );
  INVX1 U68508 ( .A(n64717), .Y(n65104) );
  XNOR2X1 U68509 ( .A(n65104), .B(n38867), .Y(n64709) );
  NAND2X1 U68510 ( .A(n64711), .B(n64710), .Y(n64715) );
  INVX1 U68511 ( .A(n64712), .Y(n64713) );
  NAND2X1 U68512 ( .A(n64713), .B(n36659), .Y(n64714) );
  NAND2X1 U68513 ( .A(n64715), .B(n64714), .Y(n64993) );
  NAND2X1 U68514 ( .A(n43903), .B(n43775), .Y(n65352) );
  NAND2X1 U68515 ( .A(n65100), .B(n65101), .Y(n64720) );
  NOR2X1 U68516 ( .A(n39826), .B(n64717), .Y(n64719) );
  NOR2X1 U68517 ( .A(n38867), .B(n64717), .Y(n64718) );
  NAND2X1 U68518 ( .A(n43896), .B(n43478), .Y(n65099) );
  NAND2X1 U68519 ( .A(n37408), .B(n65019), .Y(n65012) );
  INVX1 U68520 ( .A(n65012), .Y(n64726) );
  NAND2X1 U68521 ( .A(n65019), .B(n65010), .Y(n65015) );
  NAND2X1 U68522 ( .A(n37408), .B(n40272), .Y(n64724) );
  NAND2X1 U68523 ( .A(n65015), .B(n64724), .Y(n64725) );
  NOR2X1 U68524 ( .A(n64726), .B(n64725), .Y(n64810) );
  NAND2X1 U68525 ( .A(n64451), .B(n65025), .Y(n64728) );
  NAND2X1 U68526 ( .A(n64728), .B(n39819), .Y(n64736) );
  NAND2X1 U68527 ( .A(n64730), .B(n64729), .Y(n64731) );
  NAND2X1 U68528 ( .A(n64732), .B(n64731), .Y(n64733) );
  NAND2X1 U68529 ( .A(n41508), .B(n64734), .Y(n64735) );
  NAND2X1 U68530 ( .A(n64736), .B(n64735), .Y(n65035) );
  NAND2X1 U68531 ( .A(n43879), .B(n43486), .Y(n65014) );
  NAND2X1 U68532 ( .A(n64737), .B(n64750), .Y(n64741) );
  NAND2X1 U68533 ( .A(n64739), .B(n64738), .Y(n64740) );
  NAND2X1 U68534 ( .A(n64741), .B(n64740), .Y(n64742) );
  NOR2X1 U68535 ( .A(n65089), .B(n64742), .Y(n64749) );
  XNOR2X1 U68536 ( .A(n64768), .B(n64770), .Y(n64747) );
  NAND2X1 U68537 ( .A(n64756), .B(n64743), .Y(n64744) );
  NAND2X1 U68538 ( .A(n64744), .B(n64754), .Y(n64745) );
  NOR2X1 U68539 ( .A(n64436), .B(n64745), .Y(n64746) );
  XNOR2X1 U68540 ( .A(n64747), .B(n64746), .Y(n64753) );
  INVX1 U68541 ( .A(n64753), .Y(n65090) );
  NOR2X1 U68542 ( .A(n65090), .B(n65089), .Y(n64748) );
  NAND2X1 U68543 ( .A(n64751), .B(n64750), .Y(n64752) );
  INVX1 U68544 ( .A(n64754), .Y(n65042) );
  NOR2X1 U68545 ( .A(n64756), .B(n64755), .Y(n64757) );
  NOR2X1 U68546 ( .A(n64758), .B(n64757), .Y(n64759) );
  NOR2X1 U68547 ( .A(n65042), .B(n64759), .Y(n64765) );
  INVX1 U68548 ( .A(n65043), .Y(n64763) );
  NOR2X1 U68549 ( .A(n64761), .B(n64760), .Y(n64762) );
  NOR2X1 U68550 ( .A(n64763), .B(n64762), .Y(n64764) );
  NAND2X1 U68551 ( .A(n64765), .B(n64764), .Y(n64767) );
  NAND2X1 U68552 ( .A(n64768), .B(n64766), .Y(n65413) );
  INVX1 U68553 ( .A(n64768), .Y(n64769) );
  NAND2X1 U68554 ( .A(n64770), .B(n64769), .Y(n65039) );
  XNOR2X1 U68555 ( .A(n65086), .B(n41507), .Y(n64807) );
  NAND2X1 U68556 ( .A(n43962), .B(n43501), .Y(n65416) );
  INVX1 U68557 ( .A(n65058), .Y(n65049) );
  NOR2X1 U68558 ( .A(n64771), .B(n65049), .Y(n64784) );
  NAND2X1 U68559 ( .A(n43859), .B(n43517), .Y(n65055) );
  INVX1 U68560 ( .A(n64772), .Y(n64781) );
  NAND2X1 U68561 ( .A(n64781), .B(n43605), .Y(n66126) );
  INVX1 U68562 ( .A(n66126), .Y(n66132) );
  NAND2X1 U68563 ( .A(n64774), .B(n64773), .Y(n64775) );
  OR2X1 U68564 ( .A(n41803), .B(n64775), .Y(n64776) );
  NOR2X1 U68565 ( .A(n64777), .B(n64776), .Y(n65075) );
  XNOR2X1 U68566 ( .A(n66132), .B(n65075), .Y(n66131) );
  INVX1 U68567 ( .A(n66131), .Y(n66124) );
  XNOR2X1 U68568 ( .A(n65055), .B(n41671), .Y(n64782) );
  NOR2X1 U68569 ( .A(n41802), .B(n65385), .Y(n64779) );
  NAND2X1 U68570 ( .A(n64779), .B(n64778), .Y(n64780) );
  NAND2X1 U68571 ( .A(n64781), .B(n64780), .Y(n65081) );
  INVX1 U68572 ( .A(n65081), .Y(n65046) );
  XNOR2X1 U68573 ( .A(n64782), .B(n65046), .Y(n64792) );
  INVX1 U68574 ( .A(n64792), .Y(n64783) );
  NAND2X1 U68575 ( .A(n64784), .B(n64783), .Y(n64791) );
  NOR2X1 U68576 ( .A(n64792), .B(n64793), .Y(n64789) );
  INVX1 U68577 ( .A(n39613), .Y(n64785) );
  NOR2X1 U68578 ( .A(n64785), .B(n65058), .Y(n64787) );
  NAND2X1 U68579 ( .A(n64787), .B(n64786), .Y(n64788) );
  NAND2X1 U68580 ( .A(n64789), .B(n64788), .Y(n64790) );
  NAND2X1 U68581 ( .A(n64791), .B(n64790), .Y(n65037) );
  NAND2X1 U68582 ( .A(n65059), .B(n65058), .Y(n65056) );
  NAND2X1 U68583 ( .A(n65056), .B(n64792), .Y(n64803) );
  NOR2X1 U68584 ( .A(n64794), .B(n64793), .Y(n64796) );
  NAND2X1 U68585 ( .A(n64796), .B(n64795), .Y(n64801) );
  NAND2X1 U68586 ( .A(n65059), .B(n64799), .Y(n64800) );
  NAND2X1 U68587 ( .A(n64801), .B(n64800), .Y(n64802) );
  NOR2X1 U68588 ( .A(n64803), .B(n64802), .Y(n64805) );
  NAND2X1 U68589 ( .A(n65058), .B(n64804), .Y(n65053) );
  NOR2X1 U68590 ( .A(n65037), .B(n37397), .Y(n64806) );
  XNOR2X1 U68591 ( .A(n64807), .B(n65087), .Y(n65031) );
  NAND2X1 U68592 ( .A(n43492), .B(n43871), .Y(n65023) );
  XNOR2X1 U68593 ( .A(n65014), .B(n65009), .Y(n64808) );
  XNOR2X1 U68594 ( .A(n65035), .B(n64808), .Y(n64809) );
  XNOR2X1 U68595 ( .A(n64810), .B(n64809), .Y(n65006) );
  NOR2X1 U68596 ( .A(n64811), .B(n64997), .Y(n64813) );
  INVX1 U68597 ( .A(n64811), .Y(n64996) );
  INVX1 U68598 ( .A(n64997), .Y(n64814) );
  NAND2X1 U68599 ( .A(n43889), .B(n43484), .Y(n65001) );
  XOR2X1 U68600 ( .A(n65005), .B(n65001), .Y(n64815) );
  XNOR2X1 U68601 ( .A(n65006), .B(n64815), .Y(n65110) );
  NAND2X1 U68602 ( .A(n64818), .B(n64819), .Y(n64984) );
  INVX1 U68603 ( .A(n64819), .Y(n64821) );
  NAND2X1 U68604 ( .A(n64821), .B(n64820), .Y(n64822) );
  NAND2X1 U68605 ( .A(n64822), .B(n64823), .Y(n64986) );
  NAND2X1 U68606 ( .A(n64984), .B(n64986), .Y(n64990) );
  XNOR2X1 U68607 ( .A(n65336), .B(n39146), .Y(n64833) );
  NAND2X1 U68608 ( .A(n65338), .B(n65337), .Y(n64831) );
  NAND2X1 U68609 ( .A(n64826), .B(n64825), .Y(n64827) );
  NAND2X1 U68610 ( .A(n64827), .B(n65122), .Y(n64829) );
  NAND2X1 U68611 ( .A(n64829), .B(n64828), .Y(n64830) );
  NAND2X1 U68612 ( .A(n64831), .B(n64830), .Y(n64832) );
  INVX1 U68613 ( .A(n65338), .Y(n65334) );
  NAND2X1 U68614 ( .A(n64832), .B(n65326), .Y(n65119) );
  INVX1 U68615 ( .A(n64839), .Y(n64834) );
  NOR2X1 U68616 ( .A(n64834), .B(n64835), .Y(n64837) );
  NOR2X1 U68617 ( .A(n38564), .B(n64835), .Y(n64836) );
  NOR2X1 U68618 ( .A(n64837), .B(n64836), .Y(n64841) );
  NAND2X1 U68619 ( .A(n64839), .B(n64838), .Y(n64840) );
  NAND2X1 U68620 ( .A(n64841), .B(n64840), .Y(n65139) );
  INVX1 U68621 ( .A(n64842), .Y(n64845) );
  NOR2X1 U68622 ( .A(n41090), .B(n41145), .Y(n64846) );
  NAND2X1 U68623 ( .A(n64845), .B(n64844), .Y(n65142) );
  NAND2X1 U68624 ( .A(n64846), .B(n65142), .Y(n65845) );
  NAND2X1 U68625 ( .A(n43798), .B(n43934), .Y(n66179) );
  NAND2X1 U68626 ( .A(n43772), .B(n43943), .Y(n64979) );
  NOR2X1 U68627 ( .A(n64848), .B(n64847), .Y(n64849) );
  NOR2X1 U68628 ( .A(n64850), .B(n64849), .Y(n64854) );
  NAND2X1 U68629 ( .A(n38373), .B(n64852), .Y(n64853) );
  NAND2X1 U68630 ( .A(n36740), .B(n64853), .Y(n64981) );
  NAND2X1 U68631 ( .A(n43724), .B(n43983), .Y(n65474) );
  XNOR2X1 U68632 ( .A(n65474), .B(n42005), .Y(n64855) );
  INVX1 U68633 ( .A(n64856), .Y(n65489) );
  NOR2X1 U68634 ( .A(n64858), .B(n64857), .Y(n64860) );
  INVX1 U68635 ( .A(n64863), .Y(n64866) );
  NAND2X1 U68636 ( .A(n41602), .B(n41609), .Y(n65488) );
  NAND2X1 U68637 ( .A(n65489), .B(n65488), .Y(n65486) );
  XNOR2X1 U68638 ( .A(n64864), .B(n41999), .Y(n64865) );
  XNOR2X1 U68639 ( .A(n64866), .B(n64865), .Y(n65158) );
  XNOR2X1 U68640 ( .A(n65168), .B(n41130), .Y(n65278) );
  NAND2X1 U68641 ( .A(n40463), .B(n44018), .Y(n65504) );
  NAND2X1 U68642 ( .A(n40470), .B(n44009), .Y(n64932) );
  INVX1 U68643 ( .A(n64932), .Y(n65279) );
  XNOR2X1 U68644 ( .A(n65504), .B(n65279), .Y(n64867) );
  XNOR2X1 U68645 ( .A(n65270), .B(n64930), .Y(n64868) );
  XNOR2X1 U68646 ( .A(n65505), .B(n64868), .Y(n64869) );
  XNOR2X1 U68647 ( .A(n64870), .B(n36473), .Y(n64871) );
  XNOR2X1 U68648 ( .A(n40226), .B(n64871), .Y(n65178) );
  XNOR2X1 U68649 ( .A(n64872), .B(n65182), .Y(n64877) );
  NOR2X1 U68650 ( .A(n41079), .B(n64874), .Y(n64875) );
  NOR2X1 U68651 ( .A(n41371), .B(n64875), .Y(n64876) );
  XNOR2X1 U68652 ( .A(n64877), .B(n64876), .Y(n64910) );
  INVX1 U68653 ( .A(n64910), .Y(n64914) );
  XNOR2X1 U68654 ( .A(n43655), .B(n41153), .Y(n64879) );
  INVX1 U68655 ( .A(n64881), .Y(n64880) );
  NAND2X1 U68656 ( .A(n64880), .B(n43648), .Y(n64912) );
  NAND2X1 U68657 ( .A(n39446), .B(n64881), .Y(n64878) );
  NAND2X1 U68658 ( .A(n41365), .B(n64878), .Y(n64911) );
  XNOR2X1 U68659 ( .A(n64879), .B(n41158), .Y(n64883) );
  NAND2X1 U68660 ( .A(n43653), .B(n64881), .Y(n64882) );
  XNOR2X1 U68661 ( .A(n64908), .B(n43524), .Y(n64887) );
  NAND2X1 U68662 ( .A(n43521), .B(n64886), .Y(n65232) );
  NAND2X1 U68663 ( .A(n65234), .B(n65232), .Y(n64907) );
  XNOR2X1 U68664 ( .A(n64905), .B(n43679), .Y(n64888) );
  XNOR2X1 U68665 ( .A(n65203), .B(n43509), .Y(n64889) );
  XNOR2X1 U68666 ( .A(n41222), .B(n64889), .Y(n65205) );
  XNOR2X1 U68667 ( .A(n65205), .B(n43693), .Y(n64894) );
  NAND2X1 U68668 ( .A(n64890), .B(n43700), .Y(n65220) );
  NAND2X1 U68669 ( .A(n41454), .B(n64891), .Y(n64893) );
  NAND2X1 U68670 ( .A(n64893), .B(n64892), .Y(n65219) );
  NAND2X1 U68671 ( .A(n65220), .B(n65219), .Y(n65206) );
  XNOR2X1 U68672 ( .A(n64903), .B(n43708), .Y(n64895) );
  XNOR2X1 U68673 ( .A(n64896), .B(n64895), .Y(n64901) );
  XNOR2X1 U68674 ( .A(n64898), .B(n64897), .Y(n64899) );
  XNOR2X1 U68675 ( .A(n64899), .B(n41928), .Y(n64900) );
  MX2X1 U68676 ( .A(n64901), .B(n64900), .S0(n43720), .Y(u_muldiv_result_r[8])
         );
  NAND2X1 U68677 ( .A(u_muldiv_mult_result_q[8]), .B(n44633), .Y(n14065) );
  INVX1 U68678 ( .A(n64903), .Y(n64902) );
  NAND2X1 U68679 ( .A(n43705), .B(n64902), .Y(n65569) );
  NAND2X1 U68680 ( .A(n65569), .B(n65568), .Y(n65212) );
  NAND2X1 U68681 ( .A(n64905), .B(n43685), .Y(n65558) );
  NAND2X1 U68682 ( .A(n65558), .B(n64904), .Y(n65598) );
  INVX1 U68683 ( .A(n64905), .Y(n64906) );
  NAND2X1 U68684 ( .A(n43676), .B(n64906), .Y(n65554) );
  NAND2X1 U68685 ( .A(n65598), .B(n65554), .Y(n65202) );
  NAND2X1 U68686 ( .A(n64907), .B(n65233), .Y(n64909) );
  NAND2X1 U68687 ( .A(n43521), .B(n64908), .Y(n65229) );
  NAND2X1 U68688 ( .A(n64909), .B(n65229), .Y(n65552) );
  NAND2X1 U68689 ( .A(n40142), .B(n64910), .Y(n65924) );
  INVX1 U68690 ( .A(n64912), .Y(n64913) );
  NOR2X1 U68691 ( .A(n39475), .B(n64913), .Y(n64916) );
  NAND2X1 U68692 ( .A(n64914), .B(n43650), .Y(n64915) );
  NAND2X1 U68693 ( .A(n64916), .B(n64915), .Y(n65925) );
  XNOR2X1 U68694 ( .A(n43655), .B(n41105), .Y(n65195) );
  XNOR2X1 U68695 ( .A(n64917), .B(n36473), .Y(n64918) );
  XNOR2X1 U68696 ( .A(n40226), .B(n64918), .Y(n64922) );
  INVX1 U68697 ( .A(n64922), .Y(n64920) );
  NAND2X1 U68698 ( .A(n64920), .B(n64919), .Y(n64921) );
  NAND2X1 U68699 ( .A(n65251), .B(n64924), .Y(n64927) );
  NAND2X1 U68700 ( .A(n64929), .B(n64925), .Y(n64926) );
  OR2X1 U68701 ( .A(n64927), .B(n64926), .Y(n65260) );
  NAND2X1 U68702 ( .A(n36473), .B(n65252), .Y(n65262) );
  NAND2X1 U68703 ( .A(n65522), .B(n65523), .Y(n65172) );
  XNOR2X1 U68704 ( .A(n36727), .B(n64930), .Y(n65272) );
  NOR2X1 U68705 ( .A(n65272), .B(n39147), .Y(n64931) );
  NAND2X1 U68706 ( .A(n43821), .B(n44056), .Y(n65250) );
  INVX1 U68707 ( .A(n65250), .Y(n65257) );
  NAND2X1 U68708 ( .A(n36703), .B(n64932), .Y(n64945) );
  INVX1 U68709 ( .A(n64933), .Y(n64935) );
  NOR2X1 U68710 ( .A(n64935), .B(n64317), .Y(n64940) );
  NAND2X1 U68711 ( .A(n43995), .B(n64936), .Y(n64937) );
  NAND2X1 U68712 ( .A(n64938), .B(n64937), .Y(n64939) );
  NOR2X1 U68713 ( .A(n64940), .B(n64939), .Y(n64941) );
  NOR2X1 U68714 ( .A(n37383), .B(n64941), .Y(n64943) );
  NAND2X1 U68715 ( .A(n64943), .B(n64942), .Y(n64944) );
  NAND2X1 U68716 ( .A(n64945), .B(n64944), .Y(n65627) );
  NAND2X1 U68717 ( .A(n65279), .B(n65278), .Y(n65615) );
  NAND2X1 U68718 ( .A(n40483), .B(n44008), .Y(n65512) );
  INVX1 U68719 ( .A(n65474), .Y(n64958) );
  XNOR2X1 U68720 ( .A(n65475), .B(n64958), .Y(n64947) );
  XNOR2X1 U68721 ( .A(n38583), .B(n64947), .Y(n64948) );
  NOR2X1 U68722 ( .A(n43977), .B(n64950), .Y(n64951) );
  NOR2X1 U68723 ( .A(n64952), .B(n64951), .Y(n64956) );
  NAND2X1 U68724 ( .A(n40361), .B(n38623), .Y(n64955) );
  NAND2X1 U68725 ( .A(n64955), .B(n64956), .Y(n64957) );
  NOR2X1 U68726 ( .A(n65475), .B(n65474), .Y(n64959) );
  NOR2X1 U68727 ( .A(n41306), .B(n64959), .Y(n64965) );
  INVX1 U68728 ( .A(n65475), .Y(n64963) );
  NOR2X1 U68729 ( .A(n41572), .B(n41579), .Y(n64961) );
  NAND2X1 U68730 ( .A(n64961), .B(n64960), .Y(n64962) );
  NAND2X1 U68731 ( .A(n64963), .B(n64962), .Y(n64964) );
  NAND2X1 U68732 ( .A(n64965), .B(n64964), .Y(n65480) );
  NAND2X1 U68733 ( .A(n43787), .B(n44001), .Y(n65289) );
  INVX1 U68734 ( .A(n64966), .Y(n64976) );
  NOR2X1 U68735 ( .A(n43948), .B(n64967), .Y(n64969) );
  NOR2X1 U68736 ( .A(n43948), .B(n64970), .Y(n64968) );
  NOR2X1 U68737 ( .A(n64969), .B(n64968), .Y(n64974) );
  INVX1 U68738 ( .A(n64970), .Y(n64971) );
  NAND2X1 U68739 ( .A(n64972), .B(n64971), .Y(n64973) );
  NAND2X1 U68740 ( .A(n64974), .B(n64973), .Y(n64975) );
  NAND2X1 U68741 ( .A(n64978), .B(n64977), .Y(n65645) );
  NAND2X1 U68742 ( .A(n42632), .B(n43983), .Y(n65656) );
  INVX1 U68743 ( .A(n65656), .Y(n65470) );
  XNOR2X1 U68744 ( .A(n37319), .B(n65470), .Y(n65152) );
  INVX1 U68745 ( .A(n64979), .Y(n64980) );
  NAND2X1 U68746 ( .A(n64982), .B(n64981), .Y(n65293) );
  NAND2X1 U68747 ( .A(n42657), .B(n43934), .Y(n65305) );
  INVX1 U68748 ( .A(n64983), .Y(n64991) );
  INVX1 U68749 ( .A(n64984), .Y(n64985) );
  NOR2X1 U68750 ( .A(n64991), .B(n64985), .Y(n64987) );
  NAND2X1 U68751 ( .A(n64987), .B(n64986), .Y(n64988) );
  NAND2X1 U68752 ( .A(n64989), .B(n64988), .Y(n65452) );
  NAND2X1 U68753 ( .A(n64991), .B(n64990), .Y(n65451) );
  NAND2X1 U68754 ( .A(n64993), .B(n64992), .Y(n65355) );
  INVX1 U68755 ( .A(n65355), .Y(n64994) );
  NOR2X1 U68756 ( .A(n64995), .B(n64994), .Y(n65116) );
  NOR2X1 U68757 ( .A(n38673), .B(n38696), .Y(n64998) );
  NOR2X1 U68758 ( .A(n64997), .B(n64998), .Y(n64999) );
  NOR2X1 U68759 ( .A(n40947), .B(n64999), .Y(n65000) );
  NOR2X1 U68760 ( .A(n65000), .B(n65001), .Y(n65004) );
  INVX1 U68761 ( .A(n65006), .Y(n65002) );
  NOR2X1 U68762 ( .A(n65002), .B(n65001), .Y(n65003) );
  NOR2X1 U68763 ( .A(n65004), .B(n65003), .Y(n65008) );
  NAND2X1 U68764 ( .A(n65006), .B(n65005), .Y(n65007) );
  NAND2X1 U68765 ( .A(n65008), .B(n65007), .Y(n65361) );
  NAND2X1 U68766 ( .A(n43896), .B(n43483), .Y(n65359) );
  NAND2X1 U68767 ( .A(n65011), .B(n40272), .Y(n65013) );
  NOR2X1 U68768 ( .A(n40985), .B(n39109), .Y(n65022) );
  NAND2X1 U68769 ( .A(n65017), .B(n65016), .Y(n65018) );
  OR2X1 U68770 ( .A(n65019), .B(n65018), .Y(n65020) );
  NAND2X1 U68771 ( .A(n37408), .B(n65020), .Y(n65021) );
  NAND2X1 U68772 ( .A(n38672), .B(n65371), .Y(n65368) );
  INVX1 U68773 ( .A(n65023), .Y(n65032) );
  NAND2X1 U68774 ( .A(n65032), .B(n39819), .Y(n65024) );
  NOR2X1 U68775 ( .A(n40973), .B(n65024), .Y(n65030) );
  NAND2X1 U68776 ( .A(n65032), .B(n41508), .Y(n65027) );
  NOR2X1 U68777 ( .A(n65028), .B(n65027), .Y(n65029) );
  NOR2X1 U68778 ( .A(n65030), .B(n65029), .Y(n65034) );
  NAND2X1 U68779 ( .A(n65032), .B(n65036), .Y(n65033) );
  NAND2X1 U68780 ( .A(n65034), .B(n65033), .Y(n65366) );
  NOR2X1 U68781 ( .A(n65429), .B(n65413), .Y(n65038) );
  NOR2X1 U68782 ( .A(n65038), .B(n65416), .Y(n65432) );
  NAND2X1 U68783 ( .A(n65039), .B(n64744), .Y(n65428) );
  INVX1 U68784 ( .A(n65040), .Y(n65041) );
  NOR2X1 U68785 ( .A(n65042), .B(n65041), .Y(n65044) );
  NAND2X1 U68786 ( .A(n65044), .B(n65043), .Y(n65414) );
  INVX1 U68787 ( .A(n65414), .Y(n65430) );
  NAND2X1 U68788 ( .A(n65431), .B(n65430), .Y(n65045) );
  NAND2X1 U68789 ( .A(n65432), .B(n65045), .Y(n65763) );
  NAND2X1 U68790 ( .A(n65429), .B(n65086), .Y(n65762) );
  NAND2X1 U68791 ( .A(n43492), .B(n43880), .Y(n65737) );
  XNOR2X1 U68792 ( .A(n41671), .B(n65046), .Y(n65402) );
  NAND2X1 U68793 ( .A(n65064), .B(n65049), .Y(n65050) );
  NOR2X1 U68794 ( .A(n64412), .B(n65050), .Y(n65051) );
  NAND2X1 U68795 ( .A(n65051), .B(n39613), .Y(n65052) );
  NAND2X1 U68796 ( .A(n65059), .B(n65052), .Y(n65054) );
  NAND2X1 U68797 ( .A(n65054), .B(n65053), .Y(n65399) );
  NAND2X1 U68798 ( .A(n65402), .B(n65399), .Y(n65073) );
  INVX1 U68799 ( .A(n65055), .Y(n65072) );
  INVX1 U68800 ( .A(n65056), .Y(n65057) );
  NOR2X1 U68801 ( .A(n65402), .B(n65057), .Y(n65071) );
  NOR2X1 U68802 ( .A(n65059), .B(n65058), .Y(n65063) );
  INVX1 U68803 ( .A(n65064), .Y(n65061) );
  NOR2X1 U68804 ( .A(n65061), .B(n65060), .Y(n65062) );
  NOR2X1 U68805 ( .A(n65063), .B(n65062), .Y(n65069) );
  NAND2X1 U68806 ( .A(n65065), .B(n65064), .Y(n65066) );
  OR2X1 U68807 ( .A(n65067), .B(n65066), .Y(n65068) );
  NAND2X1 U68808 ( .A(n65069), .B(n65068), .Y(n65070) );
  NAND2X1 U68809 ( .A(n65071), .B(n65070), .Y(n65389) );
  NAND2X1 U68810 ( .A(n65072), .B(n65389), .Y(n65778) );
  NAND2X1 U68811 ( .A(n65073), .B(n65778), .Y(n65084) );
  NAND2X1 U68812 ( .A(n43962), .B(n39961), .Y(n65391) );
  NAND2X1 U68813 ( .A(n43859), .B(n43608), .Y(n65378) );
  NAND2X1 U68814 ( .A(n41490), .B(n43605), .Y(n65773) );
  INVX1 U68815 ( .A(n65773), .Y(n65074) );
  XNOR2X1 U68816 ( .A(n66132), .B(n65074), .Y(n65076) );
  XNOR2X1 U68817 ( .A(n65076), .B(n65075), .Y(n65080) );
  NAND2X1 U68818 ( .A(n65077), .B(n66132), .Y(n65079) );
  NAND2X1 U68819 ( .A(n66132), .B(n65078), .Y(n65382) );
  NAND2X1 U68820 ( .A(n65079), .B(n65382), .Y(n65772) );
  INVX1 U68821 ( .A(n65379), .Y(n65392) );
  NAND2X1 U68822 ( .A(n65081), .B(n66124), .Y(n65082) );
  NAND2X1 U68823 ( .A(n41490), .B(n65082), .Y(n65390) );
  XNOR2X1 U68824 ( .A(n65391), .B(n65388), .Y(n65083) );
  XNOR2X1 U68825 ( .A(n65084), .B(n65083), .Y(n65754) );
  NAND2X1 U68826 ( .A(n43952), .B(n43501), .Y(n65761) );
  NAND2X1 U68827 ( .A(n43870), .B(n43497), .Y(n65792) );
  XNOR2X1 U68828 ( .A(n65737), .B(n65373), .Y(n65085) );
  XNOR2X1 U68829 ( .A(n39129), .B(n65085), .Y(n65096) );
  NAND2X1 U68830 ( .A(n41221), .B(n65088), .Y(n65436) );
  NOR2X1 U68831 ( .A(n37391), .B(n41221), .Y(n65094) );
  INVX1 U68832 ( .A(n65089), .Y(n65092) );
  NAND2X1 U68833 ( .A(n40996), .B(n65090), .Y(n65091) );
  NAND2X1 U68834 ( .A(n65092), .B(n65091), .Y(n65093) );
  NAND2X1 U68835 ( .A(n65094), .B(n65093), .Y(n65095) );
  NAND2X1 U68836 ( .A(n41507), .B(n65095), .Y(n65435) );
  XNOR2X1 U68837 ( .A(n65096), .B(n40998), .Y(n65363) );
  NAND2X1 U68838 ( .A(n43889), .B(n38310), .Y(n65369) );
  XNOR2X1 U68839 ( .A(n65363), .B(n65369), .Y(n65097) );
  NAND2X1 U68840 ( .A(n65110), .B(n65098), .Y(n65346) );
  INVX1 U68841 ( .A(n65346), .Y(n65695) );
  INVX1 U68842 ( .A(n65099), .Y(n65111) );
  NAND2X1 U68843 ( .A(n65102), .B(n38867), .Y(n65103) );
  NAND2X1 U68844 ( .A(n65104), .B(n65103), .Y(n65108) );
  NAND2X1 U68845 ( .A(n65106), .B(n65105), .Y(n65107) );
  NAND2X1 U68846 ( .A(n65108), .B(n65107), .Y(n65109) );
  NAND2X1 U68847 ( .A(n65111), .B(n65109), .Y(n65347) );
  INVX1 U68848 ( .A(n65347), .Y(n65694) );
  NAND2X1 U68849 ( .A(n43909), .B(n43775), .Y(n66041) );
  NAND2X1 U68850 ( .A(n43903), .B(n43478), .Y(n65707) );
  INVX1 U68851 ( .A(n65707), .Y(n65699) );
  XNOR2X1 U68852 ( .A(n66041), .B(n65699), .Y(n65113) );
  XNOR2X1 U68853 ( .A(n39016), .B(n65113), .Y(n65114) );
  XNOR2X1 U68854 ( .A(n65708), .B(n65114), .Y(n65115) );
  XNOR2X1 U68855 ( .A(n65116), .B(n65115), .Y(n65450) );
  NAND2X1 U68856 ( .A(n43918), .B(n43796), .Y(n65449) );
  NAND2X1 U68857 ( .A(n43927), .B(n42711), .Y(n65341) );
  INVX1 U68858 ( .A(n65341), .Y(n65323) );
  XNOR2X1 U68859 ( .A(n65449), .B(n65323), .Y(n65117) );
  XNOR2X1 U68860 ( .A(n65450), .B(n65117), .Y(n65118) );
  INVX1 U68861 ( .A(n65315), .Y(n65121) );
  INVX1 U68862 ( .A(n65119), .Y(n65120) );
  NOR2X1 U68863 ( .A(n65121), .B(n65120), .Y(n65134) );
  INVX1 U68864 ( .A(n65122), .Y(n65126) );
  NOR2X1 U68865 ( .A(n65124), .B(n65123), .Y(n65125) );
  NOR2X1 U68866 ( .A(n65126), .B(n65125), .Y(n65127) );
  NOR2X1 U68867 ( .A(n39101), .B(n65127), .Y(n65128) );
  NAND2X1 U68868 ( .A(n65128), .B(n65338), .Y(n65129) );
  NAND2X1 U68869 ( .A(n65312), .B(n65129), .Y(n65317) );
  NAND2X1 U68870 ( .A(n36702), .B(n65130), .Y(n65333) );
  NAND2X1 U68871 ( .A(n65333), .B(n65334), .Y(n65318) );
  NAND2X1 U68872 ( .A(n65317), .B(n65318), .Y(n65131) );
  NOR2X1 U68873 ( .A(n65315), .B(n65131), .Y(n65132) );
  NOR2X1 U68874 ( .A(n65132), .B(n65336), .Y(n65133) );
  NOR2X1 U68875 ( .A(n65134), .B(n65133), .Y(n65303) );
  NOR2X1 U68876 ( .A(n65138), .B(n65135), .Y(n65136) );
  INVX1 U68877 ( .A(n65138), .Y(n65140) );
  INVX1 U68878 ( .A(n65307), .Y(n65295) );
  XNOR2X1 U68879 ( .A(n41435), .B(n65295), .Y(n65465) );
  NAND2X1 U68880 ( .A(n43772), .B(n43973), .Y(n65294) );
  INVX1 U68881 ( .A(n65294), .Y(n65665) );
  NAND2X1 U68882 ( .A(n43799), .B(n43943), .Y(n66183) );
  INVX1 U68883 ( .A(n66183), .Y(n65466) );
  XNOR2X1 U68884 ( .A(n65665), .B(n65466), .Y(n65149) );
  INVX1 U68885 ( .A(n66180), .Y(n65141) );
  NOR2X1 U68886 ( .A(n65141), .B(n66179), .Y(n65148) );
  NOR2X1 U68887 ( .A(n41090), .B(n41145), .Y(n65143) );
  NAND2X1 U68888 ( .A(n65143), .B(n65142), .Y(n65144) );
  NAND2X1 U68889 ( .A(n65144), .B(n66180), .Y(n65146) );
  OR2X1 U68890 ( .A(n38556), .B(n66179), .Y(n65145) );
  NAND2X1 U68891 ( .A(n65146), .B(n65145), .Y(n65147) );
  NOR2X1 U68892 ( .A(n65148), .B(n65147), .Y(n65298) );
  XNOR2X1 U68893 ( .A(n65149), .B(n65298), .Y(n65150) );
  XNOR2X1 U68894 ( .A(n65465), .B(n65150), .Y(n65151) );
  INVX1 U68895 ( .A(n65478), .Y(n65655) );
  XNOR2X1 U68896 ( .A(n65289), .B(n65287), .Y(n65153) );
  NAND2X1 U68897 ( .A(n65163), .B(n65490), .Y(n65162) );
  NAND2X1 U68898 ( .A(n41602), .B(n41609), .Y(n65156) );
  NAND2X1 U68899 ( .A(n65489), .B(n65156), .Y(n65160) );
  NAND2X1 U68900 ( .A(n65158), .B(n65157), .Y(n65159) );
  NAND2X1 U68901 ( .A(n65160), .B(n65159), .Y(n65161) );
  NAND2X1 U68902 ( .A(n65162), .B(n65161), .Y(n65165) );
  OR2X1 U68903 ( .A(n65490), .B(n65163), .Y(n65164) );
  NAND2X1 U68904 ( .A(n65165), .B(n65164), .Y(n65497) );
  INVX1 U68905 ( .A(n65497), .Y(n65510) );
  XNOR2X1 U68906 ( .A(n65513), .B(n65510), .Y(n65630) );
  INVX1 U68907 ( .A(n65630), .Y(n65530) );
  XNOR2X1 U68908 ( .A(n65619), .B(n65530), .Y(n65167) );
  NAND2X1 U68909 ( .A(n40471), .B(n44018), .Y(n65620) );
  NAND2X1 U68910 ( .A(n40464), .B(n44026), .Y(n65509) );
  XNOR2X1 U68911 ( .A(n65620), .B(n65509), .Y(n65166) );
  XNOR2X1 U68912 ( .A(n65167), .B(n65166), .Y(n65254) );
  INVX1 U68913 ( .A(n65504), .Y(n65527) );
  XNOR2X1 U68914 ( .A(n65168), .B(n65279), .Y(n65169) );
  XNOR2X1 U68915 ( .A(n65169), .B(n41130), .Y(n65170) );
  NAND2X1 U68916 ( .A(n65527), .B(n65171), .Y(n65173) );
  INVX1 U68917 ( .A(n65524), .Y(n65506) );
  AND2X1 U68918 ( .A(n65173), .B(n38929), .Y(n65255) );
  XNOR2X1 U68919 ( .A(n65254), .B(n65255), .Y(n65269) );
  XNOR2X1 U68920 ( .A(n38515), .B(n65174), .Y(n65247) );
  NAND2X1 U68921 ( .A(n43612), .B(n43759), .Y(n72153) );
  XNOR2X1 U68922 ( .A(n65247), .B(n43546), .Y(n65175) );
  XNOR2X1 U68923 ( .A(n41342), .B(n65175), .Y(n65243) );
  XNOR2X1 U68924 ( .A(n43639), .B(n65243), .Y(n65176) );
  XOR2X1 U68925 ( .A(n66519), .B(n65176), .Y(n65540) );
  XNOR2X1 U68926 ( .A(n43666), .B(n65540), .Y(n65181) );
  NAND2X1 U68927 ( .A(n65180), .B(n43636), .Y(n65903) );
  INVX1 U68928 ( .A(n65244), .Y(n65539) );
  XNOR2X1 U68929 ( .A(n65181), .B(n65539), .Y(n65194) );
  NOR2X1 U68930 ( .A(n43666), .B(n65192), .Y(n65184) );
  NOR2X1 U68931 ( .A(n41371), .B(n65184), .Y(n65191) );
  NOR2X1 U68932 ( .A(n37359), .B(n41079), .Y(n65189) );
  NAND2X1 U68933 ( .A(n40025), .B(n65185), .Y(n65186) );
  NAND2X1 U68934 ( .A(n65187), .B(n65186), .Y(n65188) );
  NAND2X1 U68935 ( .A(n65188), .B(n65189), .Y(n65190) );
  AND2X1 U68936 ( .A(n65191), .B(n65190), .Y(n65538) );
  NOR2X1 U68937 ( .A(n65538), .B(n41098), .Y(n65193) );
  XNOR2X1 U68938 ( .A(n65193), .B(n65194), .Y(n65547) );
  INVX1 U68939 ( .A(n65547), .Y(n65546) );
  XNOR2X1 U68940 ( .A(n65195), .B(n41108), .Y(n65200) );
  XNOR2X1 U68941 ( .A(n41153), .B(n41158), .Y(n65196) );
  NOR2X1 U68942 ( .A(n37927), .B(n65197), .Y(n65198) );
  NOR2X1 U68943 ( .A(n41184), .B(n65198), .Y(n65199) );
  XNOR2X1 U68944 ( .A(n65200), .B(n65199), .Y(n65553) );
  XNOR2X1 U68945 ( .A(n43677), .B(n43524), .Y(n71402) );
  XNOR2X1 U68946 ( .A(n65202), .B(n65201), .Y(n65226) );
  NAND2X1 U68947 ( .A(n43505), .B(n65203), .Y(n65588) );
  INVX1 U68948 ( .A(n65203), .Y(n65204) );
  XNOR2X1 U68949 ( .A(n65223), .B(n43693), .Y(n65210) );
  NAND2X1 U68950 ( .A(n65205), .B(n43701), .Y(n65221) );
  INVX1 U68951 ( .A(n65221), .Y(n65207) );
  NOR2X1 U68952 ( .A(n65207), .B(n65206), .Y(n65208) );
  NOR2X1 U68953 ( .A(n41226), .B(n65208), .Y(n65209) );
  XNOR2X1 U68954 ( .A(n65210), .B(n65209), .Y(n65570) );
  XNOR2X1 U68955 ( .A(n65570), .B(n43708), .Y(n65211) );
  XNOR2X1 U68956 ( .A(n65212), .B(n65211), .Y(n65217) );
  XNOR2X1 U68957 ( .A(n65214), .B(n65213), .Y(n65215) );
  XNOR2X1 U68958 ( .A(n41940), .B(n65215), .Y(n65216) );
  MX2X1 U68959 ( .A(n65217), .B(n65216), .S0(n43720), .Y(u_muldiv_result_r[9])
         );
  NAND2X1 U68960 ( .A(u_muldiv_mult_result_q[9]), .B(n44633), .Y(n14054) );
  NOR2X1 U68961 ( .A(n43702), .B(n65223), .Y(n65218) );
  NAND2X1 U68962 ( .A(n65223), .B(n43700), .Y(n65224) );
  NAND2X1 U68963 ( .A(n65226), .B(n43512), .Y(n65592) );
  NAND2X1 U68964 ( .A(n65227), .B(n65586), .Y(n65228) );
  NAND2X1 U68965 ( .A(n65592), .B(n65228), .Y(n65565) );
  NAND2X1 U68966 ( .A(n65553), .B(n43529), .Y(n65238) );
  INVX1 U68967 ( .A(n65229), .Y(n65231) );
  NOR2X1 U68968 ( .A(n43532), .B(n65553), .Y(n65230) );
  INVX1 U68969 ( .A(n65232), .Y(n65236) );
  NOR2X1 U68970 ( .A(n40344), .B(n65234), .Y(n65235) );
  NAND2X1 U68971 ( .A(n65238), .B(n65237), .Y(n65603) );
  NOR2X1 U68972 ( .A(n37927), .B(n65239), .Y(n65242) );
  NOR2X1 U68973 ( .A(n40971), .B(n43661), .Y(n65240) );
  OR2X1 U68974 ( .A(n41184), .B(n65240), .Y(n65241) );
  NOR2X1 U68975 ( .A(n65242), .B(n65241), .Y(n65931) );
  NOR2X1 U68976 ( .A(n65931), .B(n41398), .Y(n65551) );
  NAND2X1 U68977 ( .A(n65245), .B(n43638), .Y(n65899) );
  NAND2X1 U68978 ( .A(n65244), .B(n65899), .Y(n65246) );
  XNOR2X1 U68979 ( .A(n43666), .B(n41078), .Y(n65537) );
  INVX1 U68980 ( .A(n65249), .Y(n65248) );
  NAND2X1 U68981 ( .A(n65248), .B(n43548), .Y(n66516) );
  NAND2X1 U68982 ( .A(n66516), .B(n66519), .Y(n65910) );
  NAND2X1 U68983 ( .A(n43545), .B(n65249), .Y(n66514) );
  NAND2X1 U68984 ( .A(n66514), .B(n65910), .Y(n66219) );
  NOR2X1 U68985 ( .A(n65251), .B(n65250), .Y(n65253) );
  XNOR2X1 U68986 ( .A(n42067), .B(n65254), .Y(n65256) );
  NOR2X1 U68987 ( .A(n65259), .B(n65258), .Y(n65266) );
  NAND2X1 U68988 ( .A(n65261), .B(n65260), .Y(n65263) );
  NAND2X1 U68989 ( .A(n65263), .B(n65262), .Y(n65264) );
  NAND2X1 U68990 ( .A(n65264), .B(n41559), .Y(n65265) );
  NAND2X1 U68991 ( .A(n65266), .B(n65265), .Y(n65613) );
  NAND2X1 U68992 ( .A(n65269), .B(n65267), .Y(n65878) );
  INVX1 U68993 ( .A(n65270), .Y(n65276) );
  NOR2X1 U68994 ( .A(n65272), .B(n65271), .Y(n65274) );
  NAND2X1 U68995 ( .A(n65274), .B(n39947), .Y(n65275) );
  NAND2X1 U68996 ( .A(n42067), .B(n65876), .Y(n65277) );
  NAND2X1 U68997 ( .A(n65878), .B(n65277), .Y(n65880) );
  NAND2X1 U68998 ( .A(n40467), .B(n44049), .Y(n65977) );
  INVX1 U68999 ( .A(n65977), .Y(n65988) );
  NOR2X1 U69000 ( .A(n65279), .B(n65278), .Y(n65282) );
  INVX1 U69001 ( .A(n65615), .Y(n65626) );
  NOR2X1 U69002 ( .A(n65626), .B(n65280), .Y(n65281) );
  NOR2X1 U69003 ( .A(n65282), .B(n65281), .Y(n65283) );
  NOR2X1 U69004 ( .A(n65630), .B(n65283), .Y(n65284) );
  NOR2X1 U69005 ( .A(n65284), .B(n65620), .Y(n65286) );
  INVX1 U69006 ( .A(n65619), .Y(n65529) );
  NOR2X1 U69007 ( .A(n65529), .B(n65530), .Y(n65285) );
  NOR2X1 U69008 ( .A(n65286), .B(n65285), .Y(n65502) );
  INVX1 U69009 ( .A(n65289), .Y(n65291) );
  NAND2X1 U69010 ( .A(n65291), .B(n38491), .Y(n65292) );
  INVX1 U69011 ( .A(n36587), .Y(n65861) );
  XNOR2X1 U69012 ( .A(n65466), .B(n65295), .Y(n65296) );
  XNOR2X1 U69013 ( .A(n65296), .B(n41435), .Y(n65297) );
  NAND2X1 U69014 ( .A(n65299), .B(n36774), .Y(n65300) );
  NAND2X1 U69015 ( .A(n65665), .B(n36774), .Y(n65666) );
  NAND2X1 U69016 ( .A(n65300), .B(n65666), .Y(n65301) );
  NOR2X1 U69017 ( .A(n65302), .B(n65301), .Y(n65652) );
  NAND2X1 U69018 ( .A(n40259), .B(n43983), .Y(n65672) );
  INVX1 U69019 ( .A(n65672), .Y(n65664) );
  XNOR2X1 U69020 ( .A(n37320), .B(n65664), .Y(n65467) );
  XNOR2X1 U69021 ( .A(n65304), .B(n65303), .Y(n65306) );
  OR2X1 U69022 ( .A(n65306), .B(n65305), .Y(n65310) );
  NAND2X1 U69023 ( .A(n65306), .B(n65305), .Y(n65308) );
  NAND2X1 U69024 ( .A(n65308), .B(n65307), .Y(n65309) );
  NAND2X1 U69025 ( .A(n65310), .B(n65309), .Y(n65825) );
  NAND2X1 U69026 ( .A(n65326), .B(n65336), .Y(n65313) );
  NOR2X1 U69027 ( .A(n39384), .B(n65313), .Y(n65314) );
  NAND2X1 U69028 ( .A(n65314), .B(n65318), .Y(n65316) );
  NAND2X1 U69029 ( .A(n65316), .B(n65315), .Y(n65322) );
  INVX1 U69030 ( .A(n65336), .Y(n65320) );
  NAND2X1 U69031 ( .A(n65318), .B(n65317), .Y(n65319) );
  NAND2X1 U69032 ( .A(n65320), .B(n65319), .Y(n65321) );
  INVX1 U69033 ( .A(n65450), .Y(n65455) );
  INVX1 U69034 ( .A(n65449), .Y(n65456) );
  XNOR2X1 U69035 ( .A(n65453), .B(n65456), .Y(n65324) );
  XNOR2X1 U69036 ( .A(n65455), .B(n65324), .Y(n65829) );
  INVX1 U69037 ( .A(n65333), .Y(n65325) );
  NOR2X1 U69038 ( .A(n65338), .B(n65325), .Y(n65329) );
  NAND2X1 U69039 ( .A(n65327), .B(n65326), .Y(n65328) );
  NOR2X1 U69040 ( .A(n65329), .B(n65328), .Y(n65330) );
  NOR2X1 U69041 ( .A(n39146), .B(n65330), .Y(n65332) );
  NOR2X1 U69042 ( .A(n39146), .B(n65336), .Y(n65331) );
  NAND2X1 U69043 ( .A(n65334), .B(n65333), .Y(n65335) );
  NOR2X1 U69044 ( .A(n65336), .B(n65335), .Y(n65344) );
  NOR2X1 U69045 ( .A(n65337), .B(n65336), .Y(n65340) );
  NAND2X1 U69046 ( .A(n36709), .B(n65338), .Y(n65339) );
  NAND2X1 U69047 ( .A(n65340), .B(n65339), .Y(n65342) );
  NAND2X1 U69048 ( .A(n65342), .B(n65341), .Y(n65343) );
  NAND2X1 U69049 ( .A(n65834), .B(n65830), .Y(n66167) );
  NAND2X1 U69050 ( .A(n42658), .B(n43943), .Y(n65831) );
  NAND2X1 U69051 ( .A(n43799), .B(n43973), .Y(n65844) );
  INVX1 U69052 ( .A(n65844), .Y(n65843) );
  XNOR2X1 U69053 ( .A(n65831), .B(n65843), .Y(n65345) );
  XNOR2X1 U69054 ( .A(n39451), .B(n65345), .Y(n65460) );
  XNOR2X1 U69055 ( .A(n65708), .B(n65699), .Y(n65350) );
  NAND2X1 U69056 ( .A(n65347), .B(n65346), .Y(n65348) );
  NOR2X1 U69057 ( .A(n38600), .B(n65348), .Y(n65349) );
  XNOR2X1 U69058 ( .A(n65350), .B(n65349), .Y(n66044) );
  INVX1 U69059 ( .A(n66044), .Y(n65351) );
  NAND2X1 U69060 ( .A(n65351), .B(n66041), .Y(n65357) );
  INVX1 U69061 ( .A(n65352), .Y(n65354) );
  NAND2X1 U69062 ( .A(n65354), .B(n65353), .Y(n65356) );
  NAND2X1 U69063 ( .A(n65356), .B(n65355), .Y(n66043) );
  INVX1 U69064 ( .A(n66041), .Y(n65358) );
  NAND2X1 U69065 ( .A(n65360), .B(n40261), .Y(n65715) );
  INVX1 U69066 ( .A(n65359), .Y(n65362) );
  NAND2X1 U69067 ( .A(n65362), .B(n65360), .Y(n65716) );
  NAND2X1 U69068 ( .A(n65362), .B(n65361), .Y(n65717) );
  INVX1 U69069 ( .A(n65364), .Y(n65365) );
  NOR2X1 U69070 ( .A(n65366), .B(n65365), .Y(n65367) );
  NAND2X1 U69071 ( .A(n65370), .B(n65368), .Y(n65725) );
  NOR2X1 U69072 ( .A(n39479), .B(n65370), .Y(n65372) );
  NAND2X1 U69073 ( .A(n65725), .B(n65726), .Y(n65723) );
  NAND2X1 U69074 ( .A(n43903), .B(n43482), .Y(n66056) );
  INVX1 U69075 ( .A(n66056), .Y(n65720) );
  INVX1 U69076 ( .A(n65737), .Y(n65729) );
  XNOR2X1 U69077 ( .A(n39129), .B(n65373), .Y(n65374) );
  XNOR2X1 U69078 ( .A(n40998), .B(n65374), .Y(n65736) );
  NOR2X1 U69079 ( .A(n40478), .B(n65737), .Y(n65375) );
  NOR2X1 U69080 ( .A(n41000), .B(n65375), .Y(n65377) );
  NAND2X1 U69081 ( .A(n65736), .B(n65739), .Y(n65376) );
  NAND2X1 U69082 ( .A(n65377), .B(n65376), .Y(n65722) );
  NAND2X1 U69083 ( .A(n43896), .B(n38311), .Y(n65724) );
  NAND2X1 U69084 ( .A(n43492), .B(n43890), .Y(n65728) );
  INVX1 U69085 ( .A(n65378), .Y(n65381) );
  NAND2X1 U69086 ( .A(n65379), .B(n65390), .Y(n65380) );
  NAND2X1 U69087 ( .A(n65381), .B(n65380), .Y(n65780) );
  XNOR2X1 U69088 ( .A(n65780), .B(n41505), .Y(n65387) );
  NAND2X1 U69089 ( .A(n65381), .B(n43605), .Y(n65774) );
  NAND2X1 U69090 ( .A(n65382), .B(n65773), .Y(n65383) );
  OR2X1 U69091 ( .A(n66131), .B(n65383), .Y(n65384) );
  NOR2X1 U69092 ( .A(n65385), .B(n65384), .Y(n65386) );
  XNOR2X1 U69093 ( .A(n65387), .B(n41675), .Y(n65747) );
  NAND2X1 U69094 ( .A(n43869), .B(n43501), .Y(n65760) );
  INVX1 U69095 ( .A(n65760), .Y(n65769) );
  XNOR2X1 U69096 ( .A(n65747), .B(n65769), .Y(n65406) );
  INVX1 U69097 ( .A(n65391), .Y(n65401) );
  INVX1 U69098 ( .A(n65388), .Y(n65400) );
  NAND2X1 U69099 ( .A(n65401), .B(n65400), .Y(n65781) );
  INVX1 U69100 ( .A(n65781), .Y(n65398) );
  NOR2X1 U69101 ( .A(n65401), .B(n65390), .Y(n65395) );
  NAND2X1 U69102 ( .A(n65392), .B(n65391), .Y(n65393) );
  NAND2X1 U69103 ( .A(n65393), .B(n43517), .Y(n65394) );
  NOR2X1 U69104 ( .A(n65395), .B(n65394), .Y(n65396) );
  NOR2X1 U69105 ( .A(n65398), .B(n65397), .Y(n65405) );
  NAND2X1 U69106 ( .A(n65403), .B(n65402), .Y(n65404) );
  NAND2X1 U69107 ( .A(n65405), .B(n65404), .Y(n65786) );
  INVX1 U69108 ( .A(n65786), .Y(n65748) );
  XNOR2X1 U69109 ( .A(n65406), .B(n65748), .Y(n65409) );
  INVX1 U69110 ( .A(n65409), .Y(n65420) );
  INVX1 U69111 ( .A(n65754), .Y(n65749) );
  NAND2X1 U69112 ( .A(n65749), .B(n65761), .Y(n65407) );
  NOR2X1 U69113 ( .A(n65420), .B(n65407), .Y(n65411) );
  NAND2X1 U69114 ( .A(n65754), .B(n65764), .Y(n65408) );
  NOR2X1 U69115 ( .A(n65409), .B(n65408), .Y(n65410) );
  NOR2X1 U69116 ( .A(n65411), .B(n65410), .Y(n65427) );
  INVX1 U69117 ( .A(n65761), .Y(n65421) );
  NAND2X1 U69118 ( .A(n65421), .B(n65754), .Y(n65766) );
  NAND2X1 U69119 ( .A(n40005), .B(n65766), .Y(n65412) );
  NOR2X1 U69120 ( .A(n65420), .B(n65412), .Y(n65425) );
  NOR2X1 U69121 ( .A(n65415), .B(n65429), .Y(n65417) );
  NOR2X1 U69122 ( .A(n65417), .B(n65416), .Y(n65419) );
  NAND2X1 U69123 ( .A(n40313), .B(n65749), .Y(n65418) );
  NOR2X1 U69124 ( .A(n65419), .B(n65418), .Y(n65423) );
  NAND2X1 U69125 ( .A(n65421), .B(n65420), .Y(n65422) );
  NOR2X1 U69126 ( .A(n65423), .B(n65422), .Y(n65424) );
  NOR2X1 U69127 ( .A(n65425), .B(n65424), .Y(n65426) );
  NAND2X1 U69128 ( .A(n65427), .B(n65426), .Y(n65796) );
  NAND2X1 U69129 ( .A(n43879), .B(n43496), .Y(n65801) );
  INVX1 U69130 ( .A(n65801), .Y(n65804) );
  XNOR2X1 U69131 ( .A(n65728), .B(n40999), .Y(n65442) );
  NOR2X1 U69132 ( .A(n65429), .B(n65428), .Y(n65431) );
  NAND2X1 U69133 ( .A(n65432), .B(n65045), .Y(n65756) );
  NAND2X1 U69134 ( .A(n65756), .B(n40313), .Y(n65434) );
  XNOR2X1 U69135 ( .A(n65761), .B(n65754), .Y(n65433) );
  XNOR2X1 U69136 ( .A(n65434), .B(n65433), .Y(n65802) );
  NOR2X1 U69137 ( .A(n65802), .B(n65792), .Y(n65438) );
  NAND2X1 U69138 ( .A(n65436), .B(n65435), .Y(n65440) );
  NOR2X1 U69139 ( .A(n40998), .B(n65792), .Y(n65437) );
  NOR2X1 U69140 ( .A(n65438), .B(n65437), .Y(n65441) );
  INVX1 U69141 ( .A(n65802), .Y(n65439) );
  NAND2X1 U69142 ( .A(n65440), .B(n65439), .Y(n65795) );
  XNOR2X1 U69143 ( .A(n65442), .B(n41224), .Y(n65721) );
  XNOR2X1 U69144 ( .A(n65724), .B(n65721), .Y(n65443) );
  XOR2X1 U69145 ( .A(n65722), .B(n65443), .Y(n65713) );
  NAND2X1 U69146 ( .A(n43909), .B(n43478), .Y(n65693) );
  INVX1 U69147 ( .A(n65693), .Y(n65704) );
  NAND2X1 U69148 ( .A(n43918), .B(n43775), .Y(n66048) );
  INVX1 U69149 ( .A(n66048), .Y(n65690) );
  XNOR2X1 U69150 ( .A(n65704), .B(n65690), .Y(n65675) );
  NAND2X1 U69151 ( .A(n43927), .B(n43795), .Y(n65680) );
  INVX1 U69152 ( .A(n65680), .Y(n65679) );
  XNOR2X1 U69153 ( .A(n65675), .B(n65679), .Y(n65444) );
  XNOR2X1 U69154 ( .A(n40984), .B(n65444), .Y(n65447) );
  NOR2X1 U69155 ( .A(n37386), .B(n65708), .Y(n65446) );
  INVX1 U69156 ( .A(n65708), .Y(n65698) );
  NAND2X1 U69157 ( .A(n65699), .B(n65698), .Y(n65710) );
  XNOR2X1 U69158 ( .A(n65447), .B(n39113), .Y(n65448) );
  XNOR2X1 U69159 ( .A(n39117), .B(n65448), .Y(n65812) );
  NAND2X1 U69160 ( .A(n65450), .B(n65449), .Y(n65454) );
  NAND2X1 U69161 ( .A(n65452), .B(n65451), .Y(n65453) );
  NAND2X1 U69162 ( .A(n65454), .B(n65453), .Y(n65458) );
  NAND2X1 U69163 ( .A(n65456), .B(n65455), .Y(n65457) );
  NAND2X1 U69164 ( .A(n65458), .B(n65457), .Y(n65813) );
  XNOR2X1 U69165 ( .A(n65815), .B(n39013), .Y(n65459) );
  XOR2X1 U69166 ( .A(n65812), .B(n65459), .Y(n65840) );
  NOR2X1 U69167 ( .A(n38556), .B(n66179), .Y(n65461) );
  NOR2X1 U69168 ( .A(n65461), .B(n66180), .Y(n65462) );
  NOR2X1 U69169 ( .A(n41375), .B(n65462), .Y(n65464) );
  INVX1 U69170 ( .A(n65465), .Y(n66184) );
  NAND2X1 U69171 ( .A(n66184), .B(n66183), .Y(n65463) );
  NAND2X1 U69172 ( .A(n65466), .B(n65465), .Y(n66187) );
  XNOR2X1 U69173 ( .A(n41185), .B(n41376), .Y(n65671) );
  INVX1 U69174 ( .A(n65671), .Y(n65663) );
  XNOR2X1 U69175 ( .A(n65467), .B(n65663), .Y(n65468) );
  XNOR2X1 U69176 ( .A(n65652), .B(n65468), .Y(n65637) );
  NAND2X1 U69177 ( .A(n43724), .B(n44001), .Y(n66024) );
  INVX1 U69178 ( .A(n66024), .Y(n65639) );
  INVX1 U69179 ( .A(n65479), .Y(n65469) );
  NOR2X1 U69180 ( .A(n65469), .B(n65656), .Y(n65473) );
  NAND2X1 U69181 ( .A(n65470), .B(n65478), .Y(n65659) );
  NAND2X1 U69182 ( .A(n65478), .B(n65479), .Y(n65471) );
  NAND2X1 U69183 ( .A(n65659), .B(n65471), .Y(n65472) );
  NOR2X1 U69184 ( .A(n65473), .B(n65472), .Y(n65638) );
  NOR2X1 U69185 ( .A(n38583), .B(n65475), .Y(n65476) );
  OR2X1 U69186 ( .A(n41306), .B(n65476), .Y(n65477) );
  NOR2X1 U69187 ( .A(n41283), .B(n65640), .Y(n65482) );
  NAND2X1 U69188 ( .A(n65481), .B(n65480), .Y(n65641) );
  NAND2X1 U69189 ( .A(n65641), .B(n65482), .Y(n66025) );
  XNOR2X1 U69190 ( .A(n41362), .B(n40199), .Y(n66015) );
  NAND2X1 U69191 ( .A(n43787), .B(n44008), .Y(n66016) );
  NAND2X1 U69192 ( .A(n40482), .B(n44018), .Y(n66859) );
  INVX1 U69193 ( .A(n66859), .Y(n66008) );
  XNOR2X1 U69194 ( .A(n66016), .B(n66008), .Y(n65483) );
  XNOR2X1 U69195 ( .A(n66015), .B(n65483), .Y(n65484) );
  XNOR2X1 U69196 ( .A(n65861), .B(n65484), .Y(n65633) );
  INVX1 U69197 ( .A(n65512), .Y(n65485) );
  NOR2X1 U69198 ( .A(n65487), .B(n65512), .Y(n65496) );
  INVX1 U69199 ( .A(n65490), .Y(n65491) );
  NOR2X1 U69200 ( .A(n65492), .B(n65491), .Y(n65494) );
  NAND2X1 U69201 ( .A(n65494), .B(n65493), .Y(n65495) );
  NOR2X1 U69202 ( .A(n41593), .B(n41584), .Y(n65498) );
  NAND2X1 U69203 ( .A(n65497), .B(n65511), .Y(n65864) );
  NAND2X1 U69204 ( .A(n65498), .B(n65864), .Y(n66007) );
  NAND2X1 U69205 ( .A(n40472), .B(n44026), .Y(n65621) );
  INVX1 U69206 ( .A(n65621), .Y(n65499) );
  XNOR2X1 U69207 ( .A(n66007), .B(n65499), .Y(n65500) );
  XNOR2X1 U69208 ( .A(n65633), .B(n65500), .Y(n65501) );
  XNOR2X1 U69209 ( .A(n65502), .B(n65501), .Y(n65998) );
  INVX1 U69210 ( .A(n65998), .Y(n65987) );
  NAND2X1 U69211 ( .A(n43809), .B(n44056), .Y(n65874) );
  NAND2X1 U69212 ( .A(n43612), .B(n43820), .Y(n72558) );
  XNOR2X1 U69213 ( .A(n65874), .B(n43621), .Y(n65503) );
  XNOR2X1 U69214 ( .A(n41427), .B(n65503), .Y(n65534) );
  NOR2X1 U69215 ( .A(n65509), .B(n38929), .Y(n65521) );
  NOR2X1 U69216 ( .A(n65504), .B(n65509), .Y(n65508) );
  NAND2X1 U69217 ( .A(n65523), .B(n65522), .Y(n65505) );
  OR2X1 U69218 ( .A(n65506), .B(n65505), .Y(n65507) );
  NAND2X1 U69219 ( .A(n65508), .B(n65507), .Y(n65519) );
  INVX1 U69220 ( .A(n65509), .Y(n65517) );
  XNOR2X1 U69221 ( .A(n65620), .B(n65510), .Y(n65514) );
  XNOR2X1 U69222 ( .A(n65512), .B(n65511), .Y(n65513) );
  XNOR2X1 U69223 ( .A(n65514), .B(n65513), .Y(n65515) );
  XOR2X1 U69224 ( .A(n65619), .B(n65515), .Y(n65516) );
  NAND2X1 U69225 ( .A(n65517), .B(n65516), .Y(n65518) );
  NAND2X1 U69226 ( .A(n65519), .B(n65518), .Y(n65520) );
  NOR2X1 U69227 ( .A(n65521), .B(n65520), .Y(n65871) );
  NOR2X1 U69228 ( .A(n39967), .B(n40072), .Y(n65525) );
  NAND2X1 U69229 ( .A(n65525), .B(n65524), .Y(n65526) );
  NAND2X1 U69230 ( .A(n65527), .B(n65526), .Y(n65528) );
  NAND2X1 U69231 ( .A(n65528), .B(n38929), .Y(n65533) );
  INVX1 U69232 ( .A(n65620), .Y(n65625) );
  XNOR2X1 U69233 ( .A(n65531), .B(n65530), .Y(n65532) );
  NAND2X1 U69234 ( .A(n65533), .B(n65532), .Y(n65870) );
  NAND2X1 U69235 ( .A(n65871), .B(n65870), .Y(n66000) );
  INVX1 U69236 ( .A(n65875), .Y(n65608) );
  XNOR2X1 U69237 ( .A(n65534), .B(n65608), .Y(n65535) );
  XNOR2X1 U69238 ( .A(n39631), .B(n65535), .Y(n65885) );
  XNOR2X1 U69239 ( .A(n65885), .B(n43546), .Y(n65536) );
  XNOR2X1 U69240 ( .A(n36525), .B(n65536), .Y(n65911) );
  XNOR2X1 U69241 ( .A(n65537), .B(n65917), .Y(n65544) );
  XNOR2X1 U69242 ( .A(n65540), .B(n65539), .Y(n65542) );
  NAND2X1 U69243 ( .A(n43664), .B(n65542), .Y(n65541) );
  NOR2X1 U69244 ( .A(n41074), .B(n41346), .Y(n65543) );
  XNOR2X1 U69245 ( .A(n65543), .B(n65544), .Y(n65929) );
  INVX1 U69246 ( .A(n65929), .Y(n65545) );
  XNOR2X1 U69247 ( .A(n43655), .B(n43643), .Y(n71102) );
  INVX1 U69248 ( .A(n71102), .Y(n71744) );
  XNOR2X1 U69249 ( .A(n65545), .B(n71744), .Y(n65549) );
  NAND2X1 U69250 ( .A(n40142), .B(n65546), .Y(n65923) );
  NAND2X1 U69251 ( .A(n41105), .B(n65923), .Y(n65548) );
  NAND2X1 U69252 ( .A(n65547), .B(n43646), .Y(n65920) );
  XNOR2X1 U69253 ( .A(n65549), .B(n41109), .Y(n65550) );
  XNOR2X1 U69254 ( .A(n65551), .B(n65550), .Y(n65602) );
  XNOR2X1 U69255 ( .A(n65596), .B(n43679), .Y(n65563) );
  INVX1 U69256 ( .A(n65554), .Y(n65597) );
  NOR2X1 U69257 ( .A(n65597), .B(n64904), .Y(n65560) );
  NAND2X1 U69258 ( .A(n65595), .B(n65558), .Y(n65559) );
  NOR2X1 U69259 ( .A(n65560), .B(n65559), .Y(n65561) );
  NOR2X1 U69260 ( .A(n41191), .B(n65561), .Y(n65562) );
  XNOR2X1 U69261 ( .A(n65563), .B(n65562), .Y(n65594) );
  XNOR2X1 U69262 ( .A(n43512), .B(n65594), .Y(n65564) );
  XNOR2X1 U69263 ( .A(n65565), .B(n65564), .Y(n65585) );
  XNOR2X1 U69264 ( .A(n65585), .B(n43693), .Y(n65566) );
  XNOR2X1 U69265 ( .A(n37914), .B(n65566), .Y(n65583) );
  INVX1 U69266 ( .A(n65583), .Y(n65580) );
  XNOR2X1 U69267 ( .A(n43708), .B(n65580), .Y(n65574) );
  INVX1 U69268 ( .A(n65570), .Y(n65567) );
  NAND2X1 U69269 ( .A(n43705), .B(n65570), .Y(n65571) );
  INVX1 U69270 ( .A(n65581), .Y(n65573) );
  XNOR2X1 U69271 ( .A(n65574), .B(n65573), .Y(n65579) );
  XNOR2X1 U69272 ( .A(n65576), .B(n65575), .Y(n65577) );
  XNOR2X1 U69273 ( .A(n65577), .B(n41950), .Y(n65578) );
  MX2X1 U69274 ( .A(n65579), .B(n65578), .S0(n43719), .Y(u_muldiv_result_r[10]) );
  NAND2X1 U69275 ( .A(u_muldiv_mult_result_q[10]), .B(n44633), .Y(n14046) );
  NAND2X1 U69276 ( .A(n43705), .B(n65580), .Y(n65582) );
  NAND2X1 U69277 ( .A(n65582), .B(n65581), .Y(n66240) );
  NAND2X1 U69278 ( .A(n65583), .B(n43710), .Y(n66237) );
  NAND2X1 U69279 ( .A(n66237), .B(n66240), .Y(n65939) );
  NAND2X1 U69280 ( .A(n65585), .B(n43699), .Y(n65584) );
  NAND2X1 U69281 ( .A(n41470), .B(n65584), .Y(n65946) );
  NOR2X1 U69282 ( .A(n65594), .B(n43513), .Y(n65587) );
  NOR2X1 U69283 ( .A(n37404), .B(n65591), .Y(n65593) );
  NAND2X1 U69284 ( .A(n65594), .B(n43513), .Y(n65953) );
  NOR2X1 U69285 ( .A(n65597), .B(n41191), .Y(n65599) );
  NAND2X1 U69286 ( .A(n65599), .B(n65598), .Y(n65600) );
  NAND2X1 U69287 ( .A(n43522), .B(n65602), .Y(n65604) );
  NAND2X1 U69288 ( .A(n65604), .B(n65603), .Y(n65605) );
  XNOR2X1 U69289 ( .A(n65874), .B(n65988), .Y(n65607) );
  XNOR2X1 U69290 ( .A(n38193), .B(n65607), .Y(n65609) );
  XNOR2X1 U69291 ( .A(n65609), .B(n65608), .Y(n65610) );
  XNOR2X1 U69292 ( .A(n39631), .B(n65610), .Y(n65612) );
  INVX1 U69293 ( .A(n65612), .Y(n65611) );
  NAND2X1 U69294 ( .A(n65612), .B(n43628), .Y(n65614) );
  NAND2X1 U69295 ( .A(n65871), .B(n65870), .Y(n65875) );
  NAND2X1 U69296 ( .A(n38193), .B(n66000), .Y(n65994) );
  NAND2X1 U69297 ( .A(n39514), .B(n65627), .Y(n65616) );
  NOR2X1 U69298 ( .A(n65630), .B(n65616), .Y(n65618) );
  OR2X1 U69299 ( .A(n44022), .B(n65621), .Y(n65617) );
  NOR2X1 U69300 ( .A(n65620), .B(n65627), .Y(n65624) );
  NAND2X1 U69301 ( .A(n65626), .B(n65625), .Y(n65622) );
  NAND2X1 U69302 ( .A(n65622), .B(n65621), .Y(n65623) );
  NOR2X1 U69303 ( .A(n65624), .B(n65623), .Y(n65632) );
  NOR2X1 U69304 ( .A(n65626), .B(n65625), .Y(n65628) );
  NAND2X1 U69305 ( .A(n65628), .B(n65627), .Y(n65629) );
  NAND2X1 U69306 ( .A(n65630), .B(n65629), .Y(n65631) );
  NAND2X1 U69307 ( .A(n65632), .B(n65631), .Y(n65635) );
  XNOR2X1 U69308 ( .A(n66007), .B(n65633), .Y(n65634) );
  NAND2X1 U69309 ( .A(n65635), .B(n65634), .Y(n65991) );
  NAND2X1 U69310 ( .A(n40470), .B(n44049), .Y(n67180) );
  INVX1 U69311 ( .A(n67180), .Y(n66294) );
  XNOR2X1 U69312 ( .A(n42057), .B(n66294), .Y(n65868) );
  INVX1 U69313 ( .A(n66016), .Y(n65858) );
  NOR2X1 U69314 ( .A(n39029), .B(n41257), .Y(n65636) );
  NAND2X1 U69315 ( .A(n65636), .B(n66475), .Y(n66009) );
  NOR2X1 U69316 ( .A(n65640), .B(n41283), .Y(n65642) );
  NAND2X1 U69317 ( .A(n65642), .B(n65641), .Y(n65644) );
  NAND2X1 U69318 ( .A(n42632), .B(n44000), .Y(n66022) );
  NAND2X1 U69319 ( .A(n43725), .B(n44008), .Y(n66028) );
  XNOR2X1 U69320 ( .A(n66022), .B(n66028), .Y(n65854) );
  NOR2X1 U69321 ( .A(n43987), .B(n65655), .Y(n65646) );
  NOR2X1 U69322 ( .A(n65646), .B(n65657), .Y(n65649) );
  NAND2X1 U69323 ( .A(n43989), .B(n65655), .Y(n65647) );
  NAND2X1 U69324 ( .A(n37320), .B(n65647), .Y(n65648) );
  NOR2X1 U69325 ( .A(n65649), .B(n65648), .Y(n65654) );
  XNOR2X1 U69326 ( .A(n41185), .B(n65664), .Y(n65650) );
  XNOR2X1 U69327 ( .A(n65650), .B(n41376), .Y(n65651) );
  XNOR2X1 U69328 ( .A(n65652), .B(n65651), .Y(n65661) );
  NAND2X1 U69329 ( .A(n65658), .B(n65657), .Y(n65660) );
  NAND2X1 U69330 ( .A(n65660), .B(n65659), .Y(n65662) );
  NOR2X1 U69331 ( .A(n65665), .B(n36774), .Y(n65670) );
  INVX1 U69332 ( .A(n65666), .Y(n65668) );
  NOR2X1 U69333 ( .A(n65668), .B(n65667), .Y(n65669) );
  NOR2X1 U69334 ( .A(n65670), .B(n65669), .Y(n65674) );
  NAND2X1 U69335 ( .A(n65672), .B(n65671), .Y(n65673) );
  NAND2X1 U69336 ( .A(n43772), .B(n43992), .Y(n66201) );
  NAND2X1 U69337 ( .A(n43798), .B(n43983), .Y(n66178) );
  NAND2X1 U69338 ( .A(n43942), .B(n42711), .Y(n66162) );
  XNOR2X1 U69339 ( .A(n65676), .B(n39113), .Y(n65677) );
  XNOR2X1 U69340 ( .A(n39117), .B(n65677), .Y(n65681) );
  INVX1 U69341 ( .A(n65681), .Y(n65678) );
  NAND2X1 U69342 ( .A(n65679), .B(n65678), .Y(n65684) );
  NAND2X1 U69343 ( .A(n65681), .B(n65680), .Y(n65682) );
  NAND2X1 U69344 ( .A(n65682), .B(n65813), .Y(n65683) );
  NAND2X1 U69345 ( .A(n65684), .B(n65683), .Y(n66450) );
  INVX1 U69346 ( .A(n66450), .Y(n66039) );
  XNOR2X1 U69347 ( .A(n36657), .B(n65704), .Y(n65685) );
  XNOR2X1 U69348 ( .A(n65685), .B(n41171), .Y(n65686) );
  XNOR2X1 U69349 ( .A(n39113), .B(n65686), .Y(n65689) );
  INVX1 U69350 ( .A(n65689), .Y(n66049) );
  NAND2X1 U69351 ( .A(n66049), .B(n66048), .Y(n65688) );
  NAND2X1 U69352 ( .A(n65688), .B(n65687), .Y(n65691) );
  NAND2X1 U69353 ( .A(n65690), .B(n65689), .Y(n66064) );
  NAND2X1 U69354 ( .A(n65691), .B(n66064), .Y(n66036) );
  NAND2X1 U69355 ( .A(n43795), .B(n43934), .Y(n66448) );
  NAND2X1 U69356 ( .A(n65698), .B(n38914), .Y(n65692) );
  NOR2X1 U69357 ( .A(n65693), .B(n65692), .Y(n65703) );
  NOR2X1 U69358 ( .A(n65695), .B(n65694), .Y(n65697) );
  NAND2X1 U69359 ( .A(n65704), .B(n65699), .Y(n65700) );
  NOR2X1 U69360 ( .A(n65701), .B(n65700), .Y(n65702) );
  NOR2X1 U69361 ( .A(n65703), .B(n65702), .Y(n65706) );
  NAND2X1 U69362 ( .A(n65704), .B(n40984), .Y(n65705) );
  NAND2X1 U69363 ( .A(n65708), .B(n65707), .Y(n65709) );
  NAND2X1 U69364 ( .A(n65709), .B(n38914), .Y(n65711) );
  NAND2X1 U69365 ( .A(n65711), .B(n65710), .Y(n65712) );
  NAND2X1 U69366 ( .A(n40984), .B(n65712), .Y(n66078) );
  NAND2X1 U69367 ( .A(n41122), .B(n66078), .Y(n66081) );
  NAND2X1 U69368 ( .A(n65719), .B(n38622), .Y(n66055) );
  INVX1 U69369 ( .A(n65715), .Y(n65718) );
  INVX1 U69370 ( .A(n65719), .Y(n66088) );
  NAND2X1 U69371 ( .A(n43909), .B(n38313), .Y(n66087) );
  NAND2X1 U69372 ( .A(n36773), .B(n65723), .Y(n66085) );
  NAND2X1 U69373 ( .A(n65726), .B(n65725), .Y(n65727) );
  NAND2X1 U69374 ( .A(n66085), .B(n66084), .Y(n66097) );
  INVX1 U69375 ( .A(n66097), .Y(n66094) );
  XNOR2X1 U69376 ( .A(n66087), .B(n66094), .Y(n65807) );
  NOR2X1 U69377 ( .A(n65736), .B(n65739), .Y(n65731) );
  INVX1 U69378 ( .A(n65728), .Y(n65735) );
  NAND2X1 U69379 ( .A(n65735), .B(n65729), .Y(n65730) );
  NOR2X1 U69380 ( .A(n65731), .B(n65730), .Y(n65734) );
  NAND2X1 U69381 ( .A(n65735), .B(n65736), .Y(n65732) );
  NOR2X1 U69382 ( .A(n40478), .B(n65732), .Y(n65733) );
  NOR2X1 U69383 ( .A(n65734), .B(n65733), .Y(n65746) );
  NOR2X1 U69384 ( .A(n65735), .B(n41000), .Y(n65742) );
  INVX1 U69385 ( .A(n65736), .Y(n65738) );
  NAND2X1 U69386 ( .A(n65738), .B(n65737), .Y(n65740) );
  NAND2X1 U69387 ( .A(n65740), .B(n65739), .Y(n65741) );
  NAND2X1 U69388 ( .A(n65742), .B(n65741), .Y(n65744) );
  XNOR2X1 U69389 ( .A(n40999), .B(n41224), .Y(n65743) );
  NAND2X1 U69390 ( .A(n65744), .B(n65743), .Y(n65745) );
  NAND2X1 U69391 ( .A(n65746), .B(n65745), .Y(n66103) );
  NAND2X1 U69392 ( .A(n43903), .B(n43487), .Y(n67057) );
  INVX1 U69393 ( .A(n65767), .Y(n65752) );
  NOR2X1 U69394 ( .A(n65769), .B(n65752), .Y(n65750) );
  NOR2X1 U69395 ( .A(n65750), .B(n65749), .Y(n65751) );
  NAND2X1 U69396 ( .A(n65751), .B(n39129), .Y(n66144) );
  NAND2X1 U69397 ( .A(n65752), .B(n43501), .Y(n65753) );
  NOR2X1 U69398 ( .A(n43957), .B(n65753), .Y(n65759) );
  INVX1 U69399 ( .A(n65762), .Y(n65755) );
  NOR2X1 U69400 ( .A(n65755), .B(n65754), .Y(n65757) );
  NAND2X1 U69401 ( .A(n65757), .B(n65756), .Y(n65758) );
  NAND2X1 U69402 ( .A(n65759), .B(n65758), .Y(n66149) );
  NAND2X1 U69403 ( .A(n66144), .B(n66149), .Y(n65771) );
  NOR2X1 U69404 ( .A(n65761), .B(n65760), .Y(n65765) );
  NAND2X1 U69405 ( .A(n40313), .B(n65763), .Y(n65764) );
  NAND2X1 U69406 ( .A(n65765), .B(n65764), .Y(n66148) );
  NAND2X1 U69407 ( .A(n65767), .B(n65766), .Y(n65768) );
  NAND2X1 U69408 ( .A(n65769), .B(n65768), .Y(n66147) );
  NAND2X1 U69409 ( .A(n66148), .B(n66147), .Y(n65770) );
  OR2X1 U69410 ( .A(n65771), .B(n65770), .Y(n66403) );
  NAND2X1 U69411 ( .A(n43952), .B(n39653), .Y(n66123) );
  NAND2X1 U69412 ( .A(n41498), .B(n43605), .Y(n72364) );
  INVX1 U69413 ( .A(n72364), .Y(n71845) );
  OR2X1 U69414 ( .A(n66131), .B(n65772), .Y(n65775) );
  NAND2X1 U69415 ( .A(n65774), .B(n65773), .Y(n66125) );
  NOR2X1 U69416 ( .A(n65775), .B(n66125), .Y(n72367) );
  XNOR2X1 U69417 ( .A(n71845), .B(n72367), .Y(n66725) );
  INVX1 U69418 ( .A(n66725), .Y(n71847) );
  NAND2X1 U69419 ( .A(n65776), .B(n65780), .Y(n65777) );
  NAND2X1 U69420 ( .A(n41498), .B(n65777), .Y(n66139) );
  NAND2X1 U69421 ( .A(n43869), .B(n43517), .Y(n66385) );
  INVX1 U69422 ( .A(n66385), .Y(n66120) );
  XNOR2X1 U69423 ( .A(n66384), .B(n66120), .Y(n65788) );
  INVX1 U69424 ( .A(n65778), .Y(n65779) );
  NAND2X1 U69425 ( .A(n65779), .B(n41505), .Y(n65785) );
  INVX1 U69426 ( .A(n65787), .Y(n65782) );
  NAND2X1 U69427 ( .A(n65782), .B(n65781), .Y(n65783) );
  NAND2X1 U69428 ( .A(n41505), .B(n65783), .Y(n65784) );
  NAND2X1 U69429 ( .A(n65785), .B(n65784), .Y(n66116) );
  INVX1 U69430 ( .A(n66116), .Y(n66389) );
  NAND2X1 U69431 ( .A(n65787), .B(n65786), .Y(n66117) );
  NAND2X1 U69432 ( .A(n66389), .B(n66117), .Y(n66115) );
  NAND2X1 U69433 ( .A(n43879), .B(n43501), .Y(n66399) );
  INVX1 U69434 ( .A(n66399), .Y(n66100) );
  NAND2X1 U69435 ( .A(n43889), .B(n43497), .Y(n66355) );
  INVX1 U69436 ( .A(n66355), .Y(n66111) );
  XNOR2X1 U69437 ( .A(n66100), .B(n66111), .Y(n65789) );
  NAND2X1 U69438 ( .A(n43492), .B(n43899), .Y(n66411) );
  INVX1 U69439 ( .A(n66411), .Y(n66106) );
  XNOR2X1 U69440 ( .A(n65789), .B(n66106), .Y(n65790) );
  XNOR2X1 U69441 ( .A(n66400), .B(n65790), .Y(n65791) );
  XNOR2X1 U69442 ( .A(n66403), .B(n65791), .Y(n65805) );
  NOR2X1 U69443 ( .A(n65792), .B(n65796), .Y(n65794) );
  NAND2X1 U69444 ( .A(n40998), .B(n65802), .Y(n65793) );
  NAND2X1 U69445 ( .A(n65794), .B(n65793), .Y(n65800) );
  INVX1 U69446 ( .A(n65795), .Y(n65798) );
  NAND2X1 U69447 ( .A(n65801), .B(n65796), .Y(n65797) );
  NAND2X1 U69448 ( .A(n65798), .B(n65797), .Y(n65799) );
  AND2X1 U69449 ( .A(n65800), .B(n65799), .Y(n66113) );
  NOR2X1 U69450 ( .A(n43874), .B(n65801), .Y(n65803) );
  INVX1 U69451 ( .A(n66108), .Y(n66112) );
  XNOR2X1 U69452 ( .A(n65805), .B(n41220), .Y(n66093) );
  XNOR2X1 U69453 ( .A(n67057), .B(n66093), .Y(n65806) );
  XOR2X1 U69454 ( .A(n66103), .B(n65806), .Y(n66086) );
  XNOR2X1 U69455 ( .A(n65807), .B(n66086), .Y(n66077) );
  NAND2X1 U69456 ( .A(n43928), .B(n43775), .Y(n66047) );
  NAND2X1 U69457 ( .A(n43918), .B(n43478), .Y(n66321) );
  INVX1 U69458 ( .A(n66321), .Y(n66079) );
  XNOR2X1 U69459 ( .A(n66047), .B(n66079), .Y(n65808) );
  XNOR2X1 U69460 ( .A(n66077), .B(n65808), .Y(n65809) );
  XNOR2X1 U69461 ( .A(n40309), .B(n65809), .Y(n65810) );
  XNOR2X1 U69462 ( .A(n38097), .B(n65810), .Y(n66035) );
  XNOR2X1 U69463 ( .A(n66448), .B(n66035), .Y(n65811) );
  INVX1 U69464 ( .A(n65815), .Y(n65819) );
  INVX1 U69465 ( .A(n65812), .Y(n65820) );
  XNOR2X1 U69466 ( .A(n65820), .B(n39891), .Y(n65814) );
  NAND2X1 U69467 ( .A(n65819), .B(n65814), .Y(n66164) );
  NAND2X1 U69468 ( .A(n65829), .B(n65828), .Y(n65816) );
  NAND2X1 U69469 ( .A(n65834), .B(n65816), .Y(n65817) );
  NAND2X1 U69470 ( .A(n66168), .B(n65817), .Y(n65818) );
  NAND2X1 U69471 ( .A(n66164), .B(n65818), .Y(n66163) );
  NAND2X1 U69472 ( .A(n42659), .B(n43973), .Y(n66174) );
  INVX1 U69473 ( .A(n65831), .Y(n65835) );
  XNOR2X1 U69474 ( .A(n65820), .B(n65819), .Y(n65821) );
  XNOR2X1 U69475 ( .A(n65821), .B(n39891), .Y(n65822) );
  XNOR2X1 U69476 ( .A(n39451), .B(n65822), .Y(n65824) );
  INVX1 U69477 ( .A(n65824), .Y(n65823) );
  NAND2X1 U69478 ( .A(n65824), .B(n65831), .Y(n65826) );
  XOR2X1 U69479 ( .A(n66174), .B(n66176), .Y(n65827) );
  XNOR2X1 U69480 ( .A(n66178), .B(n66197), .Y(n65852) );
  NOR2X1 U69481 ( .A(n65831), .B(n65834), .Y(n65833) );
  NAND2X1 U69482 ( .A(n65829), .B(n65828), .Y(n65830) );
  NOR2X1 U69483 ( .A(n65831), .B(n65830), .Y(n65832) );
  NOR2X1 U69484 ( .A(n65833), .B(n65832), .Y(n65839) );
  INVX1 U69485 ( .A(n65834), .Y(n65836) );
  NOR2X1 U69486 ( .A(n65836), .B(n65835), .Y(n65837) );
  NAND2X1 U69487 ( .A(n65837), .B(n65830), .Y(n65838) );
  NAND2X1 U69488 ( .A(n65839), .B(n65838), .Y(n65841) );
  XNOR2X1 U69489 ( .A(n65841), .B(n65840), .Y(n65842) );
  XNOR2X1 U69490 ( .A(n39281), .B(n65842), .Y(n66189) );
  INVX1 U69491 ( .A(n66189), .Y(n66192) );
  NAND2X1 U69492 ( .A(n66189), .B(n65844), .Y(n65851) );
  INVX1 U69493 ( .A(n65845), .Y(n65846) );
  NOR2X1 U69494 ( .A(n65846), .B(n66179), .Y(n65847) );
  NOR2X1 U69495 ( .A(n65847), .B(n66180), .Y(n65848) );
  NAND2X1 U69496 ( .A(n65849), .B(n66187), .Y(n65850) );
  INVX1 U69497 ( .A(n66023), .Y(n66206) );
  XNOR2X1 U69498 ( .A(n66205), .B(n66206), .Y(n65853) );
  XNOR2X1 U69499 ( .A(n65854), .B(n65853), .Y(n65855) );
  XOR2X1 U69500 ( .A(n66031), .B(n65855), .Y(n66474) );
  NAND2X1 U69501 ( .A(n40484), .B(n44026), .Y(n66861) );
  NAND2X1 U69502 ( .A(n43787), .B(n44017), .Y(n66014) );
  INVX1 U69503 ( .A(n66014), .Y(n66021) );
  XNOR2X1 U69504 ( .A(n66861), .B(n66021), .Y(n65856) );
  XNOR2X1 U69505 ( .A(n66474), .B(n65856), .Y(n65857) );
  XNOR2X1 U69506 ( .A(n66009), .B(n65857), .Y(n65867) );
  XNOR2X1 U69507 ( .A(n65858), .B(n41362), .Y(n65859) );
  XNOR2X1 U69508 ( .A(n65859), .B(n40199), .Y(n65860) );
  NOR2X1 U69509 ( .A(n41593), .B(n41584), .Y(n65862) );
  NAND2X1 U69510 ( .A(n65862), .B(n65864), .Y(n65863) );
  NOR2X1 U69511 ( .A(n41302), .B(n40225), .Y(n65866) );
  NAND2X1 U69512 ( .A(n65498), .B(n65864), .Y(n66858) );
  NAND2X1 U69513 ( .A(n66008), .B(n66858), .Y(n65865) );
  NAND2X1 U69514 ( .A(n65866), .B(n65865), .Y(n66011) );
  XNOR2X1 U69515 ( .A(n65867), .B(n40077), .Y(n66293) );
  XNOR2X1 U69516 ( .A(n65868), .B(n39414), .Y(n65869) );
  XNOR2X1 U69517 ( .A(n38888), .B(n65869), .Y(n65978) );
  INVX1 U69518 ( .A(n65978), .Y(n65872) );
  NAND2X1 U69519 ( .A(n65988), .B(n38783), .Y(n65974) );
  XNOR2X1 U69520 ( .A(n43621), .B(n43564), .Y(n67993) );
  INVX1 U69521 ( .A(n67993), .Y(n71794) );
  XNOR2X1 U69522 ( .A(n39740), .B(n71794), .Y(n65883) );
  INVX1 U69523 ( .A(n65874), .Y(n65986) );
  NAND2X1 U69524 ( .A(n65876), .B(n44049), .Y(n65877) );
  NAND2X1 U69525 ( .A(n65878), .B(n65877), .Y(n65879) );
  OR2X1 U69526 ( .A(n65881), .B(n65879), .Y(n65984) );
  NAND2X1 U69527 ( .A(n65986), .B(n65984), .Y(n65882) );
  NAND2X1 U69528 ( .A(n65881), .B(n65880), .Y(n65981) );
  XNOR2X1 U69529 ( .A(n65883), .B(n41322), .Y(n65884) );
  INVX1 U69530 ( .A(n66224), .Y(n66222) );
  NAND2X1 U69531 ( .A(n66517), .B(n43547), .Y(n65888) );
  INVX1 U69532 ( .A(n66517), .Y(n65886) );
  NAND2X1 U69533 ( .A(n43545), .B(n65886), .Y(n65894) );
  NAND2X1 U69534 ( .A(n65888), .B(n65894), .Y(n65887) );
  NOR2X1 U69535 ( .A(n66222), .B(n65887), .Y(n65893) );
  NOR2X1 U69536 ( .A(n66222), .B(n43553), .Y(n65890) );
  NOR2X1 U69537 ( .A(n66224), .B(n65888), .Y(n65889) );
  NOR2X1 U69538 ( .A(n65890), .B(n65889), .Y(n65891) );
  NOR2X1 U69539 ( .A(n39895), .B(n65891), .Y(n65892) );
  NOR2X1 U69540 ( .A(n65893), .B(n65892), .Y(n65898) );
  OR2X1 U69541 ( .A(n66224), .B(n65894), .Y(n65896) );
  NAND2X1 U69542 ( .A(n66224), .B(n43551), .Y(n65895) );
  NAND2X1 U69543 ( .A(n65896), .B(n65895), .Y(n65897) );
  NAND2X1 U69544 ( .A(n39895), .B(n65897), .Y(n65973) );
  NAND2X1 U69545 ( .A(n65898), .B(n65973), .Y(n65972) );
  INVX1 U69546 ( .A(n65900), .Y(n65908) );
  NOR2X1 U69547 ( .A(n39266), .B(n65901), .Y(n65902) );
  NOR2X1 U69548 ( .A(n38172), .B(n65902), .Y(n65906) );
  NAND2X1 U69549 ( .A(n65904), .B(n65903), .Y(n65905) );
  NAND2X1 U69550 ( .A(n65906), .B(n65905), .Y(n65907) );
  NOR2X1 U69551 ( .A(n65908), .B(n65907), .Y(n65909) );
  NOR2X1 U69552 ( .A(n39081), .B(n65909), .Y(n65914) );
  INVX1 U69553 ( .A(n65915), .Y(n65912) );
  NAND2X1 U69554 ( .A(n65912), .B(n43638), .Y(n65913) );
  XNOR2X1 U69555 ( .A(n43639), .B(n66275), .Y(n65916) );
  XOR2X1 U69556 ( .A(n65972), .B(n65916), .Y(n65969) );
  XNOR2X1 U69557 ( .A(n41078), .B(n65917), .Y(n65918) );
  NAND2X1 U69558 ( .A(n40142), .B(n65929), .Y(n65928) );
  NOR2X1 U69559 ( .A(n43642), .B(n65929), .Y(n65922) );
  INVX1 U69560 ( .A(n65920), .Y(n65921) );
  INVX1 U69561 ( .A(n65923), .Y(n65927) );
  NAND2X1 U69562 ( .A(n65925), .B(n65924), .Y(n65926) );
  NAND2X1 U69563 ( .A(n65928), .B(n66531), .Y(n66534) );
  INVX1 U69564 ( .A(n65965), .Y(n65967) );
  XNOR2X1 U69565 ( .A(n43655), .B(n65967), .Y(n65960) );
  XNOR2X1 U69566 ( .A(n65929), .B(n43643), .Y(n65930) );
  XNOR2X1 U69567 ( .A(n41109), .B(n65930), .Y(n65932) );
  INVX1 U69568 ( .A(n65932), .Y(n65933) );
  XNOR2X1 U69569 ( .A(n43530), .B(n65966), .Y(n65934) );
  XOR2X1 U69570 ( .A(n65960), .B(n65934), .Y(n65950) );
  XNOR2X1 U69571 ( .A(n40137), .B(n65950), .Y(n66233) );
  XNOR2X1 U69572 ( .A(n43509), .B(n43679), .Y(n72583) );
  XNOR2X1 U69573 ( .A(n66233), .B(n72583), .Y(n65935) );
  XNOR2X1 U69574 ( .A(n43698), .B(n65947), .Y(n65936) );
  XNOR2X1 U69575 ( .A(n65937), .B(n65936), .Y(n66242) );
  XNOR2X1 U69576 ( .A(n43714), .B(n37911), .Y(n65938) );
  XNOR2X1 U69577 ( .A(n65939), .B(n65938), .Y(n65944) );
  XNOR2X1 U69578 ( .A(n65941), .B(n65940), .Y(n65942) );
  XOR2X1 U69579 ( .A(n41959), .B(n65942), .Y(n65943) );
  MX2X1 U69580 ( .A(n65944), .B(n65943), .S0(n43719), .Y(u_muldiv_result_r[11]) );
  NAND2X1 U69581 ( .A(u_muldiv_mult_result_q[11]), .B(n44633), .Y(n14035) );
  NOR2X1 U69582 ( .A(n65947), .B(n43702), .Y(n65945) );
  NAND2X1 U69583 ( .A(n37932), .B(n39067), .Y(n65949) );
  NAND2X1 U69584 ( .A(n65947), .B(n43700), .Y(n65948) );
  NAND2X1 U69585 ( .A(n65949), .B(n65948), .Y(n66546) );
  XNOR2X1 U69586 ( .A(n38047), .B(n40137), .Y(n65951) );
  XNOR2X1 U69587 ( .A(n65951), .B(n65950), .Y(n65952) );
  NAND2X1 U69588 ( .A(n43505), .B(n41218), .Y(n65959) );
  INVX1 U69589 ( .A(n65953), .Y(n65955) );
  NOR2X1 U69590 ( .A(n43507), .B(n41218), .Y(n65954) );
  NOR2X1 U69591 ( .A(n65955), .B(n65954), .Y(n65957) );
  NAND2X1 U69592 ( .A(n65957), .B(n65956), .Y(n65958) );
  NAND2X1 U69593 ( .A(n65959), .B(n65958), .Y(n66252) );
  NAND2X1 U69594 ( .A(n43522), .B(n65963), .Y(n65962) );
  NAND2X1 U69595 ( .A(n65961), .B(n65962), .Y(n66895) );
  INVX1 U69596 ( .A(n65963), .Y(n65964) );
  NAND2X1 U69597 ( .A(n65964), .B(n43531), .Y(n66899) );
  NAND2X1 U69598 ( .A(n65965), .B(n43660), .Y(n66261) );
  NAND2X1 U69599 ( .A(n65966), .B(n66261), .Y(n65968) );
  XNOR2X1 U69600 ( .A(n43524), .B(n41107), .Y(n66230) );
  NAND2X1 U69601 ( .A(n43664), .B(n65969), .Y(n66267) );
  NAND2X1 U69602 ( .A(n65973), .B(n43671), .Y(n65971) );
  NAND2X1 U69603 ( .A(n65971), .B(n65970), .Y(n66266) );
  NAND2X1 U69604 ( .A(n66266), .B(n66267), .Y(n66530) );
  NAND2X1 U69605 ( .A(n43632), .B(n65972), .Y(n66272) );
  NAND2X1 U69606 ( .A(n65973), .B(n43638), .Y(n66274) );
  NAND2X1 U69607 ( .A(n66274), .B(n66275), .Y(n66598) );
  XNOR2X1 U69608 ( .A(n43666), .B(n43633), .Y(n69861) );
  NOR2X1 U69609 ( .A(n39740), .B(n43560), .Y(n65983) );
  NAND2X1 U69610 ( .A(n39708), .B(n65974), .Y(n65976) );
  NOR2X1 U69611 ( .A(n65978), .B(n65977), .Y(n65979) );
  NAND2X1 U69612 ( .A(n38783), .B(n65979), .Y(n65980) );
  NOR2X1 U69613 ( .A(n65985), .B(n65981), .Y(n65982) );
  NOR2X1 U69614 ( .A(n38193), .B(n66000), .Y(n65990) );
  NAND2X1 U69615 ( .A(n65988), .B(n42057), .Y(n65989) );
  NOR2X1 U69616 ( .A(n65990), .B(n65989), .Y(n65997) );
  NAND2X1 U69617 ( .A(n65992), .B(n65991), .Y(n66005) );
  XNOR2X1 U69618 ( .A(n66005), .B(n66294), .Y(n65993) );
  XNOR2X1 U69619 ( .A(n39414), .B(n65993), .Y(n66001) );
  NOR2X1 U69620 ( .A(n42057), .B(n66001), .Y(n65995) );
  NOR2X1 U69621 ( .A(n39931), .B(n65995), .Y(n65996) );
  NAND2X1 U69622 ( .A(n44059), .B(n65998), .Y(n65999) );
  NOR2X1 U69623 ( .A(n44054), .B(n44050), .Y(n66002) );
  NOR2X1 U69624 ( .A(n40460), .B(n66002), .Y(n66003) );
  INVX1 U69625 ( .A(n66286), .Y(n66281) );
  NAND2X1 U69626 ( .A(n43613), .B(n40466), .Y(n72145) );
  NAND2X1 U69627 ( .A(n38476), .B(n66293), .Y(n66006) );
  NAND2X1 U69628 ( .A(n66294), .B(n66006), .Y(n66291) );
  NAND2X1 U69629 ( .A(n66626), .B(n66291), .Y(n66631) );
  INVX1 U69630 ( .A(n66631), .Y(n66278) );
  INVX1 U69631 ( .A(n66861), .Y(n66874) );
  INVX1 U69632 ( .A(n66474), .Y(n66478) );
  XNOR2X1 U69633 ( .A(n66009), .B(n66021), .Y(n66010) );
  XNOR2X1 U69634 ( .A(n66478), .B(n66010), .Y(n66865) );
  NAND2X1 U69635 ( .A(n39171), .B(n66011), .Y(n66492) );
  NOR2X1 U69636 ( .A(n41324), .B(n39948), .Y(n66013) );
  NAND2X1 U69637 ( .A(n66874), .B(n39171), .Y(n66012) );
  NAND2X1 U69638 ( .A(n66013), .B(n66012), .Y(n66880) );
  INVX1 U69639 ( .A(n66015), .Y(n66017) );
  NAND2X1 U69640 ( .A(n66017), .B(n66016), .Y(n66019) );
  NAND2X1 U69641 ( .A(n66021), .B(n66478), .Y(n66484) );
  NAND2X1 U69642 ( .A(n66485), .B(n66484), .Y(n66967) );
  INVX1 U69643 ( .A(n66022), .Y(n66207) );
  NOR2X1 U69644 ( .A(n40199), .B(n66024), .Y(n66027) );
  NAND2X1 U69645 ( .A(n66032), .B(n66031), .Y(n66033) );
  NAND2X1 U69646 ( .A(n40260), .B(n44000), .Y(n66659) );
  NAND2X1 U69647 ( .A(n43799), .B(n43992), .Y(n66839) );
  NAND2X1 U69648 ( .A(n42660), .B(n43983), .Y(n66819) );
  INVX1 U69649 ( .A(n66448), .Y(n66037) );
  NAND2X1 U69650 ( .A(n66037), .B(n66447), .Y(n66452) );
  NOR2X1 U69651 ( .A(n66037), .B(n66447), .Y(n66038) );
  OR2X1 U69652 ( .A(n66039), .B(n66038), .Y(n66040) );
  NAND2X1 U69653 ( .A(n66452), .B(n66040), .Y(n66161) );
  NOR2X1 U69654 ( .A(n66064), .B(n66047), .Y(n66051) );
  NOR2X1 U69655 ( .A(n36677), .B(n66041), .Y(n66042) );
  NOR2X1 U69656 ( .A(n37401), .B(n66042), .Y(n66046) );
  NAND2X1 U69657 ( .A(n66044), .B(n66043), .Y(n66045) );
  NAND2X1 U69658 ( .A(n66046), .B(n66045), .Y(n66069) );
  INVX1 U69659 ( .A(n66047), .Y(n66066) );
  NAND2X1 U69660 ( .A(n66049), .B(n66048), .Y(n66070) );
  NOR2X1 U69661 ( .A(n66051), .B(n66050), .Y(n66076) );
  INVX1 U69662 ( .A(n66057), .Y(n66052) );
  NOR2X1 U69663 ( .A(n66056), .B(n66052), .Y(n66054) );
  NAND2X1 U69664 ( .A(n66055), .B(n66321), .Y(n66053) );
  NOR2X1 U69665 ( .A(n66054), .B(n66053), .Y(n66062) );
  OR2X1 U69666 ( .A(n66321), .B(n66055), .Y(n66060) );
  NOR2X1 U69667 ( .A(n66056), .B(n66321), .Y(n66058) );
  NAND2X1 U69668 ( .A(n66058), .B(n66057), .Y(n66059) );
  NAND2X1 U69669 ( .A(n66060), .B(n66059), .Y(n66061) );
  NOR2X1 U69670 ( .A(n66062), .B(n66061), .Y(n66063) );
  XOR2X1 U69671 ( .A(n66077), .B(n66063), .Y(n66068) );
  INVX1 U69672 ( .A(n66064), .Y(n66065) );
  NOR2X1 U69673 ( .A(n66066), .B(n66065), .Y(n66067) );
  NOR2X1 U69674 ( .A(n66072), .B(n66067), .Y(n66074) );
  XNOR2X1 U69675 ( .A(n66068), .B(n38097), .Y(n66072) );
  NAND2X1 U69676 ( .A(n66070), .B(n66069), .Y(n66071) );
  NOR2X1 U69677 ( .A(n66072), .B(n66071), .Y(n66073) );
  NOR2X1 U69678 ( .A(n66074), .B(n66073), .Y(n66075) );
  NAND2X1 U69679 ( .A(n66076), .B(n66075), .Y(n66443) );
  NOR2X1 U69680 ( .A(n38922), .B(n66321), .Y(n66080) );
  NOR2X1 U69681 ( .A(n66080), .B(n39923), .Y(n66083) );
  NAND2X1 U69682 ( .A(n40336), .B(n66081), .Y(n66082) );
  INVX1 U69683 ( .A(n66084), .Y(n66345) );
  INVX1 U69684 ( .A(n66085), .Y(n66344) );
  NAND2X1 U69685 ( .A(n66089), .B(n40309), .Y(n66333) );
  NOR2X1 U69686 ( .A(n66090), .B(n66089), .Y(n66092) );
  NAND2X1 U69687 ( .A(n66333), .B(n66334), .Y(n66682) );
  INVX1 U69688 ( .A(n66103), .Y(n66417) );
  INVX1 U69689 ( .A(n66098), .Y(n66346) );
  NOR2X1 U69690 ( .A(n66346), .B(n67057), .Y(n66096) );
  NOR2X1 U69691 ( .A(n66094), .B(n67057), .Y(n66095) );
  NOR2X1 U69692 ( .A(n66096), .B(n66095), .Y(n66099) );
  NAND2X1 U69693 ( .A(n43918), .B(n38312), .Y(n66684) );
  INVX1 U69694 ( .A(n66684), .Y(n66337) );
  NAND2X1 U69695 ( .A(n43909), .B(n43486), .Y(n66340) );
  INVX1 U69696 ( .A(n66340), .Y(n66342) );
  XNOR2X1 U69697 ( .A(n66337), .B(n66342), .Y(n66155) );
  XNOR2X1 U69698 ( .A(n66400), .B(n66100), .Y(n66101) );
  XNOR2X1 U69699 ( .A(n66357), .B(n66111), .Y(n66102) );
  XNOR2X1 U69700 ( .A(n41220), .B(n66102), .Y(n66416) );
  NAND2X1 U69701 ( .A(n66416), .B(n66411), .Y(n66104) );
  NAND2X1 U69702 ( .A(n66104), .B(n66103), .Y(n66107) );
  INVX1 U69703 ( .A(n66416), .Y(n66105) );
  NAND2X1 U69704 ( .A(n66106), .B(n66105), .Y(n66415) );
  NAND2X1 U69705 ( .A(n66107), .B(n66415), .Y(n66423) );
  NOR2X1 U69706 ( .A(n66357), .B(n66108), .Y(n66109) );
  NAND2X1 U69707 ( .A(n66109), .B(n38224), .Y(n66110) );
  NAND2X1 U69708 ( .A(n66111), .B(n66110), .Y(n66114) );
  NAND2X1 U69709 ( .A(n66113), .B(n66112), .Y(n66356) );
  NAND2X1 U69710 ( .A(n66357), .B(n66356), .Y(n66360) );
  NAND2X1 U69711 ( .A(n66114), .B(n66360), .Y(n66703) );
  NAND2X1 U69712 ( .A(n66384), .B(n66115), .Y(n66122) );
  NOR2X1 U69713 ( .A(n66384), .B(n66116), .Y(n66118) );
  NAND2X1 U69714 ( .A(n66118), .B(n66117), .Y(n66119) );
  NAND2X1 U69715 ( .A(n66120), .B(n66119), .Y(n66121) );
  NAND2X1 U69716 ( .A(n66122), .B(n66121), .Y(n66745) );
  NAND2X1 U69717 ( .A(n43889), .B(n43501), .Y(n66398) );
  NAND2X1 U69718 ( .A(n43869), .B(n43608), .Y(n66366) );
  INVX1 U69719 ( .A(n66123), .Y(n66141) );
  NAND2X1 U69720 ( .A(n66141), .B(n43605), .Y(n72365) );
  INVX1 U69721 ( .A(n72365), .Y(n71844) );
  NAND2X1 U69722 ( .A(n71844), .B(n66124), .Y(n66128) );
  INVX1 U69723 ( .A(n66125), .Y(n66133) );
  NAND2X1 U69724 ( .A(n66133), .B(n66126), .Y(n66127) );
  NOR2X1 U69725 ( .A(n66128), .B(n66127), .Y(n66130) );
  NOR2X1 U69726 ( .A(n71845), .B(n72365), .Y(n66129) );
  NOR2X1 U69727 ( .A(n66130), .B(n66129), .Y(n66138) );
  NOR2X1 U69728 ( .A(n71844), .B(n72364), .Y(n66136) );
  NOR2X1 U69729 ( .A(n66132), .B(n66131), .Y(n66134) );
  NAND2X1 U69730 ( .A(n66134), .B(n66133), .Y(n66135) );
  NAND2X1 U69731 ( .A(n66136), .B(n66135), .Y(n66137) );
  NAND2X1 U69732 ( .A(n66138), .B(n66137), .Y(n71848) );
  INVX1 U69733 ( .A(n71848), .Y(n66727) );
  XNOR2X1 U69734 ( .A(n71847), .B(n66727), .Y(n67084) );
  INVX1 U69735 ( .A(n67084), .Y(n66723) );
  NAND2X1 U69736 ( .A(n66139), .B(n71847), .Y(n66140) );
  NAND2X1 U69737 ( .A(n66141), .B(n66140), .Y(n66375) );
  INVX1 U69738 ( .A(n66743), .Y(n66388) );
  NOR2X1 U69739 ( .A(n43520), .B(n43886), .Y(n66142) );
  XOR2X1 U69740 ( .A(n66388), .B(n66142), .Y(n66401) );
  XNOR2X1 U69741 ( .A(n66398), .B(n66401), .Y(n66143) );
  NAND2X1 U69742 ( .A(n66400), .B(n66399), .Y(n66404) );
  INVX1 U69743 ( .A(n66404), .Y(n66145) );
  NOR2X1 U69744 ( .A(n66145), .B(n66144), .Y(n66146) );
  NOR2X1 U69745 ( .A(n66146), .B(n66402), .Y(n66153) );
  NAND2X1 U69746 ( .A(n66150), .B(n66149), .Y(n66151) );
  NAND2X1 U69747 ( .A(n66151), .B(n66404), .Y(n66152) );
  NAND2X1 U69748 ( .A(n66153), .B(n66152), .Y(n66755) );
  NAND2X1 U69749 ( .A(n43896), .B(n43496), .Y(n66361) );
  NAND2X1 U69750 ( .A(n43492), .B(n43904), .Y(n66700) );
  XNOR2X1 U69751 ( .A(n66361), .B(n66700), .Y(n66154) );
  XNOR2X1 U69752 ( .A(n38679), .B(n66330), .Y(n66339) );
  INVX1 U69753 ( .A(n66339), .Y(n66341) );
  XNOR2X1 U69754 ( .A(n66155), .B(n66341), .Y(n66156) );
  XNOR2X1 U69755 ( .A(n41424), .B(n66156), .Y(n66322) );
  NAND2X1 U69756 ( .A(n43933), .B(n43775), .Y(n66442) );
  NAND2X1 U69757 ( .A(n43928), .B(n43478), .Y(n66323) );
  INVX1 U69758 ( .A(n66323), .Y(n66437) );
  XNOR2X1 U69759 ( .A(n66442), .B(n66437), .Y(n66157) );
  XNOR2X1 U69760 ( .A(n66322), .B(n66157), .Y(n66158) );
  XNOR2X1 U69761 ( .A(n66682), .B(n66158), .Y(n66159) );
  XNOR2X1 U69762 ( .A(n41123), .B(n66159), .Y(n66446) );
  XNOR2X1 U69763 ( .A(n66456), .B(n66446), .Y(n66160) );
  XNOR2X1 U69764 ( .A(n66462), .B(n41518), .Y(n66173) );
  INVX1 U69765 ( .A(n66162), .Y(n66166) );
  INVX1 U69766 ( .A(n66164), .Y(n66165) );
  NOR2X1 U69767 ( .A(n66166), .B(n66165), .Y(n66170) );
  NAND2X1 U69768 ( .A(n66168), .B(n66167), .Y(n66169) );
  NAND2X1 U69769 ( .A(n66170), .B(n66169), .Y(n66172) );
  INVX1 U69770 ( .A(n66319), .Y(n66820) );
  INVX1 U69771 ( .A(n66174), .Y(n66175) );
  NAND2X1 U69772 ( .A(n66177), .B(n66176), .Y(n66316) );
  INVX1 U69773 ( .A(n66314), .Y(n66836) );
  XNOR2X1 U69774 ( .A(n66839), .B(n66836), .Y(n66200) );
  INVX1 U69775 ( .A(n66178), .Y(n66196) );
  NOR2X1 U69776 ( .A(n66181), .B(n66180), .Y(n66182) );
  NOR2X1 U69777 ( .A(n41375), .B(n66182), .Y(n66186) );
  NAND2X1 U69778 ( .A(n66186), .B(n66185), .Y(n66188) );
  NAND2X1 U69779 ( .A(n66188), .B(n66187), .Y(n66191) );
  NAND2X1 U69780 ( .A(n43977), .B(n66189), .Y(n66190) );
  NAND2X1 U69781 ( .A(n66191), .B(n66190), .Y(n66194) );
  NAND2X1 U69782 ( .A(n66192), .B(n43973), .Y(n66193) );
  NAND2X1 U69783 ( .A(n66193), .B(n66194), .Y(n66195) );
  NOR2X1 U69784 ( .A(n41399), .B(n41175), .Y(n66199) );
  NAND2X1 U69785 ( .A(n66198), .B(n66197), .Y(n66311) );
  NAND2X1 U69786 ( .A(n66199), .B(n66311), .Y(n66840) );
  INVX1 U69787 ( .A(n66840), .Y(n66835) );
  XNOR2X1 U69788 ( .A(n66200), .B(n66835), .Y(n66666) );
  INVX1 U69789 ( .A(n66666), .Y(n66309) );
  INVX1 U69790 ( .A(n66201), .Y(n66202) );
  NAND2X1 U69791 ( .A(n66204), .B(n66203), .Y(n66304) );
  NAND2X1 U69792 ( .A(n43787), .B(n44026), .Y(n66473) );
  NAND2X1 U69793 ( .A(n42638), .B(n44008), .Y(n66645) );
  INVX1 U69794 ( .A(n66645), .Y(n66644) );
  NAND2X1 U69795 ( .A(n43724), .B(n44017), .Y(n66978) );
  INVX1 U69796 ( .A(n66978), .Y(n66298) );
  XNOR2X1 U69797 ( .A(n66644), .B(n66298), .Y(n66480) );
  XNOR2X1 U69798 ( .A(n66473), .B(n66480), .Y(n66208) );
  XOR2X1 U69799 ( .A(n66482), .B(n66208), .Y(n66209) );
  NAND2X1 U69800 ( .A(n40485), .B(n44049), .Y(n66868) );
  INVX1 U69801 ( .A(n66868), .Y(n66493) );
  NAND2X1 U69802 ( .A(n40473), .B(n44056), .Y(n67183) );
  INVX1 U69803 ( .A(n67183), .Y(n67186) );
  XNOR2X1 U69804 ( .A(n66288), .B(n67186), .Y(n66210) );
  INVX1 U69805 ( .A(n66285), .Y(n66284) );
  XNOR2X1 U69806 ( .A(n70752), .B(n66284), .Y(n66211) );
  XNOR2X1 U69807 ( .A(n66281), .B(n66211), .Y(n66505) );
  XNOR2X1 U69808 ( .A(n43628), .B(n66505), .Y(n66212) );
  XOR2X1 U69809 ( .A(n66504), .B(n66212), .Y(n66513) );
  XNOR2X1 U69810 ( .A(n39659), .B(n43566), .Y(n66213) );
  XNOR2X1 U69811 ( .A(n41322), .B(n66213), .Y(n66214) );
  NAND2X1 U69812 ( .A(n66215), .B(n66608), .Y(n66512) );
  XNOR2X1 U69813 ( .A(n66512), .B(n43546), .Y(n66216) );
  NAND2X1 U69814 ( .A(n43545), .B(n66519), .Y(n66217) );
  NAND2X1 U69815 ( .A(n66217), .B(n66514), .Y(n66218) );
  NOR2X1 U69816 ( .A(n41052), .B(n66218), .Y(n66221) );
  NAND2X1 U69817 ( .A(n66219), .B(n66517), .Y(n66220) );
  NAND2X1 U69818 ( .A(n66221), .B(n66220), .Y(n66223) );
  NAND2X1 U69819 ( .A(n66223), .B(n66523), .Y(n66225) );
  NAND2X1 U69820 ( .A(n43545), .B(n66224), .Y(n66525) );
  XNOR2X1 U69821 ( .A(n41071), .B(n41032), .Y(n66599) );
  INVX1 U69822 ( .A(n66599), .Y(n66271) );
  XNOR2X1 U69823 ( .A(n69861), .B(n66271), .Y(n66226) );
  XNOR2X1 U69824 ( .A(n41068), .B(n66226), .Y(n66529) );
  XNOR2X1 U69825 ( .A(n43649), .B(n66529), .Y(n66227) );
  XOR2X1 U69826 ( .A(n66530), .B(n66227), .Y(n66258) );
  NAND2X1 U69827 ( .A(n39018), .B(n43647), .Y(n66228) );
  XNOR2X1 U69828 ( .A(n66257), .B(n43654), .Y(n66229) );
  XNOR2X1 U69829 ( .A(n66230), .B(n41126), .Y(n66231) );
  XNOR2X1 U69830 ( .A(n41137), .B(n66231), .Y(n66255) );
  XNOR2X1 U69831 ( .A(n66255), .B(n43679), .Y(n66235) );
  INVX1 U69832 ( .A(n66233), .Y(n66232) );
  NAND2X1 U69833 ( .A(n66232), .B(n43685), .Y(n66576) );
  NAND2X1 U69834 ( .A(n43677), .B(n66233), .Y(n66234) );
  NAND2X1 U69835 ( .A(n66576), .B(n66577), .Y(n66254) );
  XNOR2X1 U69836 ( .A(n66251), .B(n43509), .Y(n66236) );
  INVX1 U69837 ( .A(n66554), .Y(n66551) );
  XNOR2X1 U69838 ( .A(n43709), .B(n66551), .Y(n66244) );
  INVX1 U69839 ( .A(n66237), .Y(n66239) );
  NOR2X1 U69840 ( .A(n43707), .B(n66242), .Y(n66238) );
  NOR2X1 U69841 ( .A(n66239), .B(n66238), .Y(n66241) );
  INVX1 U69842 ( .A(n66552), .Y(n66243) );
  XNOR2X1 U69843 ( .A(n66244), .B(n66243), .Y(n66249) );
  XNOR2X1 U69844 ( .A(n66246), .B(n66245), .Y(n66247) );
  XNOR2X1 U69845 ( .A(n66247), .B(n41969), .Y(n66248) );
  MX2X1 U69846 ( .A(n66249), .B(n66248), .S0(n43719), .Y(u_muldiv_result_r[12]) );
  NAND2X1 U69847 ( .A(u_muldiv_mult_result_q[12]), .B(n44632), .Y(n14027) );
  INVX1 U69848 ( .A(n66251), .Y(n66250) );
  NAND2X1 U69849 ( .A(n66251), .B(n43513), .Y(n66253) );
  NAND2X1 U69850 ( .A(n66254), .B(n66573), .Y(n66256) );
  NAND2X1 U69851 ( .A(n66255), .B(n43685), .Y(n66578) );
  XNOR2X1 U69852 ( .A(n43509), .B(n41217), .Y(n66544) );
  NOR2X1 U69853 ( .A(n41076), .B(n43661), .Y(n66260) );
  NOR2X1 U69854 ( .A(n39980), .B(n66260), .Y(n66262) );
  INVX1 U69855 ( .A(n66585), .Y(n66896) );
  XNOR2X1 U69856 ( .A(n43524), .B(n66896), .Y(n66539) );
  XNOR2X1 U69857 ( .A(n43633), .B(n41071), .Y(n66263) );
  XNOR2X1 U69858 ( .A(n66263), .B(n41032), .Y(n66264) );
  XNOR2X1 U69859 ( .A(n41068), .B(n66264), .Y(n66268) );
  INVX1 U69860 ( .A(n66268), .Y(n66265) );
  NAND2X1 U69861 ( .A(n43664), .B(n66268), .Y(n66269) );
  NOR2X1 U69862 ( .A(n40436), .B(n66271), .Y(n66273) );
  NAND2X1 U69863 ( .A(n66272), .B(n66273), .Y(n66604) );
  NAND2X1 U69864 ( .A(n66275), .B(n66274), .Y(n66276) );
  NAND2X1 U69865 ( .A(n66276), .B(n43637), .Y(n66277) );
  XNOR2X1 U69866 ( .A(n43537), .B(n66278), .Y(n66279) );
  XNOR2X1 U69867 ( .A(n66279), .B(n41347), .Y(n66280) );
  NAND2X1 U69868 ( .A(n38263), .B(n43560), .Y(n66283) );
  NAND2X1 U69869 ( .A(n66285), .B(n43538), .Y(n66287) );
  XNOR2X1 U69870 ( .A(n66488), .B(n66493), .Y(n66288) );
  XNOR2X1 U69871 ( .A(n66288), .B(n39845), .Y(n66289) );
  XNOR2X1 U69872 ( .A(n39715), .B(n66289), .Y(n67185) );
  INVX1 U69873 ( .A(n67185), .Y(n66290) );
  NOR2X1 U69874 ( .A(n66290), .B(n67183), .Y(n66297) );
  NAND2X1 U69875 ( .A(n66626), .B(n66291), .Y(n66292) );
  NAND2X1 U69876 ( .A(n67185), .B(n66292), .Y(n67187) );
  NAND2X1 U69877 ( .A(n38888), .B(n66293), .Y(n67179) );
  NAND2X1 U69878 ( .A(n66294), .B(n67179), .Y(n66627) );
  NAND2X1 U69879 ( .A(n66295), .B(n67187), .Y(n66296) );
  NOR2X1 U69880 ( .A(n66297), .B(n66296), .Y(n66611) );
  XNOR2X1 U69881 ( .A(n43537), .B(n66611), .Y(n66502) );
  NOR2X1 U69882 ( .A(n38393), .B(n39994), .Y(n66299) );
  NAND2X1 U69883 ( .A(n66298), .B(n40530), .Y(n66954) );
  NAND2X1 U69884 ( .A(n66954), .B(n36684), .Y(n66984) );
  INVX1 U69885 ( .A(n66646), .Y(n66300) );
  NOR2X1 U69886 ( .A(n66300), .B(n38522), .Y(n66301) );
  NOR2X1 U69887 ( .A(n66301), .B(n66647), .Y(n66303) );
  NAND2X1 U69888 ( .A(n66644), .B(n66646), .Y(n66302) );
  NOR2X1 U69889 ( .A(n41645), .B(n41618), .Y(n66305) );
  NAND2X1 U69890 ( .A(n66305), .B(n66304), .Y(n66668) );
  NOR2X1 U69891 ( .A(n66666), .B(n66659), .Y(n66306) );
  NOR2X1 U69892 ( .A(n66307), .B(n66306), .Y(n66310) );
  NOR2X1 U69893 ( .A(n41399), .B(n41175), .Y(n66312) );
  NAND2X1 U69894 ( .A(n66312), .B(n66311), .Y(n66315) );
  NOR2X1 U69895 ( .A(n40978), .B(n40981), .Y(n66317) );
  NAND2X1 U69896 ( .A(n66820), .B(n66318), .Y(n66822) );
  OR2X1 U69897 ( .A(n66319), .B(n66819), .Y(n66320) );
  NOR2X1 U69898 ( .A(n36682), .B(n36683), .Y(n66818) );
  NAND2X1 U69899 ( .A(n43795), .B(n43973), .Y(n66798) );
  NAND2X1 U69900 ( .A(n43942), .B(n43775), .Y(n67024) );
  NAND2X1 U69901 ( .A(n66438), .B(n66323), .Y(n67339) );
  NAND2X1 U69902 ( .A(n41196), .B(n67339), .Y(n66324) );
  NOR2X1 U69903 ( .A(n67024), .B(n66324), .Y(n66326) );
  NOR2X1 U69904 ( .A(n67024), .B(n40247), .Y(n66325) );
  NOR2X1 U69905 ( .A(n66326), .B(n66325), .Y(n66329) );
  INVX1 U69906 ( .A(n67024), .Y(n66676) );
  NOR2X1 U69907 ( .A(n66676), .B(n40287), .Y(n66327) );
  NAND2X1 U69908 ( .A(n66327), .B(n66324), .Y(n66328) );
  NAND2X1 U69909 ( .A(n66329), .B(n66328), .Y(n66436) );
  NAND2X1 U69910 ( .A(n43933), .B(n43478), .Y(n67341) );
  XNOR2X1 U69911 ( .A(n38679), .B(n66342), .Y(n66331) );
  XNOR2X1 U69912 ( .A(n66331), .B(n66330), .Y(n66332) );
  XNOR2X1 U69913 ( .A(n41424), .B(n66332), .Y(n66683) );
  NAND2X1 U69914 ( .A(n66683), .B(n66682), .Y(n67040) );
  NAND2X1 U69915 ( .A(n66334), .B(n66333), .Y(n66335) );
  OR2X1 U69916 ( .A(n66683), .B(n66335), .Y(n66336) );
  NAND2X1 U69917 ( .A(n66337), .B(n66336), .Y(n67039) );
  NAND2X1 U69918 ( .A(n67040), .B(n67039), .Y(n66681) );
  NAND2X1 U69919 ( .A(n66340), .B(n66339), .Y(n67056) );
  NAND2X1 U69920 ( .A(n38855), .B(n67056), .Y(n67062) );
  NAND2X1 U69921 ( .A(n66342), .B(n66341), .Y(n67063) );
  INVX1 U69922 ( .A(n67063), .Y(n66343) );
  NOR2X1 U69923 ( .A(n38156), .B(n66343), .Y(n66349) );
  NOR2X1 U69924 ( .A(n38857), .B(n67057), .Y(n66347) );
  NAND2X1 U69925 ( .A(n66347), .B(n67056), .Y(n66348) );
  NAND2X1 U69926 ( .A(n66349), .B(n66348), .Y(n66788) );
  NAND2X1 U69927 ( .A(n43927), .B(n43484), .Y(n67033) );
  NAND2X1 U69928 ( .A(n43903), .B(n43497), .Y(n67121) );
  INVX1 U69929 ( .A(n67121), .Y(n66768) );
  NOR2X1 U69930 ( .A(n43894), .B(n66361), .Y(n66352) );
  INVX1 U69931 ( .A(n66357), .Y(n66350) );
  NAND2X1 U69932 ( .A(n41220), .B(n66350), .Y(n66351) );
  NAND2X1 U69933 ( .A(n66352), .B(n66351), .Y(n66354) );
  INVX1 U69934 ( .A(n66361), .Y(n66413) );
  INVX1 U69935 ( .A(n66362), .Y(n66412) );
  NAND2X1 U69936 ( .A(n66413), .B(n66412), .Y(n66353) );
  NAND2X1 U69937 ( .A(n66354), .B(n66353), .Y(n66764) );
  NOR2X1 U69938 ( .A(n66362), .B(n66355), .Y(n66359) );
  OR2X1 U69939 ( .A(n66357), .B(n66356), .Y(n66358) );
  INVX1 U69940 ( .A(n66360), .Y(n66364) );
  NAND2X1 U69941 ( .A(n66362), .B(n66361), .Y(n66363) );
  NOR2X1 U69942 ( .A(n66764), .B(n66761), .Y(n66365) );
  XNOR2X1 U69943 ( .A(n66768), .B(n66365), .Y(n66697) );
  NAND2X1 U69944 ( .A(n43492), .B(n43912), .Y(n66691) );
  NAND2X1 U69945 ( .A(n66388), .B(n66745), .Y(n66381) );
  INVX1 U69946 ( .A(n66381), .Y(n66380) );
  NAND2X1 U69947 ( .A(n43889), .B(n39960), .Y(n67091) );
  INVX1 U69948 ( .A(n67091), .Y(n66742) );
  NAND2X1 U69949 ( .A(n43879), .B(n43607), .Y(n66717) );
  INVX1 U69950 ( .A(n66366), .Y(n66377) );
  NAND2X1 U69951 ( .A(n66377), .B(n43604), .Y(n72366) );
  NAND2X1 U69952 ( .A(n41853), .B(n71845), .Y(n66368) );
  INVX1 U69953 ( .A(n72366), .Y(n71843) );
  NAND2X1 U69954 ( .A(n71843), .B(n72365), .Y(n66367) );
  NAND2X1 U69955 ( .A(n66368), .B(n66367), .Y(n66373) );
  NAND2X1 U69956 ( .A(n41853), .B(n66725), .Y(n66371) );
  NOR2X1 U69957 ( .A(n71845), .B(n72366), .Y(n66369) );
  NAND2X1 U69958 ( .A(n66369), .B(n71847), .Y(n66370) );
  NAND2X1 U69959 ( .A(n66371), .B(n66370), .Y(n66372) );
  NOR2X1 U69960 ( .A(n66373), .B(n66372), .Y(n66374) );
  XNOR2X1 U69961 ( .A(n66723), .B(n66374), .Y(n67421) );
  INVX1 U69962 ( .A(n67421), .Y(n67426) );
  XNOR2X1 U69963 ( .A(n66717), .B(n67426), .Y(n66378) );
  NAND2X1 U69964 ( .A(n66375), .B(n67084), .Y(n66376) );
  NAND2X1 U69965 ( .A(n66377), .B(n66376), .Y(n66718) );
  INVX1 U69966 ( .A(n66394), .Y(n66391) );
  NOR2X1 U69967 ( .A(n66391), .B(n43882), .Y(n66379) );
  NOR2X1 U69968 ( .A(n66380), .B(n66379), .Y(n66383) );
  NOR2X1 U69969 ( .A(n66391), .B(n66381), .Y(n66382) );
  NOR2X1 U69970 ( .A(n66383), .B(n66382), .Y(n66393) );
  INVX1 U69971 ( .A(n66384), .Y(n66386) );
  NOR2X1 U69972 ( .A(n66386), .B(n66385), .Y(n66387) );
  NOR2X1 U69973 ( .A(n66388), .B(n66387), .Y(n66390) );
  NAND2X1 U69974 ( .A(n66390), .B(n66389), .Y(n66734) );
  NAND2X1 U69975 ( .A(n66734), .B(n39961), .Y(n67096) );
  INVX1 U69976 ( .A(n67096), .Y(n67406) );
  NOR2X1 U69977 ( .A(n66391), .B(n67406), .Y(n66392) );
  NOR2X1 U69978 ( .A(n66393), .B(n66392), .Y(n66397) );
  NOR2X1 U69979 ( .A(n43884), .B(n66394), .Y(n66395) );
  NAND2X1 U69980 ( .A(n67406), .B(n66395), .Y(n66396) );
  NAND2X1 U69981 ( .A(n66397), .B(n66396), .Y(n67108) );
  NAND2X1 U69982 ( .A(n43896), .B(n43501), .Y(n66753) );
  INVX1 U69983 ( .A(n66753), .Y(n67110) );
  XNOR2X1 U69984 ( .A(n67108), .B(n67110), .Y(n66409) );
  INVX1 U69985 ( .A(n66398), .Y(n66751) );
  NOR2X1 U69986 ( .A(n66400), .B(n66399), .Y(n66402) );
  NOR2X1 U69987 ( .A(n66402), .B(n66752), .Y(n66406) );
  NAND2X1 U69988 ( .A(n66404), .B(n66403), .Y(n66405) );
  NAND2X1 U69989 ( .A(n66406), .B(n66405), .Y(n66750) );
  NAND2X1 U69990 ( .A(n66751), .B(n66750), .Y(n66408) );
  NAND2X1 U69991 ( .A(n66752), .B(n66755), .Y(n66407) );
  NAND2X1 U69992 ( .A(n66408), .B(n66407), .Y(n67109) );
  XNOR2X1 U69993 ( .A(n66691), .B(n67122), .Y(n66410) );
  XOR2X1 U69994 ( .A(n66697), .B(n66410), .Y(n66786) );
  NOR2X1 U69995 ( .A(n66417), .B(n66411), .Y(n66414) );
  XNOR2X1 U69996 ( .A(n66413), .B(n66412), .Y(n66701) );
  NOR2X1 U69997 ( .A(n66414), .B(n66690), .Y(n66421) );
  INVX1 U69998 ( .A(n66415), .Y(n66419) );
  NOR2X1 U69999 ( .A(n66417), .B(n66416), .Y(n66418) );
  NOR2X1 U70000 ( .A(n66419), .B(n66418), .Y(n66420) );
  NAND2X1 U70001 ( .A(n66421), .B(n66420), .Y(n66713) );
  INVX1 U70002 ( .A(n66713), .Y(n66422) );
  NOR2X1 U70003 ( .A(n66422), .B(n66700), .Y(n66425) );
  NAND2X1 U70004 ( .A(n66690), .B(n66423), .Y(n66784) );
  NAND2X1 U70005 ( .A(n43919), .B(n38310), .Y(n66427) );
  NAND2X1 U70006 ( .A(n66784), .B(n66427), .Y(n66424) );
  NOR2X1 U70007 ( .A(n66425), .B(n66424), .Y(n66432) );
  INVX1 U70008 ( .A(n66784), .Y(n66426) );
  INVX1 U70009 ( .A(n66427), .Y(n67069) );
  NAND2X1 U70010 ( .A(n66426), .B(n67069), .Y(n66430) );
  NOR2X1 U70011 ( .A(n66700), .B(n66427), .Y(n66428) );
  NAND2X1 U70012 ( .A(n66428), .B(n66713), .Y(n66429) );
  NAND2X1 U70013 ( .A(n66430), .B(n66429), .Y(n66431) );
  NOR2X1 U70014 ( .A(n66432), .B(n66431), .Y(n66433) );
  XNOR2X1 U70015 ( .A(n66786), .B(n66433), .Y(n66680) );
  XNOR2X1 U70016 ( .A(n67033), .B(n66680), .Y(n66434) );
  INVX1 U70017 ( .A(n67344), .Y(n66675) );
  XNOR2X1 U70018 ( .A(n67341), .B(n66675), .Y(n66435) );
  XNOR2X1 U70019 ( .A(n66436), .B(n66435), .Y(n66445) );
  NAND2X1 U70020 ( .A(n40122), .B(n66442), .Y(n66441) );
  XNOR2X1 U70021 ( .A(n66438), .B(n66437), .Y(n66439) );
  XNOR2X1 U70022 ( .A(n41123), .B(n66439), .Y(n66440) );
  INVX1 U70023 ( .A(n66442), .Y(n66444) );
  NAND2X1 U70024 ( .A(n66457), .B(n66456), .Y(n66455) );
  INVX1 U70025 ( .A(n66447), .Y(n66449) );
  NAND2X1 U70026 ( .A(n66449), .B(n66448), .Y(n66451) );
  NAND2X1 U70027 ( .A(n66451), .B(n66450), .Y(n66453) );
  NAND2X1 U70028 ( .A(n66453), .B(n66452), .Y(n66454) );
  NAND2X1 U70029 ( .A(n66455), .B(n66454), .Y(n66461) );
  INVX1 U70030 ( .A(n66456), .Y(n66459) );
  INVX1 U70031 ( .A(n66457), .Y(n66458) );
  NAND2X1 U70032 ( .A(n66459), .B(n66458), .Y(n66460) );
  NAND2X1 U70033 ( .A(n66461), .B(n66460), .Y(n66799) );
  INVX1 U70034 ( .A(n66816), .Y(n66805) );
  NOR2X1 U70035 ( .A(n41205), .B(n41209), .Y(n66464) );
  NAND2X1 U70036 ( .A(n41518), .B(n66463), .Y(n66806) );
  NAND2X1 U70037 ( .A(n66464), .B(n66806), .Y(n66817) );
  INVX1 U70038 ( .A(n66817), .Y(n66465) );
  XNOR2X1 U70039 ( .A(n66805), .B(n66465), .Y(n66467) );
  NAND2X1 U70040 ( .A(n42711), .B(n43983), .Y(n66815) );
  NAND2X1 U70041 ( .A(n42661), .B(n43992), .Y(n66825) );
  INVX1 U70042 ( .A(n66825), .Y(n66831) );
  XNOR2X1 U70043 ( .A(n66815), .B(n66831), .Y(n66466) );
  XNOR2X1 U70044 ( .A(n66467), .B(n66466), .Y(n66468) );
  XNOR2X1 U70045 ( .A(n66818), .B(n66468), .Y(n66834) );
  NAND2X1 U70046 ( .A(n43772), .B(n44008), .Y(n66658) );
  NAND2X1 U70047 ( .A(n43798), .B(n44000), .Y(n66833) );
  XNOR2X1 U70048 ( .A(n66658), .B(n66833), .Y(n66469) );
  XOR2X1 U70049 ( .A(n66834), .B(n66469), .Y(n66470) );
  XNOR2X1 U70050 ( .A(n41763), .B(n66640), .Y(n66654) );
  INVX1 U70051 ( .A(n66654), .Y(n66651) );
  XNOR2X1 U70052 ( .A(n41573), .B(n66651), .Y(n66472) );
  NAND2X1 U70053 ( .A(n42639), .B(n44017), .Y(n66650) );
  NAND2X1 U70054 ( .A(n43725), .B(n44026), .Y(n66643) );
  INVX1 U70055 ( .A(n66643), .Y(n66953) );
  XNOR2X1 U70056 ( .A(n66650), .B(n66953), .Y(n66471) );
  INVX1 U70057 ( .A(n66473), .Y(n66483) );
  NAND2X1 U70058 ( .A(n44020), .B(n66474), .Y(n66477) );
  NAND2X1 U70059 ( .A(n66483), .B(n66479), .Y(n66851) );
  XNOR2X1 U70060 ( .A(n66646), .B(n66480), .Y(n66481) );
  NAND2X1 U70061 ( .A(n40486), .B(n44056), .Y(n66878) );
  NAND2X1 U70062 ( .A(n43787), .B(n44048), .Y(n66637) );
  INVX1 U70063 ( .A(n66637), .Y(n66850) );
  XNOR2X1 U70064 ( .A(n66878), .B(n66850), .Y(n66486) );
  XNOR2X1 U70065 ( .A(n66964), .B(n66486), .Y(n66487) );
  XNOR2X1 U70066 ( .A(n66972), .B(n66487), .Y(n66623) );
  XNOR2X1 U70067 ( .A(n43574), .B(n66623), .Y(n66501) );
  XNOR2X1 U70068 ( .A(n66488), .B(n39845), .Y(n66879) );
  OR2X1 U70069 ( .A(n66879), .B(n66868), .Y(n66491) );
  NAND2X1 U70070 ( .A(n66493), .B(n39171), .Y(n66489) );
  OR2X1 U70071 ( .A(n40077), .B(n66489), .Y(n66490) );
  NAND2X1 U70072 ( .A(n66491), .B(n66490), .Y(n66500) );
  OR2X1 U70073 ( .A(n66879), .B(n66492), .Y(n66498) );
  NOR2X1 U70074 ( .A(n66493), .B(n39309), .Y(n66496) );
  NAND2X1 U70075 ( .A(n66874), .B(n66873), .Y(n66495) );
  OR2X1 U70076 ( .A(n66496), .B(n66495), .Y(n66497) );
  NAND2X1 U70077 ( .A(n66498), .B(n66497), .Y(n66499) );
  NOR2X1 U70078 ( .A(n66500), .B(n66499), .Y(n66622) );
  XNOR2X1 U70079 ( .A(n66502), .B(n41366), .Y(n66503) );
  XNOR2X1 U70080 ( .A(n38606), .B(n66503), .Y(n66616) );
  INVX1 U70081 ( .A(n66215), .Y(n66509) );
  NAND2X1 U70082 ( .A(n66608), .B(n66609), .Y(n66508) );
  NOR2X1 U70083 ( .A(n66509), .B(n66508), .Y(n66510) );
  NOR2X1 U70084 ( .A(n36763), .B(n66510), .Y(n66888) );
  XNOR2X1 U70085 ( .A(n66888), .B(n43553), .Y(n66511) );
  INVX1 U70086 ( .A(n66514), .Y(n66515) );
  NOR2X1 U70087 ( .A(n41052), .B(n66515), .Y(n66522) );
  NAND2X1 U70088 ( .A(n66517), .B(n66516), .Y(n66518) );
  NAND2X1 U70089 ( .A(n66518), .B(n43550), .Y(n66520) );
  NAND2X1 U70090 ( .A(n66520), .B(n66519), .Y(n66521) );
  NAND2X1 U70091 ( .A(n66522), .B(n66521), .Y(n66524) );
  NAND2X1 U70092 ( .A(n66524), .B(n66523), .Y(n67204) );
  XNOR2X1 U70093 ( .A(n41334), .B(n41049), .Y(n66605) );
  XNOR2X1 U70094 ( .A(n66596), .B(n66527), .Y(n66587) );
  XNOR2X1 U70095 ( .A(n43650), .B(n66587), .Y(n66528) );
  XOR2X1 U70096 ( .A(n67222), .B(n66528), .Y(n66582) );
  INVX1 U70097 ( .A(n66531), .Y(n66532) );
  NAND2X1 U70098 ( .A(n66532), .B(n66535), .Y(n66533) );
  NOR2X1 U70099 ( .A(n41335), .B(n39670), .Y(n66537) );
  NAND2X1 U70100 ( .A(n66537), .B(n66589), .Y(n66581) );
  XNOR2X1 U70101 ( .A(n66581), .B(n43654), .Y(n66538) );
  XNOR2X1 U70102 ( .A(n66539), .B(n41128), .Y(n66543) );
  XNOR2X1 U70103 ( .A(n41107), .B(n41126), .Y(n66540) );
  NOR2X1 U70104 ( .A(n41106), .B(n41137), .Y(n66541) );
  NOR2X1 U70105 ( .A(n41413), .B(n66541), .Y(n66542) );
  XNOR2X1 U70106 ( .A(n66543), .B(n66542), .Y(n66580) );
  XNOR2X1 U70107 ( .A(n66544), .B(n41216), .Y(n66545) );
  XNOR2X1 U70108 ( .A(n66567), .B(n43693), .Y(n66550) );
  NAND2X1 U70109 ( .A(n43691), .B(n66548), .Y(n66547) );
  NOR2X1 U70110 ( .A(n41219), .B(n41465), .Y(n66549) );
  XNOR2X1 U70111 ( .A(n66550), .B(n66549), .Y(n66564) );
  INVX1 U70112 ( .A(n66564), .Y(n66562) );
  XNOR2X1 U70113 ( .A(n43709), .B(n66562), .Y(n66556) );
  NAND2X1 U70114 ( .A(n66551), .B(n43712), .Y(n66553) );
  NAND2X1 U70115 ( .A(n43706), .B(n66554), .Y(n66916) );
  NAND2X1 U70116 ( .A(n37908), .B(n66916), .Y(n66563) );
  INVX1 U70117 ( .A(n66563), .Y(n66555) );
  XNOR2X1 U70118 ( .A(n66556), .B(n66555), .Y(n66561) );
  XNOR2X1 U70119 ( .A(n66558), .B(n66557), .Y(n66559) );
  XNOR2X1 U70120 ( .A(n41979), .B(n66559), .Y(n66560) );
  MX2X1 U70121 ( .A(n66561), .B(n66560), .S0(n43719), .Y(u_muldiv_result_r[13]) );
  NAND2X1 U70122 ( .A(u_muldiv_mult_result_q[13]), .B(n44632), .Y(n14016) );
  NAND2X1 U70123 ( .A(n66563), .B(n66913), .Y(n66565) );
  NAND2X1 U70124 ( .A(n66565), .B(n37915), .Y(n66907) );
  INVX1 U70125 ( .A(n66567), .Y(n66566) );
  NAND2X1 U70126 ( .A(n43691), .B(n66567), .Y(n66568) );
  NAND2X1 U70127 ( .A(n37886), .B(n66568), .Y(n66919) );
  XNOR2X1 U70128 ( .A(n41217), .B(n41216), .Y(n66572) );
  NAND2X1 U70129 ( .A(n66572), .B(n43512), .Y(n66571) );
  NAND2X1 U70130 ( .A(n66921), .B(n39510), .Y(n66904) );
  NOR2X1 U70131 ( .A(n43687), .B(n66580), .Y(n66575) );
  INVX1 U70132 ( .A(n66573), .Y(n66574) );
  NAND2X1 U70133 ( .A(n66578), .B(n66577), .Y(n66579) );
  NAND2X1 U70134 ( .A(n66580), .B(n43683), .Y(n67249) );
  NAND2X1 U70135 ( .A(n66583), .B(n43659), .Y(n67584) );
  INVX1 U70136 ( .A(n66583), .Y(n66584) );
  NAND2X1 U70137 ( .A(n43655), .B(n66584), .Y(n66586) );
  NAND2X1 U70138 ( .A(n66591), .B(n66590), .Y(n66592) );
  XNOR2X1 U70139 ( .A(n43633), .B(n41334), .Y(n66594) );
  XNOR2X1 U70140 ( .A(n66594), .B(n41049), .Y(n66595) );
  XNOR2X1 U70141 ( .A(n66596), .B(n66595), .Y(n66597) );
  NAND2X1 U70142 ( .A(n67223), .B(n67222), .Y(n67273) );
  NAND2X1 U70143 ( .A(n66597), .B(n43669), .Y(n67224) );
  NAND2X1 U70144 ( .A(n67273), .B(n67224), .Y(n66932) );
  XNOR2X1 U70145 ( .A(n43667), .B(n43643), .Y(n70762) );
  NOR2X1 U70146 ( .A(n43632), .B(n41334), .Y(n66603) );
  NAND2X1 U70147 ( .A(n66598), .B(n43637), .Y(n66601) );
  NAND2X1 U70148 ( .A(n66599), .B(n43637), .Y(n66600) );
  NAND2X1 U70149 ( .A(n66601), .B(n66600), .Y(n66602) );
  NOR2X1 U70150 ( .A(n66603), .B(n66602), .Y(n66607) );
  NAND2X1 U70151 ( .A(n38466), .B(n66605), .Y(n66606) );
  NAND2X1 U70152 ( .A(n66607), .B(n66606), .Y(n67220) );
  XNOR2X1 U70153 ( .A(n66611), .B(n41366), .Y(n66620) );
  INVX1 U70154 ( .A(n66620), .Y(n66619) );
  INVX1 U70155 ( .A(n70752), .Y(n72149) );
  XNOR2X1 U70156 ( .A(n66619), .B(n72149), .Y(n66612) );
  XNOR2X1 U70157 ( .A(n66612), .B(n38606), .Y(n66613) );
  INVX1 U70158 ( .A(n66614), .Y(n66615) );
  NAND2X1 U70159 ( .A(n43620), .B(n66615), .Y(n67284) );
  NAND2X1 U70160 ( .A(n67285), .B(n67284), .Y(n67212) );
  NAND2X1 U70161 ( .A(n43536), .B(n66619), .Y(n67564) );
  NAND2X1 U70162 ( .A(n67564), .B(n67563), .Y(n67198) );
  XNOR2X1 U70163 ( .A(n67198), .B(n43566), .Y(n66886) );
  NAND2X1 U70164 ( .A(n38400), .B(n66626), .Y(n66621) );
  NOR2X1 U70165 ( .A(n67185), .B(n66621), .Y(n66625) );
  XNOR2X1 U70166 ( .A(n66623), .B(n66622), .Y(n67191) );
  NOR2X1 U70167 ( .A(n67191), .B(n43574), .Y(n66624) );
  NAND2X1 U70168 ( .A(n66625), .B(n66624), .Y(n66636) );
  INVX1 U70169 ( .A(n66626), .Y(n67182) );
  NOR2X1 U70170 ( .A(n67182), .B(n36424), .Y(n66628) );
  NOR2X1 U70171 ( .A(n66628), .B(n67183), .Y(n66629) );
  NOR2X1 U70172 ( .A(n66629), .B(n67185), .Y(n66630) );
  INVX1 U70173 ( .A(n67191), .Y(n67192) );
  NOR2X1 U70174 ( .A(n66630), .B(n67192), .Y(n66634) );
  NOR2X1 U70175 ( .A(n67186), .B(n66631), .Y(n66632) );
  NOR2X1 U70176 ( .A(n43578), .B(n66632), .Y(n66633) );
  NAND2X1 U70177 ( .A(n66634), .B(n66633), .Y(n66635) );
  NAND2X1 U70178 ( .A(n66636), .B(n66635), .Y(n66939) );
  NOR2X1 U70179 ( .A(n39310), .B(n66637), .Y(n66638) );
  INVX1 U70180 ( .A(n66650), .Y(n66655) );
  XNOR2X1 U70181 ( .A(n66655), .B(n66640), .Y(n66641) );
  XNOR2X1 U70182 ( .A(n66641), .B(n41763), .Y(n66642) );
  XNOR2X1 U70183 ( .A(n41573), .B(n66642), .Y(n66986) );
  NAND2X1 U70184 ( .A(n66986), .B(n66643), .Y(n66949) );
  NAND2X1 U70185 ( .A(n66949), .B(n40331), .Y(n66992) );
  INVX1 U70186 ( .A(n66986), .Y(n66952) );
  NAND2X1 U70187 ( .A(n66953), .B(n66952), .Y(n66990) );
  NAND2X1 U70188 ( .A(n38394), .B(n66990), .Y(n66849) );
  NOR2X1 U70189 ( .A(n66644), .B(n36619), .Y(n66649) );
  NOR2X1 U70190 ( .A(n38522), .B(n66645), .Y(n66647) );
  NOR2X1 U70191 ( .A(n66647), .B(n66646), .Y(n66648) );
  NOR2X1 U70192 ( .A(n66649), .B(n66648), .Y(n66653) );
  NAND2X1 U70193 ( .A(n66651), .B(n66650), .Y(n66652) );
  NAND2X1 U70194 ( .A(n66653), .B(n66652), .Y(n66657) );
  NAND2X1 U70195 ( .A(n66655), .B(n66654), .Y(n66656) );
  NAND2X1 U70196 ( .A(n66657), .B(n66656), .Y(n67523) );
  INVX1 U70197 ( .A(n67523), .Y(n66996) );
  INVX1 U70198 ( .A(n66658), .Y(n66672) );
  NOR2X1 U70199 ( .A(n66672), .B(n66306), .Y(n66662) );
  NAND2X1 U70200 ( .A(n66659), .B(n66666), .Y(n66660) );
  NAND2X1 U70201 ( .A(n66660), .B(n66668), .Y(n66661) );
  NAND2X1 U70202 ( .A(n66662), .B(n66661), .Y(n66663) );
  NAND2X1 U70203 ( .A(n66664), .B(n66663), .Y(n67306) );
  NOR2X1 U70204 ( .A(n44005), .B(n66666), .Y(n66667) );
  NOR2X1 U70205 ( .A(n38884), .B(n66667), .Y(n66670) );
  NAND2X1 U70206 ( .A(n66668), .B(n44000), .Y(n66669) );
  NAND2X1 U70207 ( .A(n66670), .B(n66669), .Y(n66671) );
  NAND2X1 U70208 ( .A(n66672), .B(n66671), .Y(n67305) );
  NAND2X1 U70209 ( .A(n42640), .B(n44025), .Y(n67521) );
  INVX1 U70210 ( .A(n67521), .Y(n67520) );
  NAND2X1 U70211 ( .A(n42711), .B(n43992), .Y(n67493) );
  NAND2X1 U70212 ( .A(n43796), .B(n43983), .Y(n67329) );
  NAND2X1 U70213 ( .A(n66676), .B(n67026), .Y(n67030) );
  INVX1 U70214 ( .A(n67030), .Y(n66679) );
  INVX1 U70215 ( .A(n67341), .Y(n67345) );
  XNOR2X1 U70216 ( .A(n66792), .B(n67345), .Y(n66674) );
  XNOR2X1 U70217 ( .A(n66675), .B(n66674), .Y(n67025) );
  INVX1 U70218 ( .A(n67025), .Y(n66677) );
  NAND2X1 U70219 ( .A(n66677), .B(n67026), .Y(n67029) );
  NAND2X1 U70220 ( .A(n39461), .B(n67029), .Y(n66678) );
  NOR2X1 U70221 ( .A(n66679), .B(n66678), .Y(n66797) );
  INVX1 U70222 ( .A(n66686), .Y(n67042) );
  NAND2X1 U70223 ( .A(n67042), .B(n67041), .Y(n67035) );
  INVX1 U70224 ( .A(n67033), .Y(n67043) );
  NOR2X1 U70225 ( .A(n66683), .B(n66682), .Y(n66685) );
  NOR2X1 U70226 ( .A(n66685), .B(n66684), .Y(n66688) );
  NAND2X1 U70227 ( .A(n67040), .B(n66686), .Y(n66687) );
  OR2X1 U70228 ( .A(n66688), .B(n66687), .Y(n67031) );
  NAND2X1 U70229 ( .A(n67043), .B(n67031), .Y(n66689) );
  INVX1 U70230 ( .A(n66690), .Y(n66693) );
  INVX1 U70231 ( .A(n66691), .Y(n66706) );
  INVX1 U70232 ( .A(n66700), .Y(n66714) );
  NAND2X1 U70233 ( .A(n66706), .B(n66714), .Y(n66692) );
  NOR2X1 U70234 ( .A(n66693), .B(n66692), .Y(n66696) );
  INVX1 U70235 ( .A(n67122), .Y(n66766) );
  NAND2X1 U70236 ( .A(n66706), .B(n66766), .Y(n66694) );
  NOR2X1 U70237 ( .A(n66697), .B(n66694), .Y(n66695) );
  NOR2X1 U70238 ( .A(n66696), .B(n66695), .Y(n66712) );
  INVX1 U70239 ( .A(n66697), .Y(n66715) );
  NAND2X1 U70240 ( .A(n66706), .B(n67122), .Y(n66698) );
  NOR2X1 U70241 ( .A(n66715), .B(n66698), .Y(n66710) );
  NAND2X1 U70242 ( .A(n66703), .B(n66700), .Y(n66699) );
  NOR2X1 U70243 ( .A(n66701), .B(n66699), .Y(n66705) );
  NAND2X1 U70244 ( .A(n66701), .B(n66700), .Y(n66702) );
  NOR2X1 U70245 ( .A(n66703), .B(n66702), .Y(n66704) );
  NOR2X1 U70246 ( .A(n66705), .B(n66704), .Y(n66707) );
  NAND2X1 U70247 ( .A(n66707), .B(n66706), .Y(n66708) );
  NOR2X1 U70248 ( .A(n38679), .B(n66708), .Y(n66709) );
  NOR2X1 U70249 ( .A(n66710), .B(n66709), .Y(n66711) );
  NAND2X1 U70250 ( .A(n66712), .B(n66711), .Y(n67441) );
  NAND2X1 U70251 ( .A(n66714), .B(n66713), .Y(n66785) );
  NAND2X1 U70252 ( .A(n66785), .B(n66784), .Y(n66716) );
  XNOR2X1 U70253 ( .A(n66766), .B(n66715), .Y(n67077) );
  NAND2X1 U70254 ( .A(n43928), .B(n38311), .Y(n67054) );
  NAND2X1 U70255 ( .A(n43903), .B(n43501), .Y(n67395) );
  INVX1 U70256 ( .A(n67395), .Y(n67106) );
  INVX1 U70257 ( .A(n66717), .Y(n66720) );
  NAND2X1 U70258 ( .A(n66718), .B(n67426), .Y(n66719) );
  NAND2X1 U70259 ( .A(n66720), .B(n66719), .Y(n67088) );
  XNOR2X1 U70260 ( .A(n67088), .B(n41509), .Y(n66733) );
  NAND2X1 U70261 ( .A(n66720), .B(n43604), .Y(n72372) );
  NAND2X1 U70262 ( .A(n41880), .B(n71844), .Y(n66722) );
  INVX1 U70263 ( .A(n72372), .Y(n72370) );
  NAND2X1 U70264 ( .A(n72370), .B(n72366), .Y(n66721) );
  NAND2X1 U70265 ( .A(n66722), .B(n66721), .Y(n66731) );
  NAND2X1 U70266 ( .A(n41880), .B(n66723), .Y(n66729) );
  NAND2X1 U70267 ( .A(n72370), .B(n72364), .Y(n66724) );
  NOR2X1 U70268 ( .A(n66725), .B(n66724), .Y(n66726) );
  NAND2X1 U70269 ( .A(n66727), .B(n66726), .Y(n66728) );
  NAND2X1 U70270 ( .A(n66729), .B(n66728), .Y(n66730) );
  NOR2X1 U70271 ( .A(n66731), .B(n66730), .Y(n66732) );
  XNOR2X1 U70272 ( .A(n67426), .B(n66732), .Y(n67746) );
  INVX1 U70273 ( .A(n67746), .Y(n67083) );
  XNOR2X1 U70274 ( .A(n66733), .B(n67083), .Y(n67094) );
  XNOR2X1 U70275 ( .A(n67094), .B(n41708), .Y(n66749) );
  INVX1 U70276 ( .A(n66734), .Y(n66739) );
  NOR2X1 U70277 ( .A(n43884), .B(n67091), .Y(n66737) );
  NAND2X1 U70278 ( .A(n67090), .B(n43880), .Y(n66735) );
  NOR2X1 U70279 ( .A(n36706), .B(n66735), .Y(n66736) );
  NOR2X1 U70280 ( .A(n66737), .B(n66736), .Y(n66738) );
  NOR2X1 U70281 ( .A(n66739), .B(n66738), .Y(n66741) );
  NAND2X1 U70282 ( .A(n66742), .B(n67090), .Y(n67095) );
  INVX1 U70283 ( .A(n67095), .Y(n66740) );
  NOR2X1 U70284 ( .A(n66741), .B(n66740), .Y(n66748) );
  NOR2X1 U70285 ( .A(n66742), .B(n67090), .Y(n66744) );
  NOR2X1 U70286 ( .A(n66744), .B(n66743), .Y(n66746) );
  NAND2X1 U70287 ( .A(n66746), .B(n66745), .Y(n66747) );
  NAND2X1 U70288 ( .A(n66748), .B(n66747), .Y(n67098) );
  INVX1 U70289 ( .A(n67385), .Y(n67396) );
  INVX1 U70290 ( .A(n66752), .Y(n66754) );
  NOR2X1 U70291 ( .A(n66754), .B(n66753), .Y(n66756) );
  NAND2X1 U70292 ( .A(n66756), .B(n66755), .Y(n66757) );
  NAND2X1 U70293 ( .A(n67110), .B(n67108), .Y(n67102) );
  NAND2X1 U70294 ( .A(n66757), .B(n67102), .Y(n66758) );
  NOR2X1 U70295 ( .A(n66759), .B(n66758), .Y(n66760) );
  NAND2X1 U70296 ( .A(n67109), .B(n67108), .Y(n67384) );
  XNOR2X1 U70297 ( .A(n41248), .B(n41240), .Y(n67379) );
  NOR2X1 U70298 ( .A(n66766), .B(n66764), .Y(n66762) );
  INVX1 U70299 ( .A(n66761), .Y(n66765) );
  NAND2X1 U70300 ( .A(n66762), .B(n66765), .Y(n66767) );
  NAND2X1 U70301 ( .A(n43491), .B(n43920), .Y(n67079) );
  NAND2X1 U70302 ( .A(n66767), .B(n66770), .Y(n66763) );
  OR2X1 U70303 ( .A(n67121), .B(n66763), .Y(n66776) );
  NOR2X1 U70304 ( .A(n67379), .B(n66776), .Y(n66774) );
  NAND2X1 U70305 ( .A(n66766), .B(n67118), .Y(n67072) );
  NOR2X1 U70306 ( .A(n39557), .B(n67379), .Y(n66769) );
  NAND2X1 U70307 ( .A(n66768), .B(n66767), .Y(n67073) );
  NAND2X1 U70308 ( .A(n66769), .B(n41227), .Y(n66772) );
  NAND2X1 U70309 ( .A(n39557), .B(n66770), .Y(n66775) );
  OR2X1 U70310 ( .A(n67379), .B(n66775), .Y(n66771) );
  NAND2X1 U70311 ( .A(n66772), .B(n66771), .Y(n66773) );
  NOR2X1 U70312 ( .A(n66774), .B(n66773), .Y(n66782) );
  NAND2X1 U70313 ( .A(n66775), .B(n67379), .Y(n66778) );
  INVX1 U70314 ( .A(n66776), .Y(n66777) );
  NOR2X1 U70315 ( .A(n66778), .B(n66777), .Y(n66780) );
  NAND2X1 U70316 ( .A(n41227), .B(n67072), .Y(n66779) );
  NAND2X1 U70317 ( .A(n66780), .B(n66779), .Y(n66781) );
  NAND2X1 U70318 ( .A(n66782), .B(n66781), .Y(n67052) );
  XNOR2X1 U70319 ( .A(n67054), .B(n67052), .Y(n66783) );
  XOR2X1 U70320 ( .A(n67076), .B(n66783), .Y(n67134) );
  XNOR2X1 U70321 ( .A(n66786), .B(n40994), .Y(n67066) );
  NAND2X1 U70322 ( .A(n39968), .B(n67066), .Y(n66787) );
  INVX1 U70323 ( .A(n67066), .Y(n66789) );
  INVX1 U70324 ( .A(n67053), .Y(n67136) );
  XNOR2X1 U70325 ( .A(n67134), .B(n67136), .Y(n67047) );
  NAND2X1 U70326 ( .A(n43942), .B(n43477), .Y(n67147) );
  NAND2X1 U70327 ( .A(n43933), .B(n43483), .Y(n67046) );
  INVX1 U70328 ( .A(n67046), .Y(n67135) );
  XNOR2X1 U70329 ( .A(n67147), .B(n67135), .Y(n66790) );
  XNOR2X1 U70330 ( .A(n67047), .B(n66790), .Y(n66791) );
  XNOR2X1 U70331 ( .A(n41203), .B(n66791), .Y(n67028) );
  NAND2X1 U70332 ( .A(n67344), .B(n66792), .Y(n67146) );
  NAND2X1 U70333 ( .A(n67345), .B(n66793), .Y(n66794) );
  NAND2X1 U70334 ( .A(n67146), .B(n66794), .Y(n67139) );
  XNOR2X1 U70335 ( .A(n67028), .B(n66795), .Y(n66796) );
  XNOR2X1 U70336 ( .A(n66797), .B(n66796), .Y(n67018) );
  INVX1 U70337 ( .A(n67018), .Y(n67333) );
  XNOR2X1 U70338 ( .A(n67333), .B(n67329), .Y(n66804) );
  NAND2X1 U70339 ( .A(n41407), .B(n66799), .Y(n67019) );
  INVX1 U70340 ( .A(n67019), .Y(n66802) );
  INVX1 U70341 ( .A(n66798), .Y(n66800) );
  NAND2X1 U70342 ( .A(n66800), .B(n41407), .Y(n67021) );
  NAND2X1 U70343 ( .A(n67020), .B(n67021), .Y(n66801) );
  NOR2X1 U70344 ( .A(n66802), .B(n66801), .Y(n66803) );
  XNOR2X1 U70345 ( .A(n66804), .B(n66803), .Y(n67494) );
  INVX1 U70346 ( .A(n67494), .Y(n67491) );
  XNOR2X1 U70347 ( .A(n67493), .B(n67491), .Y(n66814) );
  NOR2X1 U70348 ( .A(n66805), .B(n66815), .Y(n66810) );
  NOR2X1 U70349 ( .A(n41205), .B(n41209), .Y(n66807) );
  NAND2X1 U70350 ( .A(n66807), .B(n66806), .Y(n66811) );
  INVX1 U70351 ( .A(n66811), .Y(n66808) );
  NOR2X1 U70352 ( .A(n66808), .B(n66815), .Y(n66809) );
  NOR2X1 U70353 ( .A(n66810), .B(n66809), .Y(n66813) );
  NAND2X1 U70354 ( .A(n66811), .B(n66816), .Y(n66812) );
  NAND2X1 U70355 ( .A(n66813), .B(n66812), .Y(n67495) );
  INVX1 U70356 ( .A(n67495), .Y(n67156) );
  XNOR2X1 U70357 ( .A(n66814), .B(n67156), .Y(n67017) );
  NAND2X1 U70358 ( .A(n42661), .B(n44000), .Y(n67014) );
  NOR2X1 U70359 ( .A(n66829), .B(n66818), .Y(n66828) );
  NOR2X1 U70360 ( .A(n36769), .B(n66819), .Y(n66824) );
  INVX1 U70361 ( .A(n66819), .Y(n66821) );
  NAND2X1 U70362 ( .A(n66821), .B(n66820), .Y(n66823) );
  NOR2X1 U70363 ( .A(n36670), .B(n36671), .Y(n66826) );
  NOR2X1 U70364 ( .A(n66826), .B(n66825), .Y(n66827) );
  INVX1 U70365 ( .A(n66829), .Y(n66830) );
  NAND2X1 U70366 ( .A(n66832), .B(n66834), .Y(n67002) );
  INVX1 U70367 ( .A(n66833), .Y(n66845) );
  NAND2X1 U70368 ( .A(n66845), .B(n66834), .Y(n67003) );
  INVX1 U70369 ( .A(n67003), .Y(n67167) );
  NOR2X1 U70370 ( .A(n66836), .B(n66835), .Y(n66838) );
  NOR2X1 U70371 ( .A(n66836), .B(n66839), .Y(n66837) );
  NOR2X1 U70372 ( .A(n66838), .B(n66837), .Y(n66843) );
  INVX1 U70373 ( .A(n66839), .Y(n66841) );
  NAND2X1 U70374 ( .A(n66841), .B(n66840), .Y(n66842) );
  NAND2X1 U70375 ( .A(n66843), .B(n66842), .Y(n66844) );
  NAND2X1 U70376 ( .A(n66845), .B(n66844), .Y(n67168) );
  NAND2X1 U70377 ( .A(n43799), .B(n44008), .Y(n67507) );
  NAND2X1 U70378 ( .A(n43772), .B(n44017), .Y(n67008) );
  XNOR2X1 U70379 ( .A(n67507), .B(n67008), .Y(n66846) );
  XNOR2X1 U70380 ( .A(n66996), .B(n41633), .Y(n66995) );
  NAND2X1 U70381 ( .A(n43788), .B(n44055), .Y(n66966) );
  NAND2X1 U70382 ( .A(n43725), .B(n44048), .Y(n66983) );
  XNOR2X1 U70383 ( .A(n66966), .B(n66983), .Y(n66847) );
  NAND2X1 U70384 ( .A(n43613), .B(n40487), .Y(n72182) );
  XNOR2X1 U70385 ( .A(n66972), .B(n66850), .Y(n66855) );
  NAND2X1 U70386 ( .A(n66852), .B(n66851), .Y(n66853) );
  NOR2X1 U70387 ( .A(n38368), .B(n66853), .Y(n66854) );
  XNOR2X1 U70388 ( .A(n66855), .B(n66854), .Y(n67545) );
  INVX1 U70389 ( .A(n66878), .Y(n66857) );
  NOR2X1 U70390 ( .A(n66879), .B(n66868), .Y(n66856) );
  NOR2X1 U70391 ( .A(n66857), .B(n66856), .Y(n66872) );
  NOR2X1 U70392 ( .A(n41291), .B(n66858), .Y(n66860) );
  NOR2X1 U70393 ( .A(n66860), .B(n66859), .Y(n66864) );
  NAND2X1 U70394 ( .A(n66862), .B(n66861), .Y(n66863) );
  NOR2X1 U70395 ( .A(n66864), .B(n66863), .Y(n66867) );
  NOR2X1 U70396 ( .A(n41324), .B(n39171), .Y(n66866) );
  NOR2X1 U70397 ( .A(n66867), .B(n66866), .Y(n66870) );
  NAND2X1 U70398 ( .A(n66879), .B(n66868), .Y(n66869) );
  NAND2X1 U70399 ( .A(n66870), .B(n66869), .Y(n66871) );
  INVX1 U70400 ( .A(n66946), .Y(n66882) );
  NOR2X1 U70401 ( .A(n44052), .B(n66878), .Y(n66877) );
  NOR2X1 U70402 ( .A(n39948), .B(n39309), .Y(n66875) );
  NAND2X1 U70403 ( .A(n66875), .B(n66495), .Y(n66876) );
  NOR2X1 U70404 ( .A(n66879), .B(n66878), .Y(n66881) );
  NOR2X1 U70405 ( .A(n66882), .B(n67548), .Y(n66883) );
  XNOR2X1 U70406 ( .A(n66883), .B(n66884), .Y(n67653) );
  XNOR2X1 U70407 ( .A(n43542), .B(n67653), .Y(n66885) );
  XOR2X1 U70408 ( .A(n66939), .B(n66885), .Y(n67199) );
  XNOR2X1 U70409 ( .A(n66886), .B(n67199), .Y(n66936) );
  XNOR2X1 U70410 ( .A(n66888), .B(n66887), .Y(n67208) );
  NOR2X1 U70411 ( .A(n67208), .B(n43552), .Y(n66889) );
  NOR2X1 U70412 ( .A(n37362), .B(n66889), .Y(n66892) );
  NAND2X1 U70413 ( .A(n67203), .B(n66890), .Y(n66891) );
  XNOR2X1 U70414 ( .A(n40414), .B(n41368), .Y(n67221) );
  XNOR2X1 U70415 ( .A(n70762), .B(n67221), .Y(n66893) );
  XNOR2X1 U70416 ( .A(n66929), .B(n43654), .Y(n66894) );
  XNOR2X1 U70417 ( .A(n43524), .B(n36381), .Y(n67232) );
  NOR2X1 U70418 ( .A(n41106), .B(n66895), .Y(n66898) );
  NOR2X1 U70419 ( .A(n43523), .B(n40969), .Y(n66897) );
  INVX1 U70420 ( .A(n66899), .Y(n66900) );
  NAND2X1 U70421 ( .A(n43522), .B(n40969), .Y(n67260) );
  NAND2X1 U70422 ( .A(n67260), .B(n36488), .Y(n67231) );
  XNOR2X1 U70423 ( .A(n67231), .B(n43679), .Y(n66901) );
  XNOR2X1 U70424 ( .A(n66901), .B(n67232), .Y(n66902) );
  XNOR2X1 U70425 ( .A(n43512), .B(n66922), .Y(n66903) );
  XNOR2X1 U70426 ( .A(n66904), .B(n66903), .Y(n66918) );
  XNOR2X1 U70427 ( .A(n36362), .B(n43693), .Y(n66905) );
  XNOR2X1 U70428 ( .A(n66917), .B(n43708), .Y(n66906) );
  XNOR2X1 U70429 ( .A(n66907), .B(n66906), .Y(n66912) );
  XNOR2X1 U70430 ( .A(n66909), .B(n66908), .Y(n66910) );
  XNOR2X1 U70431 ( .A(n66910), .B(n41988), .Y(n66911) );
  MX2X1 U70432 ( .A(n66912), .B(n66911), .S0(n43719), .Y(u_muldiv_result_r[14]) );
  NAND2X1 U70433 ( .A(u_muldiv_mult_result_q[14]), .B(n44632), .Y(n14008) );
  NAND2X1 U70434 ( .A(n66913), .B(n39519), .Y(n66915) );
  OR2X1 U70435 ( .A(n37922), .B(n43715), .Y(n66914) );
  NAND2X1 U70436 ( .A(n36362), .B(n43698), .Y(n66920) );
  NAND2X1 U70437 ( .A(n66920), .B(n66919), .Y(n67608) );
  NAND2X1 U70438 ( .A(n67607), .B(n67608), .Y(n67595) );
  INVX1 U70439 ( .A(n66921), .Y(n66924) );
  NOR2X1 U70440 ( .A(n66924), .B(n66923), .Y(n66925) );
  NAND2X1 U70441 ( .A(n39518), .B(n67591), .Y(n67237) );
  XNOR2X1 U70442 ( .A(n38047), .B(n41096), .Y(n67230) );
  INVX1 U70443 ( .A(n66929), .Y(n66927) );
  NAND2X1 U70444 ( .A(n43655), .B(n66927), .Y(n67581) );
  NAND2X1 U70445 ( .A(n66928), .B(n67581), .Y(n66930) );
  NAND2X1 U70446 ( .A(n66929), .B(n43660), .Y(n67583) );
  NAND2X1 U70447 ( .A(n66930), .B(n67583), .Y(n67256) );
  XNOR2X1 U70448 ( .A(n43667), .B(n40414), .Y(n66933) );
  XNOR2X1 U70449 ( .A(n66933), .B(n41368), .Y(n66934) );
  NAND2X1 U70450 ( .A(n43620), .B(n66938), .Y(n67283) );
  NAND2X1 U70451 ( .A(n67282), .B(n67862), .Y(n67576) );
  INVX1 U70452 ( .A(n39797), .Y(n67658) );
  INVX1 U70453 ( .A(n67567), .Y(n66940) );
  NAND2X1 U70454 ( .A(n43536), .B(n66940), .Y(n66941) );
  NOR2X1 U70455 ( .A(n67565), .B(n66941), .Y(n66945) );
  INVX1 U70456 ( .A(n67565), .Y(n66943) );
  NAND2X1 U70457 ( .A(n67658), .B(n43541), .Y(n66942) );
  NOR2X1 U70458 ( .A(n66943), .B(n66942), .Y(n66944) );
  NOR2X1 U70459 ( .A(n66945), .B(n66944), .Y(n67197) );
  NAND2X1 U70460 ( .A(n41319), .B(n43587), .Y(n67549) );
  INVX1 U70461 ( .A(n66949), .Y(n66959) );
  NAND2X1 U70462 ( .A(n66951), .B(n66950), .Y(n66957) );
  NAND2X1 U70463 ( .A(n66953), .B(n66952), .Y(n66955) );
  NAND2X1 U70464 ( .A(n66955), .B(n66954), .Y(n66956) );
  NOR2X1 U70465 ( .A(n66957), .B(n66956), .Y(n66958) );
  NOR2X1 U70466 ( .A(n66959), .B(n66958), .Y(n66962) );
  INVX1 U70467 ( .A(n66983), .Y(n66991) );
  XNOR2X1 U70468 ( .A(n66991), .B(n66996), .Y(n66960) );
  XNOR2X1 U70469 ( .A(n66960), .B(n41633), .Y(n66961) );
  XNOR2X1 U70470 ( .A(n66962), .B(n66961), .Y(n66973) );
  NOR2X1 U70471 ( .A(n39310), .B(n66966), .Y(n66965) );
  NAND2X1 U70472 ( .A(n66965), .B(n66964), .Y(n67536) );
  INVX1 U70473 ( .A(n66966), .Y(n66974) );
  NOR2X1 U70474 ( .A(n39929), .B(n39300), .Y(n66970) );
  NAND2X1 U70475 ( .A(n66968), .B(n66967), .Y(n66969) );
  NAND2X1 U70476 ( .A(n66970), .B(n66969), .Y(n66971) );
  NAND2X1 U70477 ( .A(n66974), .B(n66973), .Y(n67537) );
  NAND2X1 U70478 ( .A(n66975), .B(n67537), .Y(n66976) );
  NOR2X1 U70479 ( .A(n39633), .B(n66976), .Y(n67178) );
  NOR2X1 U70480 ( .A(n66977), .B(n36627), .Y(n66979) );
  NOR2X1 U70481 ( .A(n66979), .B(n66978), .Y(n66980) );
  NOR2X1 U70482 ( .A(n39924), .B(n66980), .Y(n66982) );
  NAND2X1 U70483 ( .A(n66991), .B(n44025), .Y(n66981) );
  NOR2X1 U70484 ( .A(n66982), .B(n66981), .Y(n66989) );
  NOR2X1 U70485 ( .A(n66986), .B(n66983), .Y(n66985) );
  NOR2X1 U70486 ( .A(n44029), .B(n66986), .Y(n66987) );
  NAND2X1 U70487 ( .A(n66993), .B(n66992), .Y(n66994) );
  NOR2X1 U70488 ( .A(n66996), .B(n67521), .Y(n66998) );
  XNOR2X1 U70489 ( .A(n39535), .B(n66997), .Y(n67522) );
  NOR2X1 U70490 ( .A(n66998), .B(n67524), .Y(n67000) );
  INVX1 U70491 ( .A(n67522), .Y(n67519) );
  NAND2X1 U70492 ( .A(n67519), .B(n67523), .Y(n66999) );
  INVX1 U70493 ( .A(n67507), .Y(n67001) );
  XNOR2X1 U70494 ( .A(n67508), .B(n67001), .Y(n67007) );
  INVX1 U70495 ( .A(n67168), .Y(n67005) );
  NAND2X1 U70496 ( .A(n67003), .B(n67002), .Y(n67004) );
  NOR2X1 U70497 ( .A(n67005), .B(n67004), .Y(n67006) );
  XNOR2X1 U70498 ( .A(n67007), .B(n67006), .Y(n67310) );
  INVX1 U70499 ( .A(n67310), .Y(n67307) );
  NOR2X1 U70500 ( .A(n67307), .B(n67008), .Y(n67010) );
  NOR2X1 U70501 ( .A(n39535), .B(n67008), .Y(n67009) );
  NOR2X1 U70502 ( .A(n67010), .B(n67009), .Y(n67013) );
  NAND2X1 U70503 ( .A(n67310), .B(n67011), .Y(n67012) );
  NAND2X1 U70504 ( .A(n67013), .B(n67012), .Y(n67315) );
  INVX1 U70505 ( .A(n67014), .Y(n67015) );
  INVX1 U70506 ( .A(n67814), .Y(n67514) );
  NAND2X1 U70507 ( .A(n42661), .B(n44008), .Y(n67817) );
  INVX1 U70508 ( .A(n67817), .Y(n67321) );
  NAND2X1 U70509 ( .A(n43799), .B(n44017), .Y(n67829) );
  INVX1 U70510 ( .A(n67829), .Y(n67515) );
  XNOR2X1 U70511 ( .A(n67321), .B(n67515), .Y(n67313) );
  NAND2X1 U70512 ( .A(n42711), .B(n44000), .Y(n67502) );
  NAND2X1 U70513 ( .A(n38603), .B(n67018), .Y(n67332) );
  NAND2X1 U70514 ( .A(n67022), .B(n67328), .Y(n67023) );
  NAND2X1 U70515 ( .A(n67332), .B(n67023), .Y(n67323) );
  NAND2X1 U70516 ( .A(n67025), .B(n67024), .Y(n67027) );
  NAND2X1 U70517 ( .A(n67027), .B(n67026), .Y(n67466) );
  INVX1 U70518 ( .A(n67139), .Y(n67357) );
  NAND2X1 U70519 ( .A(n67684), .B(n67465), .Y(n67155) );
  INVX1 U70520 ( .A(n67047), .Y(n67034) );
  NAND2X1 U70521 ( .A(n67034), .B(n67031), .Y(n67032) );
  NOR2X1 U70522 ( .A(n67033), .B(n67032), .Y(n67038) );
  NOR2X1 U70523 ( .A(n67135), .B(n67034), .Y(n67036) );
  NOR2X1 U70524 ( .A(n67036), .B(n67035), .Y(n67037) );
  NOR2X1 U70525 ( .A(n67038), .B(n67037), .Y(n67051) );
  NAND2X1 U70526 ( .A(n67040), .B(n67039), .Y(n67041) );
  NOR2X1 U70527 ( .A(n67042), .B(n67041), .Y(n67045) );
  NAND2X1 U70528 ( .A(n67135), .B(n67043), .Y(n67044) );
  NOR2X1 U70529 ( .A(n67045), .B(n67044), .Y(n67049) );
  NOR2X1 U70530 ( .A(n67047), .B(n67046), .Y(n67048) );
  NOR2X1 U70531 ( .A(n67049), .B(n67048), .Y(n67050) );
  NAND2X1 U70532 ( .A(n67051), .B(n67050), .Y(n67371) );
  XNOR2X1 U70533 ( .A(n41719), .B(n41718), .Y(n67132) );
  NAND2X1 U70534 ( .A(n67055), .B(n67053), .Y(n67459) );
  NOR2X1 U70535 ( .A(n37369), .B(n67055), .Y(n67071) );
  INVX1 U70536 ( .A(n67056), .Y(n67061) );
  INVX1 U70537 ( .A(n67057), .Y(n67059) );
  NAND2X1 U70538 ( .A(n67059), .B(n67058), .Y(n67060) );
  NOR2X1 U70539 ( .A(n67061), .B(n67060), .Y(n67065) );
  NAND2X1 U70540 ( .A(n67063), .B(n67062), .Y(n67064) );
  NOR2X1 U70541 ( .A(n67065), .B(n67064), .Y(n67067) );
  NAND2X1 U70542 ( .A(n67067), .B(n67066), .Y(n67068) );
  NAND2X1 U70543 ( .A(n67069), .B(n67068), .Y(n67070) );
  NAND2X1 U70544 ( .A(n67073), .B(n67072), .Y(n67376) );
  XNOR2X1 U70545 ( .A(n41711), .B(n41248), .Y(n67074) );
  XNOR2X1 U70546 ( .A(n67074), .B(n41240), .Y(n67075) );
  NAND2X1 U70547 ( .A(n67442), .B(n67076), .Y(n67436) );
  OR2X1 U70548 ( .A(n67442), .B(n67077), .Y(n67078) );
  NOR2X1 U70549 ( .A(n67441), .B(n67078), .Y(n67080) );
  NOR2X1 U70550 ( .A(n67080), .B(n67079), .Y(n67445) );
  NOR2X1 U70551 ( .A(n67441), .B(n67442), .Y(n67081) );
  NAND2X1 U70552 ( .A(n67081), .B(n40994), .Y(n67082) );
  NAND2X1 U70553 ( .A(n67445), .B(n67082), .Y(n67437) );
  NAND2X1 U70554 ( .A(n67436), .B(n67437), .Y(n67439) );
  NAND2X1 U70555 ( .A(n43896), .B(n43607), .Y(n67415) );
  NAND2X1 U70556 ( .A(n41509), .B(n43604), .Y(n72383) );
  XNOR2X1 U70557 ( .A(n72383), .B(n67083), .Y(n67087) );
  NAND2X1 U70558 ( .A(n67084), .B(n72365), .Y(n67085) );
  NAND2X1 U70559 ( .A(n71843), .B(n67085), .Y(n72373) );
  NAND2X1 U70560 ( .A(n72373), .B(n67426), .Y(n67086) );
  NAND2X1 U70561 ( .A(n72370), .B(n67086), .Y(n72382) );
  INVX1 U70562 ( .A(n72382), .Y(n72386) );
  XNOR2X1 U70563 ( .A(n67087), .B(n72386), .Y(n68107) );
  INVX1 U70564 ( .A(n68107), .Y(n67752) );
  NAND2X1 U70565 ( .A(n67746), .B(n67088), .Y(n67089) );
  NAND2X1 U70566 ( .A(n41509), .B(n67089), .Y(n67416) );
  NAND2X1 U70567 ( .A(n43903), .B(n43518), .Y(n67761) );
  INVX1 U70568 ( .A(n67761), .Y(n67760) );
  XNOR2X1 U70569 ( .A(n67762), .B(n67760), .Y(n67101) );
  INVX1 U70570 ( .A(n67094), .Y(n67099) );
  NOR2X1 U70571 ( .A(n67090), .B(n67099), .Y(n67092) );
  NAND2X1 U70572 ( .A(n67092), .B(n67091), .Y(n67093) );
  NAND2X1 U70573 ( .A(n41708), .B(n67093), .Y(n67407) );
  NAND2X1 U70574 ( .A(n67095), .B(n67094), .Y(n67405) );
  INVX1 U70575 ( .A(n67405), .Y(n67097) );
  NAND2X1 U70576 ( .A(n67099), .B(n67098), .Y(n67410) );
  NAND2X1 U70577 ( .A(n67100), .B(n67410), .Y(n68113) );
  NAND2X1 U70578 ( .A(n43909), .B(n43501), .Y(n67738) );
  INVX1 U70579 ( .A(n67738), .Y(n67393) );
  XNOR2X1 U70580 ( .A(n67402), .B(n67393), .Y(n67117) );
  INVX1 U70581 ( .A(n67102), .Y(n67389) );
  NOR2X1 U70582 ( .A(n67389), .B(n67385), .Y(n67103) );
  NOR2X1 U70583 ( .A(n67103), .B(n67395), .Y(n67105) );
  NAND2X1 U70584 ( .A(n67110), .B(n67109), .Y(n67387) );
  NOR2X1 U70585 ( .A(n67395), .B(n67387), .Y(n67104) );
  NOR2X1 U70586 ( .A(n67105), .B(n67104), .Y(n67116) );
  NOR2X1 U70587 ( .A(n67106), .B(n67385), .Y(n67107) );
  NOR2X1 U70588 ( .A(n67107), .B(n67384), .Y(n67114) );
  NOR2X1 U70589 ( .A(n67109), .B(n67108), .Y(n67112) );
  NAND2X1 U70590 ( .A(n67110), .B(n67385), .Y(n67111) );
  NOR2X1 U70591 ( .A(n67112), .B(n67111), .Y(n67113) );
  NOR2X1 U70592 ( .A(n67114), .B(n67113), .Y(n67115) );
  NAND2X1 U70593 ( .A(n67116), .B(n67115), .Y(n67403) );
  INVX1 U70594 ( .A(n67403), .Y(n67735) );
  XNOR2X1 U70595 ( .A(n67117), .B(n67735), .Y(n67772) );
  NAND2X1 U70596 ( .A(n43918), .B(n43496), .Y(n67771) );
  INVX1 U70597 ( .A(n67771), .Y(n67377) );
  XNOR2X1 U70598 ( .A(n67772), .B(n67377), .Y(n67129) );
  INVX1 U70599 ( .A(n67379), .Y(n67124) );
  NAND2X1 U70600 ( .A(n67124), .B(n67376), .Y(n67128) );
  INVX1 U70601 ( .A(n67118), .Y(n67119) );
  NOR2X1 U70602 ( .A(n67119), .B(n67121), .Y(n67120) );
  NOR2X1 U70603 ( .A(n39557), .B(n67120), .Y(n67126) );
  NOR2X1 U70604 ( .A(n67122), .B(n67121), .Y(n67123) );
  NOR2X1 U70605 ( .A(n67124), .B(n67123), .Y(n67125) );
  NAND2X1 U70606 ( .A(n67126), .B(n67125), .Y(n67127) );
  NAND2X1 U70607 ( .A(n41711), .B(n67127), .Y(n67375) );
  NAND2X1 U70608 ( .A(n67128), .B(n67375), .Y(n67773) );
  XNOR2X1 U70609 ( .A(n67129), .B(n38168), .Y(n67440) );
  NAND2X1 U70610 ( .A(n43491), .B(n43929), .Y(n67724) );
  INVX1 U70611 ( .A(n67724), .Y(n67448) );
  XNOR2X1 U70612 ( .A(n67440), .B(n67448), .Y(n67130) );
  XNOR2X1 U70613 ( .A(n38736), .B(n67130), .Y(n67715) );
  NAND2X1 U70614 ( .A(n43933), .B(n43487), .Y(n67455) );
  XNOR2X1 U70615 ( .A(n67715), .B(n67455), .Y(n67131) );
  XNOR2X1 U70616 ( .A(n67714), .B(n67131), .Y(n67370) );
  INVX1 U70617 ( .A(n67370), .Y(n67372) );
  XNOR2X1 U70618 ( .A(n67132), .B(n67372), .Y(n67133) );
  XNOR2X1 U70619 ( .A(n67371), .B(n67133), .Y(n67152) );
  XNOR2X1 U70620 ( .A(n67135), .B(n67134), .Y(n67137) );
  XNOR2X1 U70621 ( .A(n67137), .B(n67136), .Y(n67138) );
  XNOR2X1 U70622 ( .A(n41203), .B(n67138), .Y(n67358) );
  NOR2X1 U70623 ( .A(n67344), .B(n67339), .Y(n67145) );
  NAND2X1 U70624 ( .A(n67141), .B(n67140), .Y(n67142) );
  NAND2X1 U70625 ( .A(n67142), .B(n40247), .Y(n67143) );
  NOR2X1 U70626 ( .A(n67344), .B(n67143), .Y(n67144) );
  INVX1 U70627 ( .A(n67146), .Y(n67349) );
  INVX1 U70628 ( .A(n67147), .Y(n67359) );
  NOR2X1 U70629 ( .A(n67363), .B(n40140), .Y(n67149) );
  NAND2X1 U70630 ( .A(n67359), .B(n67358), .Y(n67148) );
  NAND2X1 U70631 ( .A(n67149), .B(n67148), .Y(n67150) );
  NOR2X1 U70632 ( .A(n39979), .B(n67150), .Y(n67151) );
  XNOR2X1 U70633 ( .A(n67152), .B(n67151), .Y(n67682) );
  NAND2X1 U70634 ( .A(n43795), .B(n43992), .Y(n67322) );
  NAND2X1 U70635 ( .A(n43982), .B(n43774), .Y(n67689) );
  XNOR2X1 U70636 ( .A(n67322), .B(n67689), .Y(n67153) );
  XNOR2X1 U70637 ( .A(n67682), .B(n67153), .Y(n67154) );
  INVX1 U70638 ( .A(n67503), .Y(n67499) );
  XNOR2X1 U70639 ( .A(n67502), .B(n67499), .Y(n67162) );
  NOR2X1 U70640 ( .A(n67494), .B(n67156), .Y(n67160) );
  INVX1 U70641 ( .A(n67493), .Y(n67492) );
  NAND2X1 U70642 ( .A(n67492), .B(n67491), .Y(n67158) );
  NAND2X1 U70643 ( .A(n67492), .B(n67495), .Y(n67157) );
  NAND2X1 U70644 ( .A(n67158), .B(n67157), .Y(n67159) );
  NOR2X1 U70645 ( .A(n67160), .B(n67159), .Y(n67161) );
  XNOR2X1 U70646 ( .A(n67162), .B(n67161), .Y(n67813) );
  INVX1 U70647 ( .A(n67813), .Y(n67512) );
  XNOR2X1 U70648 ( .A(n67163), .B(n67512), .Y(n67164) );
  XNOR2X1 U70649 ( .A(n67514), .B(n67164), .Y(n67172) );
  NOR2X1 U70650 ( .A(n40128), .B(n67507), .Y(n67166) );
  NOR2X1 U70651 ( .A(n67508), .B(n67507), .Y(n67165) );
  NOR2X1 U70652 ( .A(n67166), .B(n67165), .Y(n67170) );
  NOR2X1 U70653 ( .A(n38139), .B(n67167), .Y(n67169) );
  NAND2X1 U70654 ( .A(n67170), .B(n67510), .Y(n67833) );
  INVX1 U70655 ( .A(n40307), .Y(n67171) );
  XNOR2X1 U70656 ( .A(n67172), .B(n67171), .Y(n67173) );
  NAND2X1 U70657 ( .A(n43725), .B(n44055), .Y(n67299) );
  NAND2X1 U70658 ( .A(n42632), .B(n44048), .Y(n67527) );
  INVX1 U70659 ( .A(n67527), .Y(n67532) );
  XNOR2X1 U70660 ( .A(n67299), .B(n67532), .Y(n67174) );
  XNOR2X1 U70661 ( .A(n67531), .B(n67174), .Y(n67175) );
  XNOR2X1 U70662 ( .A(n41119), .B(n67175), .Y(n67540) );
  NAND2X1 U70663 ( .A(n43613), .B(n43788), .Y(n72168) );
  XNOR2X1 U70664 ( .A(n67540), .B(n43569), .Y(n67176) );
  XNOR2X1 U70665 ( .A(n67303), .B(n67176), .Y(n67177) );
  XNOR2X1 U70666 ( .A(n67178), .B(n67177), .Y(n67554) );
  INVX1 U70667 ( .A(n67655), .Y(n67661) );
  NOR2X1 U70668 ( .A(n38209), .B(n67180), .Y(n67181) );
  NOR2X1 U70669 ( .A(n67182), .B(n67181), .Y(n67184) );
  NOR2X1 U70670 ( .A(n67184), .B(n67183), .Y(n67190) );
  NAND2X1 U70671 ( .A(n67186), .B(n67185), .Y(n67188) );
  NAND2X1 U70672 ( .A(n67188), .B(n67187), .Y(n67189) );
  NAND2X1 U70673 ( .A(n67192), .B(n43572), .Y(n67555) );
  NOR2X1 U70674 ( .A(n67657), .B(n67193), .Y(n67195) );
  XNOR2X1 U70675 ( .A(n67647), .B(n43565), .Y(n67196) );
  XNOR2X1 U70676 ( .A(n67197), .B(n67196), .Y(n67287) );
  XNOR2X1 U70677 ( .A(n67287), .B(n43621), .Y(n67202) );
  NAND2X1 U70678 ( .A(n67200), .B(n43559), .Y(n67294) );
  NOR2X1 U70679 ( .A(n67200), .B(n43560), .Y(n67201) );
  OR2X1 U70680 ( .A(n67201), .B(n66937), .Y(n67291) );
  XNOR2X1 U70681 ( .A(n67202), .B(n40953), .Y(n67575) );
  INVX1 U70682 ( .A(n67203), .Y(n67205) );
  NOR2X1 U70683 ( .A(n67205), .B(n67204), .Y(n67206) );
  NOR2X1 U70684 ( .A(n43545), .B(n67206), .Y(n67207) );
  NOR2X1 U70685 ( .A(n67208), .B(n43551), .Y(n67211) );
  NOR2X1 U70686 ( .A(n40492), .B(n43553), .Y(n67210) );
  NOR2X1 U70687 ( .A(n67211), .B(n67210), .Y(n67215) );
  XNOR2X1 U70688 ( .A(n67640), .B(n43633), .Y(n67216) );
  NAND2X1 U70689 ( .A(n67219), .B(n43636), .Y(n67278) );
  INVX1 U70690 ( .A(n67278), .Y(n67874) );
  NAND2X1 U70691 ( .A(n67872), .B(n67220), .Y(n67279) );
  INVX1 U70692 ( .A(n67632), .Y(n67272) );
  INVX1 U70693 ( .A(n70762), .Y(n72088) );
  XNOR2X1 U70694 ( .A(n67272), .B(n72088), .Y(n67227) );
  NAND2X1 U70695 ( .A(n67221), .B(n43671), .Y(n67274) );
  NAND2X1 U70696 ( .A(n43664), .B(n36425), .Y(n67631) );
  NAND2X1 U70697 ( .A(n67223), .B(n67222), .Y(n67225) );
  NAND2X1 U70698 ( .A(n67225), .B(n67224), .Y(n67226) );
  NAND2X1 U70699 ( .A(n67631), .B(n67226), .Y(n67275) );
  XNOR2X1 U70700 ( .A(n67227), .B(n41064), .Y(n67228) );
  XNOR2X1 U70701 ( .A(n43655), .B(n36472), .Y(n67255) );
  XNOR2X1 U70702 ( .A(n43528), .B(n67255), .Y(n67229) );
  XOR2X1 U70703 ( .A(n67256), .B(n67229), .Y(n67246) );
  XNOR2X1 U70704 ( .A(n67230), .B(n67246), .Y(n67235) );
  XNOR2X1 U70705 ( .A(n67235), .B(n67234), .Y(n67590) );
  XNOR2X1 U70706 ( .A(n43512), .B(n67590), .Y(n67236) );
  XNOR2X1 U70707 ( .A(n67237), .B(n67236), .Y(n67606) );
  XNOR2X1 U70708 ( .A(n67244), .B(n43708), .Y(n67238) );
  XNOR2X1 U70709 ( .A(n37907), .B(n67238), .Y(n67243) );
  XNOR2X1 U70710 ( .A(n67240), .B(n67239), .Y(n67241) );
  XNOR2X1 U70711 ( .A(n42001), .B(n67241), .Y(n67242) );
  MX2X1 U70712 ( .A(n67243), .B(n67242), .S0(n43719), .Y(u_muldiv_result_r[15]) );
  NAND2X1 U70713 ( .A(u_muldiv_mult_result_q[15]), .B(n44632), .Y(n13997) );
  NAND2X1 U70714 ( .A(n37909), .B(n43712), .Y(n67245) );
  XNOR2X1 U70715 ( .A(n41096), .B(n67246), .Y(n67251) );
  NAND2X1 U70716 ( .A(n67251), .B(n43682), .Y(n67893) );
  NOR2X1 U70717 ( .A(n43678), .B(n67247), .Y(n67250) );
  INVX1 U70718 ( .A(n67251), .Y(n67252) );
  NAND2X1 U70719 ( .A(n43677), .B(n67252), .Y(n67253) );
  NAND2X1 U70720 ( .A(n67253), .B(n67254), .Y(n67892) );
  INVX1 U70721 ( .A(n67264), .Y(n67257) );
  NAND2X1 U70722 ( .A(n67257), .B(n43528), .Y(n67616) );
  NOR2X1 U70723 ( .A(n38003), .B(n67259), .Y(n67263) );
  NAND2X1 U70724 ( .A(n67261), .B(n67260), .Y(n67262) );
  XNOR2X1 U70725 ( .A(n38047), .B(n41059), .Y(n67588) );
  XNOR2X1 U70726 ( .A(n43666), .B(n41300), .Y(n67265) );
  XNOR2X1 U70727 ( .A(n67265), .B(n40504), .Y(n67266) );
  XNOR2X1 U70728 ( .A(n41064), .B(n67266), .Y(n67269) );
  INVX1 U70729 ( .A(n67269), .Y(n67267) );
  NOR2X1 U70730 ( .A(n67268), .B(n41316), .Y(n67271) );
  NAND2X1 U70731 ( .A(n67269), .B(n43648), .Y(n67270) );
  NAND2X1 U70732 ( .A(n43664), .B(n67273), .Y(n67634) );
  NOR2X1 U70733 ( .A(n40504), .B(n43639), .Y(n67281) );
  INVX1 U70734 ( .A(n67640), .Y(n67643) );
  XNOR2X1 U70735 ( .A(n67643), .B(n67276), .Y(n67277) );
  NAND2X1 U70736 ( .A(n43631), .B(n67277), .Y(n67878) );
  INVX1 U70737 ( .A(n67277), .Y(n67875) );
  NAND2X1 U70738 ( .A(n67278), .B(n67279), .Y(n67280) );
  NOR2X1 U70739 ( .A(n36750), .B(n38959), .Y(n67630) );
  NOR2X1 U70740 ( .A(n36647), .B(n67286), .Y(n67289) );
  NAND2X1 U70741 ( .A(n43620), .B(n67290), .Y(n67863) );
  INVX1 U70742 ( .A(n67291), .Y(n67295) );
  INVX1 U70743 ( .A(n67647), .Y(n67646) );
  NOR2X1 U70744 ( .A(n67646), .B(n43560), .Y(n67292) );
  NAND2X1 U70745 ( .A(n67295), .B(n67292), .Y(n67293) );
  NAND2X1 U70746 ( .A(n67294), .B(n43559), .Y(n67297) );
  OR2X1 U70747 ( .A(n67295), .B(n36668), .Y(n67296) );
  XNOR2X1 U70748 ( .A(n43621), .B(n67628), .Y(n67572) );
  XNOR2X1 U70749 ( .A(n67531), .B(n67532), .Y(n67298) );
  XNOR2X1 U70750 ( .A(n41119), .B(n67298), .Y(n67302) );
  NOR2X1 U70751 ( .A(n67302), .B(n67299), .Y(n67301) );
  NOR2X1 U70752 ( .A(n39586), .B(n67299), .Y(n67300) );
  INVX1 U70753 ( .A(n67302), .Y(n67304) );
  NAND2X1 U70754 ( .A(n42632), .B(n44055), .Y(n67665) );
  XNOR2X1 U70755 ( .A(n67665), .B(n43593), .Y(n67534) );
  NOR2X1 U70756 ( .A(n41378), .B(n67307), .Y(n67309) );
  NOR2X1 U70757 ( .A(n44020), .B(n41378), .Y(n67308) );
  NOR2X1 U70758 ( .A(n67309), .B(n67308), .Y(n67312) );
  NAND2X1 U70759 ( .A(n67310), .B(n44017), .Y(n67311) );
  XNOR2X1 U70760 ( .A(n67313), .B(n67512), .Y(n67314) );
  NAND2X1 U70761 ( .A(n42183), .B(n67316), .Y(n67680) );
  INVX1 U70762 ( .A(n67680), .Y(n68039) );
  NOR2X1 U70763 ( .A(n68039), .B(n39543), .Y(n67317) );
  NAND2X1 U70764 ( .A(n67316), .B(n67315), .Y(n67676) );
  NAND2X1 U70765 ( .A(n67512), .B(n67318), .Y(n67812) );
  NOR2X1 U70766 ( .A(n41178), .B(n41146), .Y(n67320) );
  NAND2X1 U70767 ( .A(n67321), .B(n67815), .Y(n67809) );
  NAND2X1 U70768 ( .A(n43799), .B(n44025), .Y(n68284) );
  INVX1 U70769 ( .A(n68284), .Y(n68055) );
  XNOR2X1 U70770 ( .A(n67825), .B(n68055), .Y(n67505) );
  INVX1 U70771 ( .A(n67322), .Y(n67331) );
  NAND2X1 U70772 ( .A(n67331), .B(n67323), .Y(n67793) );
  INVX1 U70773 ( .A(n67689), .Y(n67683) );
  INVX1 U70774 ( .A(n67682), .Y(n67690) );
  XNOR2X1 U70775 ( .A(n67683), .B(n67690), .Y(n67327) );
  NOR2X1 U70776 ( .A(n39971), .B(n41165), .Y(n67324) );
  NAND2X1 U70777 ( .A(n67324), .B(n41155), .Y(n67325) );
  NAND2X1 U70778 ( .A(n67479), .B(n67325), .Y(n67326) );
  NAND2X1 U70779 ( .A(n67326), .B(n67684), .Y(n67473) );
  INVX1 U70780 ( .A(n67328), .Y(n67334) );
  NOR2X1 U70781 ( .A(n67334), .B(n67329), .Y(n67330) );
  NOR2X1 U70782 ( .A(n67331), .B(n67330), .Y(n67336) );
  NAND2X1 U70783 ( .A(n67336), .B(n67335), .Y(n67337) );
  NAND2X1 U70784 ( .A(n67338), .B(n67337), .Y(n67794) );
  NAND2X1 U70785 ( .A(n67793), .B(n67794), .Y(n67789) );
  NOR2X1 U70786 ( .A(n40247), .B(n67341), .Y(n67343) );
  NAND2X1 U70787 ( .A(n41127), .B(n40327), .Y(n67340) );
  NOR2X1 U70788 ( .A(n67341), .B(n67340), .Y(n67342) );
  NOR2X1 U70789 ( .A(n67343), .B(n67342), .Y(n67347) );
  NAND2X1 U70790 ( .A(n67345), .B(n67344), .Y(n67346) );
  NAND2X1 U70791 ( .A(n67347), .B(n67346), .Y(n67348) );
  NOR2X1 U70792 ( .A(n67349), .B(n67348), .Y(n67350) );
  INVX1 U70793 ( .A(n67358), .Y(n67356) );
  NAND2X1 U70794 ( .A(n67350), .B(n67356), .Y(n67351) );
  NAND2X1 U70795 ( .A(n67359), .B(n67351), .Y(n67353) );
  NAND2X1 U70796 ( .A(n67353), .B(n67352), .Y(n67354) );
  NAND2X1 U70797 ( .A(n41718), .B(n67354), .Y(n67369) );
  XNOR2X1 U70798 ( .A(n41719), .B(n40267), .Y(n67355) );
  XNOR2X1 U70799 ( .A(n67355), .B(n67372), .Y(n67367) );
  NOR2X1 U70800 ( .A(n67357), .B(n67356), .Y(n67362) );
  NAND2X1 U70801 ( .A(n67148), .B(n67360), .Y(n67361) );
  NOR2X1 U70802 ( .A(n67362), .B(n67361), .Y(n67365) );
  NOR2X1 U70803 ( .A(n41718), .B(n67363), .Y(n67364) );
  NAND2X1 U70804 ( .A(n67365), .B(n67364), .Y(n67366) );
  NAND2X1 U70805 ( .A(n67367), .B(n67366), .Y(n67368) );
  NAND2X1 U70806 ( .A(n67369), .B(n67368), .Y(n67703) );
  NAND2X1 U70807 ( .A(n67371), .B(n67370), .Y(n67707) );
  NAND2X1 U70808 ( .A(n40267), .B(n67372), .Y(n67373) );
  NAND2X1 U70809 ( .A(n41719), .B(n67373), .Y(n67708) );
  NAND2X1 U70810 ( .A(n67707), .B(n67708), .Y(n67706) );
  NAND2X1 U70811 ( .A(n67440), .B(n67439), .Y(n67730) );
  NOR2X1 U70812 ( .A(n38168), .B(n67772), .Y(n67374) );
  NOR2X1 U70813 ( .A(n41006), .B(n67374), .Y(n67383) );
  NOR2X1 U70814 ( .A(n67771), .B(n67375), .Y(n67381) );
  NAND2X1 U70815 ( .A(n67377), .B(n67376), .Y(n67378) );
  NOR2X1 U70816 ( .A(n67379), .B(n67378), .Y(n67380) );
  NOR2X1 U70817 ( .A(n67381), .B(n67380), .Y(n67382) );
  NAND2X1 U70818 ( .A(n67383), .B(n67382), .Y(n67778) );
  INVX1 U70819 ( .A(n67778), .Y(n67727) );
  INVX1 U70820 ( .A(n67384), .Y(n67386) );
  NOR2X1 U70821 ( .A(n67386), .B(n67385), .Y(n67391) );
  INVX1 U70822 ( .A(n67387), .Y(n67388) );
  NOR2X1 U70823 ( .A(n67389), .B(n67388), .Y(n67390) );
  NAND2X1 U70824 ( .A(n67391), .B(n67390), .Y(n67392) );
  NAND2X1 U70825 ( .A(n67393), .B(n67392), .Y(n67394) );
  NOR2X1 U70826 ( .A(n67395), .B(n67394), .Y(n67401) );
  INVX1 U70827 ( .A(n67402), .Y(n67739) );
  NAND2X1 U70828 ( .A(n41240), .B(n67739), .Y(n67398) );
  NAND2X1 U70829 ( .A(n67739), .B(n67396), .Y(n67397) );
  NAND2X1 U70830 ( .A(n67398), .B(n67397), .Y(n67399) );
  NOR2X1 U70831 ( .A(n67738), .B(n67399), .Y(n67400) );
  NOR2X1 U70832 ( .A(n67401), .B(n67400), .Y(n67404) );
  NAND2X1 U70833 ( .A(n67403), .B(n67402), .Y(n67734) );
  NAND2X1 U70834 ( .A(n67404), .B(n67734), .Y(n67733) );
  INVX1 U70835 ( .A(n67733), .Y(n68092) );
  INVX1 U70836 ( .A(n67762), .Y(n67759) );
  NAND2X1 U70837 ( .A(n67759), .B(n68113), .Y(n67414) );
  NOR2X1 U70838 ( .A(n67406), .B(n67405), .Y(n67408) );
  NOR2X1 U70839 ( .A(n67408), .B(n67407), .Y(n67409) );
  NOR2X1 U70840 ( .A(n67759), .B(n67409), .Y(n67411) );
  NAND2X1 U70841 ( .A(n67411), .B(n67410), .Y(n67412) );
  NAND2X1 U70842 ( .A(n67760), .B(n67412), .Y(n67413) );
  NAND2X1 U70843 ( .A(n67414), .B(n67413), .Y(n67758) );
  INVX1 U70844 ( .A(n67758), .Y(n68118) );
  INVX1 U70845 ( .A(n67415), .Y(n67418) );
  NAND2X1 U70846 ( .A(n67416), .B(n68107), .Y(n67417) );
  NAND2X1 U70847 ( .A(n67418), .B(n67417), .Y(n67755) );
  XNOR2X1 U70848 ( .A(n67755), .B(n41705), .Y(n67431) );
  INVX1 U70849 ( .A(n72383), .Y(n72387) );
  NAND2X1 U70850 ( .A(n67418), .B(n43604), .Y(n72310) );
  NAND2X1 U70851 ( .A(n41900), .B(n72370), .Y(n67420) );
  INVX1 U70852 ( .A(n72310), .Y(n72333) );
  NAND2X1 U70853 ( .A(n72333), .B(n72383), .Y(n67419) );
  NAND2X1 U70854 ( .A(n67420), .B(n67419), .Y(n67425) );
  NAND2X1 U70855 ( .A(n41900), .B(n67421), .Y(n67423) );
  INVX1 U70856 ( .A(n72373), .Y(n72371) );
  NAND2X1 U70857 ( .A(n41900), .B(n41685), .Y(n67422) );
  NAND2X1 U70858 ( .A(n67423), .B(n67422), .Y(n67424) );
  NOR2X1 U70859 ( .A(n67425), .B(n67424), .Y(n67430) );
  NAND2X1 U70860 ( .A(n72372), .B(n67426), .Y(n67427) );
  NOR2X1 U70861 ( .A(n72371), .B(n67427), .Y(n67428) );
  NAND2X1 U70862 ( .A(n72333), .B(n67428), .Y(n67429) );
  XNOR2X1 U70863 ( .A(n67752), .B(n41684), .Y(n68367) );
  INVX1 U70864 ( .A(n68367), .Y(n68653) );
  XNOR2X1 U70865 ( .A(n67431), .B(n68653), .Y(n68119) );
  XNOR2X1 U70866 ( .A(n68119), .B(n41713), .Y(n67432) );
  XNOR2X1 U70867 ( .A(n68118), .B(n67432), .Y(n68094) );
  XNOR2X1 U70868 ( .A(n68094), .B(n41714), .Y(n67433) );
  XNOR2X1 U70869 ( .A(n68092), .B(n67433), .Y(n67779) );
  NAND2X1 U70870 ( .A(n43491), .B(n43934), .Y(n68142) );
  XNOR2X1 U70871 ( .A(n68142), .B(n41514), .Y(n67434) );
  XNOR2X1 U70872 ( .A(n67779), .B(n67434), .Y(n67435) );
  XNOR2X1 U70873 ( .A(n67727), .B(n67435), .Y(n67450) );
  INVX1 U70874 ( .A(n67440), .Y(n67725) );
  NAND2X1 U70875 ( .A(n67450), .B(n67731), .Y(n67438) );
  NOR2X1 U70876 ( .A(n67723), .B(n67438), .Y(n67454) );
  OR2X1 U70877 ( .A(n67450), .B(n67730), .Y(n67452) );
  NOR2X1 U70878 ( .A(n67442), .B(n67441), .Y(n67443) );
  NAND2X1 U70879 ( .A(n67443), .B(n40994), .Y(n67444) );
  NAND2X1 U70880 ( .A(n67445), .B(n67444), .Y(n67446) );
  NAND2X1 U70881 ( .A(n41001), .B(n67446), .Y(n67447) );
  NAND2X1 U70882 ( .A(n67448), .B(n67447), .Y(n67449) );
  OR2X1 U70883 ( .A(n67450), .B(n67449), .Y(n67451) );
  NAND2X1 U70884 ( .A(n67452), .B(n67451), .Y(n67453) );
  NOR2X1 U70885 ( .A(n67454), .B(n67453), .Y(n67713) );
  XNOR2X1 U70886 ( .A(n67713), .B(n41519), .Y(n67705) );
  INVX1 U70887 ( .A(n67715), .Y(n67457) );
  NAND2X1 U70888 ( .A(n67459), .B(n67456), .Y(n67714) );
  INVX1 U70889 ( .A(n67455), .Y(n67718) );
  INVX1 U70890 ( .A(n67456), .Y(n67458) );
  NOR2X1 U70891 ( .A(n67458), .B(n67457), .Y(n67460) );
  NAND2X1 U70892 ( .A(n67460), .B(n67459), .Y(n67461) );
  NAND2X1 U70893 ( .A(n43972), .B(n38312), .Y(n67710) );
  INVX1 U70894 ( .A(n67710), .Y(n67462) );
  XNOR2X1 U70895 ( .A(n67712), .B(n67462), .Y(n67463) );
  XNOR2X1 U70896 ( .A(n67705), .B(n67463), .Y(n67464) );
  NAND2X1 U70897 ( .A(n43774), .B(n43992), .Y(n67693) );
  INVX1 U70898 ( .A(n67693), .Y(n67478) );
  NOR2X1 U70899 ( .A(n67478), .B(n41165), .Y(n67469) );
  NAND2X1 U70900 ( .A(n67466), .B(n39461), .Y(n67467) );
  NOR2X1 U70901 ( .A(n67478), .B(n67467), .Y(n67468) );
  NOR2X1 U70902 ( .A(n67469), .B(n67468), .Y(n67470) );
  NOR2X1 U70903 ( .A(n39486), .B(n67470), .Y(n67472) );
  NAND2X1 U70904 ( .A(n67683), .B(n67682), .Y(n67471) );
  NAND2X1 U70905 ( .A(n67472), .B(n67471), .Y(n67476) );
  NOR2X1 U70906 ( .A(n67690), .B(n67693), .Y(n67474) );
  NAND2X1 U70907 ( .A(n67474), .B(n67473), .Y(n67475) );
  NAND2X1 U70908 ( .A(n67476), .B(n67475), .Y(n67487) );
  NAND2X1 U70909 ( .A(n67693), .B(n67689), .Y(n67477) );
  NOR2X1 U70910 ( .A(n67682), .B(n67477), .Y(n67482) );
  NAND2X1 U70911 ( .A(n41522), .B(n67479), .Y(n67480) );
  NOR2X1 U70912 ( .A(n39779), .B(n67480), .Y(n67481) );
  NOR2X1 U70913 ( .A(n67482), .B(n67481), .Y(n67485) );
  NAND2X1 U70914 ( .A(n67690), .B(n67684), .Y(n67483) );
  NAND2X1 U70915 ( .A(n41522), .B(n67483), .Y(n67484) );
  NAND2X1 U70916 ( .A(n67485), .B(n67484), .Y(n67486) );
  NOR2X1 U70917 ( .A(n67487), .B(n67486), .Y(n67488) );
  XNOR2X1 U70918 ( .A(n40563), .B(n67488), .Y(n67796) );
  NAND2X1 U70919 ( .A(n43795), .B(n44000), .Y(n67795) );
  NAND2X1 U70920 ( .A(n42711), .B(n44008), .Y(n67792) );
  INVX1 U70921 ( .A(n67792), .Y(n67802) );
  XNOR2X1 U70922 ( .A(n67795), .B(n67802), .Y(n67489) );
  XNOR2X1 U70923 ( .A(n67796), .B(n67489), .Y(n67490) );
  XNOR2X1 U70924 ( .A(n67789), .B(n67490), .Y(n67806) );
  NOR2X1 U70925 ( .A(n67492), .B(n67491), .Y(n67498) );
  NOR2X1 U70926 ( .A(n67494), .B(n67493), .Y(n67496) );
  NOR2X1 U70927 ( .A(n67496), .B(n67495), .Y(n67497) );
  NOR2X1 U70928 ( .A(n67498), .B(n67497), .Y(n67501) );
  NAND2X1 U70929 ( .A(n67499), .B(n67502), .Y(n67500) );
  INVX1 U70930 ( .A(n67502), .Y(n67504) );
  NAND2X1 U70931 ( .A(n42651), .B(n44017), .Y(n67816) );
  XNOR2X1 U70932 ( .A(n67505), .B(n67826), .Y(n67678) );
  OR2X1 U70933 ( .A(n67508), .B(n67507), .Y(n67509) );
  NAND2X1 U70934 ( .A(n67510), .B(n67509), .Y(n67511) );
  XNOR2X1 U70935 ( .A(n67817), .B(n67815), .Y(n67513) );
  XNOR2X1 U70936 ( .A(n67514), .B(n67513), .Y(n67834) );
  NOR2X1 U70937 ( .A(n41403), .B(n67832), .Y(n67516) );
  NAND2X1 U70938 ( .A(n67834), .B(n67833), .Y(n67824) );
  NAND2X1 U70939 ( .A(n67516), .B(n67824), .Y(n67677) );
  XNOR2X1 U70940 ( .A(n67677), .B(n37416), .Y(n67517) );
  XNOR2X1 U70941 ( .A(n67678), .B(n67517), .Y(n67518) );
  XNOR2X1 U70942 ( .A(n41377), .B(n67518), .Y(n67672) );
  NOR2X1 U70943 ( .A(n67520), .B(n67519), .Y(n67526) );
  NOR2X1 U70944 ( .A(n67522), .B(n67521), .Y(n67524) );
  NOR2X1 U70945 ( .A(n67524), .B(n67523), .Y(n67525) );
  NOR2X1 U70946 ( .A(n67526), .B(n67525), .Y(n67530) );
  INVX1 U70947 ( .A(n67531), .Y(n67528) );
  NAND2X1 U70948 ( .A(n67528), .B(n67527), .Y(n67529) );
  NAND2X1 U70949 ( .A(n67530), .B(n67529), .Y(n67667) );
  NAND2X1 U70950 ( .A(n67532), .B(n67531), .Y(n67666) );
  NAND2X1 U70951 ( .A(n67667), .B(n67666), .Y(n67671) );
  XNOR2X1 U70952 ( .A(n67672), .B(n67671), .Y(n67533) );
  XNOR2X1 U70953 ( .A(n67534), .B(n67533), .Y(n67535) );
  XOR2X1 U70954 ( .A(n68012), .B(n67535), .Y(n68010) );
  INVX1 U70955 ( .A(n68010), .Y(n68019) );
  NAND2X1 U70956 ( .A(n67536), .B(n67537), .Y(n67538) );
  NAND2X1 U70957 ( .A(n43567), .B(n67849), .Y(n67847) );
  NAND2X1 U70958 ( .A(n43567), .B(n67847), .Y(n67541) );
  NOR2X1 U70959 ( .A(n67850), .B(n67541), .Y(n67542) );
  NOR2X1 U70960 ( .A(n67543), .B(n67542), .Y(n67544) );
  XNOR2X1 U70961 ( .A(n68019), .B(n67544), .Y(n67856) );
  NOR2X1 U70962 ( .A(n67545), .B(n43589), .Y(n67547) );
  NAND2X1 U70963 ( .A(n67550), .B(n38212), .Y(n67553) );
  NOR2X1 U70964 ( .A(n67554), .B(n43588), .Y(n67551) );
  NAND2X1 U70965 ( .A(n43576), .B(n67661), .Y(n67557) );
  NAND2X1 U70966 ( .A(n67556), .B(n67555), .Y(n67657) );
  NOR2X1 U70967 ( .A(n67557), .B(n67558), .Y(n67562) );
  NAND2X1 U70968 ( .A(n67655), .B(n39958), .Y(n67560) );
  NAND2X1 U70969 ( .A(n67658), .B(n67558), .Y(n67559) );
  NOR2X1 U70970 ( .A(n67560), .B(n67559), .Y(n67561) );
  XNOR2X1 U70971 ( .A(n68264), .B(n43537), .Y(n67571) );
  NOR2X1 U70972 ( .A(n39798), .B(n43541), .Y(n67566) );
  NAND2X1 U70973 ( .A(n67564), .B(n36405), .Y(n67565) );
  OR2X1 U70974 ( .A(n67566), .B(n67565), .Y(n67569) );
  NAND2X1 U70975 ( .A(n67569), .B(n67567), .Y(n67568) );
  NOR2X1 U70976 ( .A(n36751), .B(n67650), .Y(n67570) );
  XNOR2X1 U70977 ( .A(n67571), .B(n67570), .Y(n68585) );
  XNOR2X1 U70978 ( .A(n67572), .B(n36705), .Y(n67573) );
  INVX1 U70979 ( .A(n67638), .Y(n67637) );
  XNOR2X1 U70980 ( .A(n43633), .B(n43546), .Y(n71810) );
  XNOR2X1 U70981 ( .A(n71810), .B(n43666), .Y(n67574) );
  XNOR2X1 U70982 ( .A(n67637), .B(n67574), .Y(n67578) );
  NOR2X1 U70983 ( .A(n43545), .B(n67642), .Y(n67577) );
  NAND2X1 U70984 ( .A(n43545), .B(n67642), .Y(n67639) );
  XNOR2X1 U70985 ( .A(n67578), .B(n67870), .Y(n67579) );
  XNOR2X1 U70986 ( .A(n67630), .B(n67579), .Y(n67623) );
  XNOR2X1 U70987 ( .A(n67623), .B(n43643), .Y(n67580) );
  XNOR2X1 U70988 ( .A(n43655), .B(n67626), .Y(n67618) );
  NOR2X1 U70989 ( .A(n43653), .B(n67585), .Y(n67582) );
  NAND2X1 U70990 ( .A(n67584), .B(n67583), .Y(n67940) );
  NAND2X1 U70991 ( .A(n43653), .B(n67585), .Y(n67939) );
  NAND2X1 U70992 ( .A(n67586), .B(n67939), .Y(n67625) );
  XNOR2X1 U70993 ( .A(n43528), .B(n38924), .Y(n67587) );
  XOR2X1 U70994 ( .A(n67618), .B(n67587), .Y(n67890) );
  XNOR2X1 U70995 ( .A(n67588), .B(n67890), .Y(n67589) );
  XNOR2X1 U70996 ( .A(n41094), .B(n67589), .Y(n67898) );
  XNOR2X1 U70997 ( .A(n67898), .B(n43509), .Y(n67594) );
  INVX1 U70998 ( .A(n67590), .Y(n67592) );
  NAND2X1 U70999 ( .A(n43506), .B(n67592), .Y(n67922) );
  NAND2X1 U71000 ( .A(n67922), .B(n67923), .Y(n67899) );
  XNOR2X1 U71001 ( .A(n67613), .B(n43693), .Y(n67598) );
  NOR2X1 U71002 ( .A(n67610), .B(n67595), .Y(n67596) );
  NOR2X1 U71003 ( .A(n36791), .B(n67596), .Y(n67597) );
  XNOR2X1 U71004 ( .A(n67598), .B(n67597), .Y(n67605) );
  XNOR2X1 U71005 ( .A(n67605), .B(n43708), .Y(n67599) );
  XNOR2X1 U71006 ( .A(n67601), .B(n67600), .Y(n67602) );
  XNOR2X1 U71007 ( .A(n67602), .B(n42012), .Y(n67603) );
  MX2X1 U71008 ( .A(n67604), .B(n67603), .S0(n43719), .Y(u_muldiv_result_r[16]) );
  NAND2X1 U71009 ( .A(u_muldiv_mult_result_q[16]), .B(n44632), .Y(n13989) );
  NAND2X1 U71010 ( .A(n67605), .B(n43711), .Y(n67917) );
  NOR2X1 U71011 ( .A(n67606), .B(n43696), .Y(n67610) );
  NOR2X1 U71012 ( .A(n67610), .B(n67609), .Y(n67612) );
  NOR2X1 U71013 ( .A(n67612), .B(n67611), .Y(n67615) );
  NOR2X1 U71014 ( .A(n67613), .B(n43696), .Y(n67614) );
  OR2X1 U71015 ( .A(n67615), .B(n67614), .Y(n68539) );
  NAND2X1 U71016 ( .A(n67617), .B(n67616), .Y(n67619) );
  NAND2X1 U71017 ( .A(n43522), .B(n67620), .Y(n67927) );
  NAND2X1 U71018 ( .A(n67619), .B(n67927), .Y(n67622) );
  INVX1 U71019 ( .A(n67620), .Y(n67621) );
  NAND2X1 U71020 ( .A(n67621), .B(n43530), .Y(n67926) );
  INVX1 U71021 ( .A(n67886), .Y(n67883) );
  NAND2X1 U71022 ( .A(n67883), .B(n43660), .Y(n67938) );
  NAND2X1 U71023 ( .A(n38924), .B(n67938), .Y(n67627) );
  NAND2X1 U71024 ( .A(n43655), .B(n67626), .Y(n67936) );
  NAND2X1 U71025 ( .A(n67627), .B(n67936), .Y(n67930) );
  XNOR2X1 U71026 ( .A(n43633), .B(n67870), .Y(n67629) );
  XNOR2X1 U71027 ( .A(n43621), .B(n43546), .Y(n70560) );
  XNOR2X1 U71028 ( .A(n67628), .B(n36705), .Y(n67861) );
  NAND2X1 U71029 ( .A(n39057), .B(n41320), .Y(n67953) );
  INVX1 U71030 ( .A(n67631), .Y(n67633) );
  NOR2X1 U71031 ( .A(n67633), .B(n67632), .Y(n67635) );
  NAND2X1 U71032 ( .A(n67635), .B(n67634), .Y(n67636) );
  NAND2X1 U71033 ( .A(n43664), .B(n67636), .Y(n67954) );
  NAND2X1 U71034 ( .A(n43664), .B(n41320), .Y(n67955) );
  NAND2X1 U71035 ( .A(n43544), .B(n67637), .Y(n67973) );
  NOR2X1 U71036 ( .A(n43547), .B(n67640), .Y(n67641) );
  NOR2X1 U71037 ( .A(n39637), .B(n67641), .Y(n67645) );
  NAND2X1 U71038 ( .A(n67643), .B(n67642), .Y(n67644) );
  INVX1 U71039 ( .A(n71810), .Y(n72587) );
  XNOR2X1 U71040 ( .A(n72587), .B(n72088), .Y(n67867) );
  NAND2X1 U71041 ( .A(n68585), .B(n43559), .Y(n67649) );
  NAND2X1 U71042 ( .A(n67647), .B(n43559), .Y(n67648) );
  NAND2X1 U71043 ( .A(n67649), .B(n68495), .Y(n67991) );
  NAND2X1 U71044 ( .A(n67989), .B(n67991), .Y(n67980) );
  NAND2X1 U71045 ( .A(n43535), .B(n68264), .Y(n67652) );
  NAND2X1 U71046 ( .A(n67653), .B(n67657), .Y(n67654) );
  NOR2X1 U71047 ( .A(n67655), .B(n67654), .Y(n67656) );
  NOR2X1 U71048 ( .A(n67656), .B(n43574), .Y(n68000) );
  INVX1 U71049 ( .A(n67657), .Y(n67659) );
  NAND2X1 U71050 ( .A(n67659), .B(n67658), .Y(n67660) );
  NOR2X1 U71051 ( .A(n67661), .B(n67660), .Y(n67662) );
  NAND2X1 U71052 ( .A(n67662), .B(n67663), .Y(n67998) );
  NOR2X1 U71053 ( .A(n68000), .B(n40216), .Y(n67664) );
  NAND2X1 U71054 ( .A(n67664), .B(n67999), .Y(n68198) );
  XNOR2X1 U71055 ( .A(n43580), .B(n43583), .Y(n70726) );
  INVX1 U71056 ( .A(n67665), .Y(n67674) );
  XNOR2X1 U71057 ( .A(n67672), .B(n67674), .Y(n67668) );
  XNOR2X1 U71058 ( .A(n67668), .B(n41112), .Y(n67669) );
  NAND2X1 U71059 ( .A(n43593), .B(n67669), .Y(n68024) );
  NAND2X1 U71060 ( .A(n68011), .B(n68012), .Y(n68023) );
  NAND2X1 U71061 ( .A(n68024), .B(n68023), .Y(n68479) );
  INVX1 U71062 ( .A(n68479), .Y(n68487) );
  INVX1 U71063 ( .A(n67672), .Y(n67670) );
  NAND2X1 U71064 ( .A(n67671), .B(n67670), .Y(n67675) );
  NAND2X1 U71065 ( .A(n41112), .B(n67672), .Y(n67673) );
  NAND2X1 U71066 ( .A(n67675), .B(n39297), .Y(n68464) );
  INVX1 U71067 ( .A(n67676), .Y(n68047) );
  NAND2X1 U71068 ( .A(n67680), .B(n36731), .Y(n68045) );
  NAND2X1 U71069 ( .A(n37416), .B(n68045), .Y(n67681) );
  INVX1 U71070 ( .A(n68037), .Y(n68032) );
  NAND2X1 U71071 ( .A(n43796), .B(n44008), .Y(n68178) );
  XNOR2X1 U71072 ( .A(n68178), .B(n41527), .Y(n67788) );
  NOR2X1 U71073 ( .A(n67690), .B(n67689), .Y(n67687) );
  NOR2X1 U71074 ( .A(n67683), .B(n67682), .Y(n67685) );
  NAND2X1 U71075 ( .A(n67467), .B(n41165), .Y(n67684) );
  NOR2X1 U71076 ( .A(n67685), .B(n67684), .Y(n67686) );
  NOR2X1 U71077 ( .A(n39779), .B(n67688), .Y(n67692) );
  NAND2X1 U71078 ( .A(n67690), .B(n67689), .Y(n67691) );
  NOR2X1 U71079 ( .A(n39436), .B(n67693), .Y(n67695) );
  NOR2X1 U71080 ( .A(n40563), .B(n67693), .Y(n67694) );
  NOR2X1 U71081 ( .A(n67702), .B(n67698), .Y(n67701) );
  INVX1 U71082 ( .A(n67703), .Y(n67699) );
  NOR2X1 U71083 ( .A(n67699), .B(n67698), .Y(n67700) );
  INVX1 U71084 ( .A(n67702), .Y(n67704) );
  INVX1 U71085 ( .A(n68165), .Y(n67787) );
  NAND2X1 U71086 ( .A(n67709), .B(n67706), .Y(n68161) );
  OR2X1 U71087 ( .A(n67711), .B(n67710), .Y(n68160) );
  NAND2X1 U71088 ( .A(n68161), .B(n68160), .Y(n68082) );
  NAND2X1 U71089 ( .A(n67713), .B(n67712), .Y(n68322) );
  NOR2X1 U71090 ( .A(n39119), .B(n67713), .Y(n67720) );
  INVX1 U71091 ( .A(n67714), .Y(n67716) );
  NAND2X1 U71092 ( .A(n67716), .B(n67715), .Y(n67717) );
  NAND2X1 U71093 ( .A(n67718), .B(n67717), .Y(n67719) );
  NAND2X1 U71094 ( .A(n67720), .B(n67719), .Y(n67721) );
  NAND2X1 U71095 ( .A(n41519), .B(n67721), .Y(n68321) );
  NAND2X1 U71096 ( .A(n68322), .B(n68321), .Y(n68086) );
  INVX1 U71097 ( .A(n68142), .Y(n67729) );
  INVX1 U71098 ( .A(n67730), .Y(n67723) );
  NOR2X1 U71099 ( .A(n38736), .B(n67724), .Y(n67722) );
  NOR2X1 U71100 ( .A(n67725), .B(n67724), .Y(n67728) );
  XNOR2X1 U71101 ( .A(n67779), .B(n41514), .Y(n67726) );
  XNOR2X1 U71102 ( .A(n67727), .B(n67726), .Y(n68133) );
  INVX1 U71103 ( .A(n68133), .Y(n67732) );
  NAND2X1 U71104 ( .A(n67729), .B(n68140), .Y(n68407) );
  NAND2X1 U71105 ( .A(n67731), .B(n67730), .Y(n68136) );
  NAND2X1 U71106 ( .A(n68136), .B(n67732), .Y(n68397) );
  NAND2X1 U71107 ( .A(n68407), .B(n68397), .Y(n68085) );
  NAND2X1 U71108 ( .A(n43491), .B(n43943), .Y(n68138) );
  INVX1 U71109 ( .A(n68138), .Y(n68132) );
  INVX1 U71110 ( .A(n68094), .Y(n67740) );
  NAND2X1 U71111 ( .A(n67740), .B(n67733), .Y(n67745) );
  INVX1 U71112 ( .A(n67734), .Y(n67737) );
  NOR2X1 U71113 ( .A(n67735), .B(n67738), .Y(n67736) );
  NOR2X1 U71114 ( .A(n67737), .B(n67736), .Y(n67743) );
  NOR2X1 U71115 ( .A(n67739), .B(n67738), .Y(n67741) );
  NOR2X1 U71116 ( .A(n67741), .B(n67740), .Y(n67742) );
  NAND2X1 U71117 ( .A(n67743), .B(n67742), .Y(n67744) );
  NAND2X1 U71118 ( .A(n41714), .B(n67744), .Y(n68091) );
  NAND2X1 U71119 ( .A(n67745), .B(n68091), .Y(n68383) );
  NAND2X1 U71120 ( .A(n43928), .B(n43501), .Y(n68381) );
  INVX1 U71121 ( .A(n68381), .Y(n68099) );
  NAND2X1 U71122 ( .A(n43909), .B(n39653), .Y(n68103) );
  NAND2X1 U71123 ( .A(n41705), .B(n43604), .Y(n72334) );
  INVX1 U71124 ( .A(n72334), .Y(n72303) );
  NOR2X1 U71125 ( .A(n72333), .B(n72303), .Y(n67749) );
  NAND2X1 U71126 ( .A(n72382), .B(n67746), .Y(n67747) );
  NAND2X1 U71127 ( .A(n72387), .B(n67747), .Y(n72309) );
  NAND2X1 U71128 ( .A(n72303), .B(n72333), .Y(n67750) );
  NOR2X1 U71129 ( .A(n72309), .B(n67750), .Y(n67748) );
  NOR2X1 U71130 ( .A(n68107), .B(n67750), .Y(n67754) );
  NAND2X1 U71131 ( .A(n72309), .B(n72334), .Y(n67751) );
  NOR2X1 U71132 ( .A(n67752), .B(n67751), .Y(n67753) );
  XNOR2X1 U71133 ( .A(n68653), .B(n71853), .Y(n68377) );
  INVX1 U71134 ( .A(n68377), .Y(n68650) );
  XNOR2X1 U71135 ( .A(n68103), .B(n68650), .Y(n67757) );
  NAND2X1 U71136 ( .A(n68653), .B(n67755), .Y(n67756) );
  XNOR2X1 U71137 ( .A(n67757), .B(n41503), .Y(n68124) );
  NAND2X1 U71138 ( .A(n43918), .B(n39960), .Y(n68353) );
  INVX1 U71139 ( .A(n68353), .Y(n68117) );
  XNOR2X1 U71140 ( .A(n68124), .B(n68117), .Y(n67769) );
  NAND2X1 U71141 ( .A(n68119), .B(n67758), .Y(n67768) );
  INVX1 U71142 ( .A(n68114), .Y(n67765) );
  NAND2X1 U71143 ( .A(n67762), .B(n67761), .Y(n67763) );
  NAND2X1 U71144 ( .A(n67763), .B(n68113), .Y(n67764) );
  NAND2X1 U71145 ( .A(n67765), .B(n67764), .Y(n67766) );
  NAND2X1 U71146 ( .A(n41713), .B(n67766), .Y(n67767) );
  NAND2X1 U71147 ( .A(n67768), .B(n67767), .Y(n68125) );
  INVX1 U71148 ( .A(n68125), .Y(n68354) );
  XNOR2X1 U71149 ( .A(n67769), .B(n68354), .Y(n68382) );
  INVX1 U71150 ( .A(n68382), .Y(n68090) );
  XNOR2X1 U71151 ( .A(n68099), .B(n68090), .Y(n68088) );
  NAND2X1 U71152 ( .A(n43933), .B(n43496), .Y(n68342) );
  INVX1 U71153 ( .A(n68342), .Y(n68340) );
  XNOR2X1 U71154 ( .A(n68088), .B(n68340), .Y(n67770) );
  XNOR2X1 U71155 ( .A(n68383), .B(n67770), .Y(n67780) );
  NOR2X1 U71156 ( .A(n41006), .B(n67779), .Y(n67776) );
  NAND2X1 U71157 ( .A(n67772), .B(n67771), .Y(n67774) );
  NAND2X1 U71158 ( .A(n67774), .B(n67773), .Y(n67775) );
  NAND2X1 U71159 ( .A(n67776), .B(n67775), .Y(n67777) );
  NAND2X1 U71160 ( .A(n41514), .B(n67777), .Y(n68338) );
  NAND2X1 U71161 ( .A(n67779), .B(n67778), .Y(n68341) );
  NAND2X1 U71162 ( .A(n68338), .B(n68341), .Y(n68089) );
  XNOR2X1 U71163 ( .A(n67780), .B(n38788), .Y(n68139) );
  INVX1 U71164 ( .A(n68139), .Y(n68131) );
  XNOR2X1 U71165 ( .A(n68132), .B(n68131), .Y(n68084) );
  NAND2X1 U71166 ( .A(n43972), .B(n38310), .Y(n68325) );
  INVX1 U71167 ( .A(n68325), .Y(n67781) );
  XNOR2X1 U71168 ( .A(n68084), .B(n67781), .Y(n67782) );
  XNOR2X1 U71169 ( .A(n68085), .B(n67782), .Y(n67783) );
  NAND2X1 U71170 ( .A(n43774), .B(n44000), .Y(n68074) );
  NAND2X1 U71171 ( .A(n43477), .B(n43992), .Y(n68167) );
  NAND2X1 U71172 ( .A(n43982), .B(n38313), .Y(n68163) );
  INVX1 U71173 ( .A(n68163), .Y(n68421) );
  XNOR2X1 U71174 ( .A(n68074), .B(n68075), .Y(n67784) );
  XOR2X1 U71175 ( .A(n68419), .B(n67784), .Y(n67785) );
  XOR2X1 U71176 ( .A(n41207), .B(n67785), .Y(n67786) );
  INVX1 U71177 ( .A(n68179), .Y(n68171) );
  XNOR2X1 U71178 ( .A(n67788), .B(n68171), .Y(n67791) );
  NAND2X1 U71179 ( .A(n67796), .B(n67789), .Y(n68174) );
  INVX1 U71180 ( .A(n67795), .Y(n68173) );
  NAND2X1 U71181 ( .A(n68174), .B(n68175), .Y(n68067) );
  INVX1 U71182 ( .A(n68067), .Y(n67790) );
  XNOR2X1 U71183 ( .A(n67791), .B(n67790), .Y(n67803) );
  NOR2X1 U71184 ( .A(n40134), .B(n67792), .Y(n67800) );
  NAND2X1 U71185 ( .A(n67794), .B(n67793), .Y(n67798) );
  XNOR2X1 U71186 ( .A(n67796), .B(n67795), .Y(n67797) );
  XNOR2X1 U71187 ( .A(n67798), .B(n67797), .Y(n68068) );
  INVX1 U71188 ( .A(n68068), .Y(n67801) );
  NAND2X1 U71189 ( .A(n67801), .B(n39972), .Y(n68070) );
  INVX1 U71190 ( .A(n68070), .Y(n67799) );
  INVX1 U71191 ( .A(n68310), .Y(n68049) );
  NAND2X1 U71192 ( .A(n42653), .B(n44025), .Y(n68311) );
  INVX1 U71193 ( .A(n68311), .Y(n68064) );
  XNOR2X1 U71194 ( .A(n68049), .B(n68064), .Y(n67805) );
  NAND2X1 U71195 ( .A(n43772), .B(n44055), .Y(n68042) );
  INVX1 U71196 ( .A(n68042), .Y(n68038) );
  XNOR2X1 U71197 ( .A(n42995), .B(n68038), .Y(n67804) );
  XNOR2X1 U71198 ( .A(n67805), .B(n67804), .Y(n67823) );
  XNOR2X1 U71199 ( .A(n40134), .B(n67806), .Y(n67811) );
  NAND2X1 U71200 ( .A(n67807), .B(n67812), .Y(n67808) );
  NAND2X1 U71201 ( .A(n67816), .B(n67809), .Y(n67810) );
  NOR2X1 U71202 ( .A(n41187), .B(n41441), .Y(n67822) );
  NOR2X1 U71203 ( .A(n67816), .B(n67812), .Y(n67821) );
  INVX1 U71204 ( .A(n67813), .Y(n67815) );
  NOR2X1 U71205 ( .A(n67815), .B(n67814), .Y(n67819) );
  OR2X1 U71206 ( .A(n67817), .B(n67816), .Y(n67818) );
  NOR2X1 U71207 ( .A(n67819), .B(n67818), .Y(n67820) );
  NOR2X1 U71208 ( .A(n67821), .B(n67820), .Y(n68062) );
  NAND2X1 U71209 ( .A(n67822), .B(n68062), .Y(n68309) );
  INVX1 U71210 ( .A(n68309), .Y(n68051) );
  XNOR2X1 U71211 ( .A(n67823), .B(n68051), .Y(n67844) );
  INVX1 U71212 ( .A(n67824), .Y(n67827) );
  INVX1 U71213 ( .A(n67841), .Y(n67828) );
  NOR2X1 U71214 ( .A(n67828), .B(n68284), .Y(n67839) );
  INVX1 U71215 ( .A(n67834), .Y(n67830) );
  NOR2X1 U71216 ( .A(n67830), .B(n67829), .Y(n67831) );
  NOR2X1 U71217 ( .A(n67832), .B(n67831), .Y(n67836) );
  NAND2X1 U71218 ( .A(n67834), .B(n40307), .Y(n67835) );
  NAND2X1 U71219 ( .A(n67836), .B(n67835), .Y(n67837) );
  NAND2X1 U71220 ( .A(n67837), .B(n37356), .Y(n68282) );
  NAND2X1 U71221 ( .A(n43798), .B(n44048), .Y(n68059) );
  NAND2X1 U71222 ( .A(n68282), .B(n68059), .Y(n67838) );
  OR2X1 U71223 ( .A(n68059), .B(n68282), .Y(n67843) );
  NOR2X1 U71224 ( .A(n68284), .B(n68059), .Y(n67840) );
  NAND2X1 U71225 ( .A(n67841), .B(n67840), .Y(n67842) );
  XNOR2X1 U71226 ( .A(n67844), .B(n68052), .Y(n67845) );
  XNOR2X1 U71227 ( .A(n68032), .B(n67845), .Y(n68022) );
  XNOR2X1 U71228 ( .A(n43569), .B(n43594), .Y(n71079) );
  XNOR2X1 U71229 ( .A(n68022), .B(n71079), .Y(n67846) );
  XNOR2X1 U71230 ( .A(n70726), .B(n68007), .Y(n67854) );
  NAND2X1 U71231 ( .A(n43567), .B(n67850), .Y(n67848) );
  NAND2X1 U71232 ( .A(n67848), .B(n67847), .Y(n68018) );
  NAND2X1 U71233 ( .A(n67850), .B(n67849), .Y(n68009) );
  NOR2X1 U71234 ( .A(n68010), .B(n68009), .Y(n67852) );
  NOR2X1 U71235 ( .A(n68010), .B(n40670), .Y(n67851) );
  OR2X1 U71236 ( .A(n67852), .B(n67851), .Y(n67853) );
  NOR2X1 U71237 ( .A(n68018), .B(n67853), .Y(n68006) );
  XNOR2X1 U71238 ( .A(n67854), .B(n68006), .Y(n68197) );
  NAND2X1 U71239 ( .A(n67856), .B(n38100), .Y(n68008) );
  NAND2X1 U71240 ( .A(n43581), .B(n67856), .Y(n68004) );
  XNOR2X1 U71241 ( .A(n43542), .B(n40317), .Y(n67857) );
  XNOR2X1 U71242 ( .A(n67993), .B(n67983), .Y(n67858) );
  XOR2X1 U71243 ( .A(n40210), .B(n67858), .Y(n67859) );
  NAND2X1 U71244 ( .A(n38725), .B(n67860), .Y(n67981) );
  INVX1 U71245 ( .A(n67981), .Y(n67865) );
  NAND2X1 U71246 ( .A(n40085), .B(n67863), .Y(n67864) );
  NAND2X1 U71247 ( .A(n43619), .B(n67864), .Y(n67982) );
  NAND2X1 U71248 ( .A(n39952), .B(n67982), .Y(n67961) );
  NOR2X1 U71249 ( .A(n67865), .B(n67961), .Y(n67866) );
  XNOR2X1 U71250 ( .A(n67962), .B(n67866), .Y(n68255) );
  INVX1 U71251 ( .A(n68255), .Y(n67971) );
  XNOR2X1 U71252 ( .A(n67867), .B(n67971), .Y(n67868) );
  XNOR2X1 U71253 ( .A(n38913), .B(n67868), .Y(n67881) );
  XNOR2X1 U71254 ( .A(n67870), .B(n67869), .Y(n67880) );
  INVX1 U71255 ( .A(n67880), .Y(n67871) );
  NOR2X1 U71256 ( .A(n40414), .B(n36426), .Y(n67873) );
  NOR2X1 U71257 ( .A(n67874), .B(n67873), .Y(n67877) );
  NAND2X1 U71258 ( .A(n67875), .B(n43635), .Y(n67876) );
  NAND2X1 U71259 ( .A(n67876), .B(n67877), .Y(n67879) );
  NAND2X1 U71260 ( .A(n43631), .B(n67880), .Y(n67966) );
  XNOR2X1 U71261 ( .A(n67881), .B(n41057), .Y(n67882) );
  XNOR2X1 U71262 ( .A(n68210), .B(n67882), .Y(n67935) );
  NAND2X1 U71263 ( .A(n67885), .B(n67884), .Y(n68236) );
  NAND2X1 U71264 ( .A(n40142), .B(n67886), .Y(n68235) );
  NAND2X1 U71265 ( .A(n68236), .B(n68235), .Y(n67934) );
  XNOR2X1 U71266 ( .A(n43658), .B(n67934), .Y(n67887) );
  XOR2X1 U71267 ( .A(n67935), .B(n67887), .Y(n67931) );
  XNOR2X1 U71268 ( .A(n43528), .B(n67931), .Y(n67888) );
  XNOR2X1 U71269 ( .A(n67930), .B(n67888), .Y(n67889) );
  XNOR2X1 U71270 ( .A(n68219), .B(n43679), .Y(n67897) );
  XNOR2X1 U71271 ( .A(n41059), .B(n67890), .Y(n67891) );
  INVX1 U71272 ( .A(n68218), .Y(n67895) );
  NAND2X1 U71273 ( .A(n67893), .B(n67892), .Y(n67894) );
  NOR2X1 U71274 ( .A(n67895), .B(n67894), .Y(n67896) );
  XNOR2X1 U71275 ( .A(n67925), .B(n43508), .Y(n67902) );
  NOR2X1 U71276 ( .A(n41163), .B(n67899), .Y(n67900) );
  NOR2X1 U71277 ( .A(n41416), .B(n67900), .Y(n67901) );
  XNOR2X1 U71278 ( .A(n67902), .B(n67901), .Y(n67918) );
  XNOR2X1 U71279 ( .A(n67918), .B(n43693), .Y(n67903) );
  XNOR2X1 U71280 ( .A(n43715), .B(n36392), .Y(n67904) );
  XNOR2X1 U71281 ( .A(n67905), .B(n67904), .Y(n67910) );
  XNOR2X1 U71282 ( .A(n67907), .B(n67906), .Y(n67908) );
  XOR2X1 U71283 ( .A(n42022), .B(n67908), .Y(n67909) );
  MX2X1 U71284 ( .A(n67910), .B(n67909), .S0(n43719), .Y(u_muldiv_result_r[17]) );
  NAND2X1 U71285 ( .A(u_muldiv_mult_result_q[17]), .B(n44632), .Y(n13978) );
  OR2X1 U71286 ( .A(n43715), .B(n67915), .Y(n67911) );
  NAND2X1 U71287 ( .A(n67912), .B(n67911), .Y(n67913) );
  NAND2X1 U71288 ( .A(n36392), .B(n43711), .Y(n67916) );
  NAND2X1 U71289 ( .A(n43691), .B(n67918), .Y(n67920) );
  NAND2X1 U71290 ( .A(n68540), .B(n36402), .Y(n67919) );
  NAND2X1 U71291 ( .A(n67920), .B(n69225), .Y(n68229) );
  NOR2X1 U71292 ( .A(n43508), .B(n67925), .Y(n67921) );
  NOR2X1 U71293 ( .A(n41204), .B(n37994), .Y(n68222) );
  INVX1 U71294 ( .A(n67926), .Y(n67929) );
  INVX1 U71295 ( .A(n67932), .Y(n67933) );
  NAND2X1 U71296 ( .A(n43523), .B(n67933), .Y(n68232) );
  NAND2X1 U71297 ( .A(n36427), .B(n68232), .Y(n68824) );
  INVX1 U71298 ( .A(n67936), .Y(n67937) );
  NOR2X1 U71299 ( .A(n67947), .B(n67937), .Y(n67945) );
  INVX1 U71300 ( .A(n67938), .Y(n67942) );
  NOR2X1 U71301 ( .A(n67942), .B(n67941), .Y(n67944) );
  NAND2X1 U71302 ( .A(n36472), .B(n43659), .Y(n67943) );
  NAND2X1 U71303 ( .A(n67944), .B(n67943), .Y(n67946) );
  NAND2X1 U71304 ( .A(n43658), .B(n67946), .Y(n67950) );
  INVX1 U71305 ( .A(n67947), .Y(n67948) );
  NAND2X1 U71306 ( .A(n67948), .B(n43659), .Y(n67949) );
  NAND2X1 U71307 ( .A(n67950), .B(n67949), .Y(n68515) );
  NOR2X1 U71308 ( .A(n39888), .B(n68515), .Y(n68215) );
  XNOR2X1 U71309 ( .A(n71810), .B(n68255), .Y(n67951) );
  XOR2X1 U71310 ( .A(n67952), .B(n67951), .Y(n68207) );
  XNOR2X1 U71311 ( .A(n41057), .B(n68207), .Y(n67958) );
  INVX1 U71312 ( .A(n67953), .Y(n67957) );
  NAND2X1 U71313 ( .A(n67955), .B(n67954), .Y(n67956) );
  NOR2X1 U71314 ( .A(n67957), .B(n67956), .Y(n67960) );
  NAND2X1 U71315 ( .A(n43665), .B(n67958), .Y(n67959) );
  NAND2X1 U71316 ( .A(n67960), .B(n67959), .Y(n68247) );
  NAND2X1 U71317 ( .A(n68248), .B(n68247), .Y(n68241) );
  XNOR2X1 U71318 ( .A(n67963), .B(n67962), .Y(n67964) );
  XNOR2X1 U71319 ( .A(n39160), .B(n67964), .Y(n67969) );
  NOR2X1 U71320 ( .A(n67969), .B(n43639), .Y(n67968) );
  NAND2X1 U71321 ( .A(n67966), .B(n67965), .Y(n67967) );
  INVX1 U71322 ( .A(n67969), .Y(n67970) );
  NAND2X1 U71323 ( .A(n67971), .B(n43550), .Y(n68256) );
  INVX1 U71324 ( .A(n67972), .Y(n67975) );
  INVX1 U71325 ( .A(n67973), .Y(n67974) );
  NOR2X1 U71326 ( .A(n67975), .B(n67974), .Y(n67977) );
  NAND2X1 U71327 ( .A(n43544), .B(n68255), .Y(n67976) );
  NAND2X1 U71328 ( .A(n67977), .B(n67976), .Y(n67978) );
  NAND2X1 U71329 ( .A(n68256), .B(n67978), .Y(n68566) );
  XNOR2X1 U71330 ( .A(n43560), .B(n68200), .Y(n67979) );
  NOR2X1 U71331 ( .A(n71794), .B(n68583), .Y(n67988) );
  NAND2X1 U71332 ( .A(n67990), .B(n67989), .Y(n67984) );
  NOR2X1 U71333 ( .A(n68495), .B(n67984), .Y(n67986) );
  NAND2X1 U71334 ( .A(n43562), .B(n71794), .Y(n67985) );
  NOR2X1 U71335 ( .A(n67986), .B(n67985), .Y(n67987) );
  NOR2X1 U71336 ( .A(n67988), .B(n67987), .Y(n67995) );
  INVX1 U71337 ( .A(n67989), .Y(n68497) );
  INVX1 U71338 ( .A(n67990), .Y(n68496) );
  INVX1 U71339 ( .A(n68495), .Y(n68584) );
  NAND2X1 U71340 ( .A(n43559), .B(n67991), .Y(n68501) );
  NAND2X1 U71341 ( .A(n68582), .B(n68501), .Y(n67992) );
  NAND2X1 U71342 ( .A(n67993), .B(n67992), .Y(n67994) );
  NAND2X1 U71343 ( .A(n67995), .B(n67994), .Y(n68204) );
  XNOR2X1 U71344 ( .A(n43589), .B(n68007), .Y(n67996) );
  XOR2X1 U71345 ( .A(n67997), .B(n68196), .Y(n68001) );
  NOR2X1 U71346 ( .A(n68000), .B(n39635), .Y(n68002) );
  NAND2X1 U71347 ( .A(n68002), .B(n68001), .Y(n68491) );
  NAND2X1 U71348 ( .A(n68491), .B(n40002), .Y(n68003) );
  XNOR2X1 U71349 ( .A(n43580), .B(n68003), .Y(n68195) );
  NAND2X1 U71350 ( .A(n68008), .B(n43587), .Y(n68271) );
  XNOR2X1 U71351 ( .A(n68599), .B(n43582), .Y(n68194) );
  NOR2X1 U71352 ( .A(n43568), .B(n67852), .Y(n68017) );
  NAND2X1 U71353 ( .A(n68012), .B(n68011), .Y(n68015) );
  XNOR2X1 U71354 ( .A(n68022), .B(n43594), .Y(n68013) );
  XOR2X1 U71355 ( .A(n68015), .B(n68014), .Y(n68020) );
  NOR2X1 U71356 ( .A(n43568), .B(n68020), .Y(n68016) );
  NOR2X1 U71357 ( .A(n68017), .B(n68016), .Y(n68021) );
  NAND2X1 U71358 ( .A(n68277), .B(n68021), .Y(n68278) );
  XNOR2X1 U71359 ( .A(n68278), .B(n43569), .Y(n68193) );
  NOR2X1 U71360 ( .A(n68477), .B(n42993), .Y(n68026) );
  NAND2X1 U71361 ( .A(n68024), .B(n68023), .Y(n68025) );
  NOR2X1 U71362 ( .A(n68026), .B(n68025), .Y(n68027) );
  NOR2X1 U71363 ( .A(n68027), .B(n41622), .Y(n68192) );
  XNOR2X1 U71364 ( .A(n68311), .B(n68038), .Y(n68029) );
  XNOR2X1 U71365 ( .A(n68309), .B(n68049), .Y(n68028) );
  XNOR2X1 U71366 ( .A(n68029), .B(n68028), .Y(n68030) );
  XNOR2X1 U71367 ( .A(n68030), .B(n68052), .Y(n68031) );
  INVX1 U71368 ( .A(n68465), .Y(n68468) );
  NOR2X1 U71369 ( .A(n43618), .B(n68468), .Y(n68033) );
  NAND2X1 U71370 ( .A(n68033), .B(n68464), .Y(n68036) );
  NOR2X1 U71371 ( .A(n68465), .B(n42996), .Y(n68034) );
  NAND2X1 U71372 ( .A(n40027), .B(n68034), .Y(n68035) );
  NAND2X1 U71373 ( .A(n68036), .B(n68035), .Y(n68483) );
  NAND2X1 U71374 ( .A(n68038), .B(n68037), .Y(n68458) );
  NOR2X1 U71375 ( .A(n68047), .B(n68038), .Y(n68041) );
  NOR2X1 U71376 ( .A(n39543), .B(n68039), .Y(n68040) );
  NAND2X1 U71377 ( .A(n68041), .B(n68040), .Y(n68044) );
  NAND2X1 U71378 ( .A(n68042), .B(n38928), .Y(n68043) );
  XNOR2X1 U71379 ( .A(n68311), .B(n68049), .Y(n68050) );
  XNOR2X1 U71380 ( .A(n68051), .B(n68050), .Y(n68060) );
  XNOR2X1 U71381 ( .A(n68060), .B(n68052), .Y(n68053) );
  NAND2X1 U71382 ( .A(n68054), .B(n68053), .Y(n68459) );
  NAND2X1 U71383 ( .A(n68459), .B(n68458), .Y(n68189) );
  NAND2X1 U71384 ( .A(n68060), .B(n68059), .Y(n68058) );
  NAND2X1 U71385 ( .A(n68055), .B(n68283), .Y(n68056) );
  NAND2X1 U71386 ( .A(n68056), .B(n68282), .Y(n68057) );
  NAND2X1 U71387 ( .A(n68058), .B(n68057), .Y(n68061) );
  INVX1 U71388 ( .A(n68059), .Y(n68289) );
  INVX1 U71389 ( .A(n68060), .Y(n68288) );
  NAND2X1 U71390 ( .A(n68289), .B(n68288), .Y(n68281) );
  NAND2X1 U71391 ( .A(n68061), .B(n68281), .Y(n68306) );
  NAND2X1 U71392 ( .A(n68064), .B(n68310), .Y(n68300) );
  NAND2X1 U71393 ( .A(n68064), .B(n68063), .Y(n68301) );
  NAND2X1 U71394 ( .A(n68300), .B(n68301), .Y(n68065) );
  NOR2X1 U71395 ( .A(n37387), .B(n68065), .Y(n68066) );
  XNOR2X1 U71396 ( .A(n41728), .B(n68066), .Y(n68186) );
  NAND2X1 U71397 ( .A(n41527), .B(n68739), .Y(n68294) );
  INVX1 U71398 ( .A(n68294), .Y(n68737) );
  NAND2X1 U71399 ( .A(n40134), .B(n68068), .Y(n68069) );
  NAND2X1 U71400 ( .A(n68069), .B(n44008), .Y(n68071) );
  NAND2X1 U71401 ( .A(n68071), .B(n68070), .Y(n68072) );
  NAND2X1 U71402 ( .A(n41527), .B(n68072), .Y(n68295) );
  INVX1 U71403 ( .A(n68295), .Y(n68736) );
  NOR2X1 U71404 ( .A(n68737), .B(n68736), .Y(n68073) );
  NAND2X1 U71405 ( .A(n68073), .B(n68740), .Y(n68445) );
  NAND2X1 U71406 ( .A(n43795), .B(n44017), .Y(n68442) );
  INVX1 U71407 ( .A(n68074), .Y(n68077) );
  INVX1 U71408 ( .A(n68419), .Y(n68162) );
  XNOR2X1 U71409 ( .A(n68075), .B(n68162), .Y(n68076) );
  NOR2X1 U71410 ( .A(n41439), .B(n41384), .Y(n68080) );
  NAND2X1 U71411 ( .A(n68079), .B(n68078), .Y(n68435) );
  NAND2X1 U71412 ( .A(n68435), .B(n68080), .Y(n68081) );
  XNOR2X1 U71413 ( .A(n68081), .B(n42034), .Y(n68170) );
  NAND2X1 U71414 ( .A(n43477), .B(n44000), .Y(n68430) );
  NOR2X1 U71415 ( .A(n68324), .B(n68086), .Y(n68087) );
  OR2X1 U71416 ( .A(n68087), .B(n68325), .Y(n68151) );
  NAND2X1 U71417 ( .A(n68149), .B(n68151), .Y(n68320) );
  NAND2X1 U71418 ( .A(n68339), .B(n68089), .Y(n68636) );
  NAND2X1 U71419 ( .A(n68090), .B(n68383), .Y(n68102) );
  INVX1 U71420 ( .A(n68091), .Y(n68096) );
  NAND2X1 U71421 ( .A(n68092), .B(n68382), .Y(n68093) );
  NOR2X1 U71422 ( .A(n68096), .B(n68093), .Y(n68098) );
  NAND2X1 U71423 ( .A(n68382), .B(n68094), .Y(n68095) );
  NOR2X1 U71424 ( .A(n68096), .B(n68095), .Y(n68097) );
  NOR2X1 U71425 ( .A(n68098), .B(n68097), .Y(n68100) );
  NAND2X1 U71426 ( .A(n68100), .B(n68099), .Y(n68101) );
  NAND2X1 U71427 ( .A(n68102), .B(n68101), .Y(n68388) );
  INVX1 U71428 ( .A(n68388), .Y(n68333) );
  INVX1 U71429 ( .A(n68103), .Y(n68106) );
  NAND2X1 U71430 ( .A(n68106), .B(n68377), .Y(n68105) );
  NAND2X1 U71431 ( .A(n68106), .B(n41503), .Y(n68104) );
  NAND2X1 U71432 ( .A(n68105), .B(n68104), .Y(n68364) );
  XNOR2X1 U71433 ( .A(n68364), .B(n68650), .Y(n68112) );
  NAND2X1 U71434 ( .A(n68106), .B(n43604), .Y(n72400) );
  INVX1 U71435 ( .A(n72400), .Y(n72397) );
  XNOR2X1 U71436 ( .A(n41510), .B(n72397), .Y(n68110) );
  NAND2X1 U71437 ( .A(n72303), .B(n68367), .Y(n68109) );
  NAND2X1 U71438 ( .A(n72309), .B(n68107), .Y(n68108) );
  NAND2X1 U71439 ( .A(n72333), .B(n68108), .Y(n68654) );
  INVX1 U71440 ( .A(n68654), .Y(n72302) );
  NAND2X1 U71441 ( .A(n72302), .B(n72303), .Y(n72304) );
  NAND2X1 U71442 ( .A(n68109), .B(n72304), .Y(n72396) );
  INVX1 U71443 ( .A(n72396), .Y(n72401) );
  XNOR2X1 U71444 ( .A(n68110), .B(n72401), .Y(n68111) );
  XNOR2X1 U71445 ( .A(n68112), .B(n68111), .Y(n68358) );
  NOR2X1 U71446 ( .A(n68114), .B(n68113), .Y(n68116) );
  NAND2X1 U71447 ( .A(n68117), .B(n43912), .Y(n68115) );
  NOR2X1 U71448 ( .A(n68116), .B(n68115), .Y(n68123) );
  NAND2X1 U71449 ( .A(n68117), .B(n68124), .Y(n68357) );
  NOR2X1 U71450 ( .A(n68118), .B(n68353), .Y(n68120) );
  NAND2X1 U71451 ( .A(n68120), .B(n68119), .Y(n68121) );
  NAND2X1 U71452 ( .A(n68357), .B(n68121), .Y(n68122) );
  NOR2X1 U71453 ( .A(n68123), .B(n68122), .Y(n68126) );
  NAND2X1 U71454 ( .A(n68125), .B(n68124), .Y(n68352) );
  NAND2X1 U71455 ( .A(n68126), .B(n68352), .Y(n68351) );
  NAND2X1 U71456 ( .A(n43942), .B(n43497), .Y(n68631) );
  XNOR2X1 U71457 ( .A(n68631), .B(n41716), .Y(n68127) );
  XNOR2X1 U71458 ( .A(n68379), .B(n68127), .Y(n68128) );
  XNOR2X1 U71459 ( .A(n68333), .B(n68128), .Y(n68398) );
  NAND2X1 U71460 ( .A(n38481), .B(n68398), .Y(n68402) );
  NAND2X1 U71461 ( .A(n68340), .B(n68635), .Y(n68334) );
  NAND2X1 U71462 ( .A(n39466), .B(n68398), .Y(n68401) );
  NAND2X1 U71463 ( .A(n68636), .B(n68334), .Y(n68129) );
  OR2X1 U71464 ( .A(n68398), .B(n68129), .Y(n68130) );
  NOR2X1 U71465 ( .A(n68133), .B(n68138), .Y(n68135) );
  NOR2X1 U71466 ( .A(n68139), .B(n68133), .Y(n68134) );
  NOR2X1 U71467 ( .A(n41003), .B(n68137), .Y(n68144) );
  NAND2X1 U71468 ( .A(n68139), .B(n68138), .Y(n68396) );
  NAND2X1 U71469 ( .A(n68140), .B(n68396), .Y(n68141) );
  OR2X1 U71470 ( .A(n68142), .B(n68141), .Y(n68143) );
  NAND2X1 U71471 ( .A(n68144), .B(n68143), .Y(n68394) );
  XNOR2X1 U71472 ( .A(n68394), .B(n41523), .Y(n68145) );
  XNOR2X1 U71473 ( .A(n41236), .B(n68145), .Y(n68146) );
  NAND2X1 U71474 ( .A(n39396), .B(n68146), .Y(n68417) );
  INVX1 U71475 ( .A(n68417), .Y(n68148) );
  INVX1 U71476 ( .A(n68146), .Y(n68154) );
  NAND2X1 U71477 ( .A(n68154), .B(n68320), .Y(n68416) );
  NAND2X1 U71478 ( .A(n68416), .B(n68150), .Y(n68147) );
  NOR2X1 U71479 ( .A(n68148), .B(n68147), .Y(n68158) );
  OR2X1 U71480 ( .A(n68150), .B(n68416), .Y(n68156) );
  NOR2X1 U71481 ( .A(n39332), .B(n68150), .Y(n68152) );
  NAND2X1 U71482 ( .A(n68152), .B(n68151), .Y(n68153) );
  OR2X1 U71483 ( .A(n68154), .B(n68153), .Y(n68155) );
  NAND2X1 U71484 ( .A(n68156), .B(n68155), .Y(n68157) );
  NOR2X1 U71485 ( .A(n68158), .B(n68157), .Y(n68428) );
  XNOR2X1 U71486 ( .A(n68430), .B(n68428), .Y(n68159) );
  XNOR2X1 U71487 ( .A(n68427), .B(n68159), .Y(n68169) );
  XNOR2X1 U71488 ( .A(n68163), .B(n68162), .Y(n68164) );
  XNOR2X1 U71489 ( .A(n41207), .B(n68164), .Y(n68166) );
  NAND2X1 U71490 ( .A(n68166), .B(n68165), .Y(n68709) );
  NOR2X1 U71491 ( .A(n68166), .B(n68165), .Y(n68168) );
  OR2X1 U71492 ( .A(n68168), .B(n68167), .Y(n68712) );
  NAND2X1 U71493 ( .A(n68709), .B(n68712), .Y(n68429) );
  INVX1 U71494 ( .A(n68436), .Y(n68622) );
  XNOR2X1 U71495 ( .A(n68170), .B(n68622), .Y(n68441) );
  INVX1 U71496 ( .A(n68441), .Y(n68443) );
  XNOR2X1 U71497 ( .A(n68442), .B(n68443), .Y(n68183) );
  NAND2X1 U71498 ( .A(n68171), .B(n68178), .Y(n68177) );
  NAND2X1 U71499 ( .A(n68173), .B(n68172), .Y(n68175) );
  NAND2X1 U71500 ( .A(n68175), .B(n68174), .Y(n68176) );
  NAND2X1 U71501 ( .A(n68177), .B(n68176), .Y(n68182) );
  INVX1 U71502 ( .A(n68178), .Y(n68180) );
  NAND2X1 U71503 ( .A(n68180), .B(n68179), .Y(n68181) );
  NAND2X1 U71504 ( .A(n68182), .B(n68181), .Y(n68440) );
  INVX1 U71505 ( .A(n68440), .Y(n68444) );
  XNOR2X1 U71506 ( .A(n68183), .B(n68444), .Y(n68446) );
  INVX1 U71507 ( .A(n68446), .Y(n68743) );
  XNOR2X1 U71508 ( .A(n68445), .B(n68743), .Y(n68185) );
  NAND2X1 U71509 ( .A(n42654), .B(n44048), .Y(n68314) );
  NAND2X1 U71510 ( .A(n42712), .B(n44025), .Y(n68744) );
  XNOR2X1 U71511 ( .A(n68314), .B(n68744), .Y(n68184) );
  XNOR2X1 U71512 ( .A(n68185), .B(n68184), .Y(n68305) );
  XNOR2X1 U71513 ( .A(n68186), .B(n68305), .Y(n68187) );
  NAND2X1 U71514 ( .A(n43613), .B(n43772), .Y(n72536) );
  XNOR2X1 U71515 ( .A(n68768), .B(n40683), .Y(n68188) );
  XNOR2X1 U71516 ( .A(n68189), .B(n68188), .Y(n68482) );
  XNOR2X1 U71517 ( .A(n68482), .B(n43593), .Y(n68190) );
  XNOR2X1 U71518 ( .A(n68483), .B(n68190), .Y(n68191) );
  XNOR2X1 U71519 ( .A(n68192), .B(n68191), .Y(n68279) );
  INVX1 U71520 ( .A(n68276), .Y(n68272) );
  XNOR2X1 U71521 ( .A(n68194), .B(n68272), .Y(n69174) );
  INVX1 U71522 ( .A(n69174), .Y(n68796) );
  XNOR2X1 U71523 ( .A(n68195), .B(n68796), .Y(n68804) );
  NAND2X1 U71524 ( .A(n43535), .B(n68265), .Y(n68199) );
  NOR2X1 U71525 ( .A(n68199), .B(n40210), .Y(n68201) );
  NOR2X1 U71526 ( .A(n68202), .B(n68201), .Y(n68203) );
  XNOR2X1 U71527 ( .A(n40093), .B(n68203), .Y(n68588) );
  XNOR2X1 U71528 ( .A(n68204), .B(n68588), .Y(n68205) );
  XNOR2X1 U71529 ( .A(n71810), .B(n68567), .Y(n68206) );
  XNOR2X1 U71530 ( .A(n39470), .B(n68242), .Y(n68249) );
  XNOR2X1 U71531 ( .A(n43655), .B(n68516), .Y(n68213) );
  XNOR2X1 U71532 ( .A(n43666), .B(n68207), .Y(n68208) );
  XNOR2X1 U71533 ( .A(n68208), .B(n41057), .Y(n68209) );
  XNOR2X1 U71534 ( .A(n68210), .B(n68209), .Y(n68211) );
  NAND2X1 U71535 ( .A(n40168), .B(n68239), .Y(n68212) );
  NAND2X1 U71536 ( .A(n68211), .B(n39301), .Y(n68237) );
  XNOR2X1 U71537 ( .A(n68213), .B(n41036), .Y(n68214) );
  XNOR2X1 U71538 ( .A(n68215), .B(n68214), .Y(n68521) );
  XNOR2X1 U71539 ( .A(n39973), .B(n68522), .Y(n69542) );
  XNOR2X1 U71540 ( .A(n69542), .B(n38047), .Y(n68216) );
  XNOR2X1 U71541 ( .A(n43509), .B(n68216), .Y(n68220) );
  NOR2X1 U71542 ( .A(n43686), .B(n68219), .Y(n68217) );
  NAND2X1 U71543 ( .A(n68219), .B(n43684), .Y(n68860) );
  XNOR2X1 U71544 ( .A(n68220), .B(n36444), .Y(n68221) );
  XNOR2X1 U71545 ( .A(n68222), .B(n68221), .Y(n69226) );
  XNOR2X1 U71546 ( .A(n69226), .B(n43693), .Y(n68223) );
  XNOR2X1 U71547 ( .A(n68225), .B(n68224), .Y(n68226) );
  XNOR2X1 U71548 ( .A(n68226), .B(n42036), .Y(n68227) );
  MX2X1 U71549 ( .A(n68228), .B(n68227), .S0(n43719), .Y(u_muldiv_result_r[18]) );
  NAND2X1 U71550 ( .A(u_muldiv_mult_result_q[18]), .B(n44632), .Y(n13970) );
  NAND2X1 U71551 ( .A(n69226), .B(n43698), .Y(n68541) );
  NAND2X1 U71552 ( .A(n68541), .B(n68229), .Y(n68546) );
  NAND2X1 U71553 ( .A(n43677), .B(n69542), .Y(n68835) );
  NAND2X1 U71554 ( .A(n36523), .B(n43683), .Y(n68230) );
  NAND2X1 U71555 ( .A(n41095), .B(n68230), .Y(n68834) );
  NAND2X1 U71556 ( .A(n68521), .B(n43529), .Y(n68823) );
  NOR2X1 U71557 ( .A(n68521), .B(n43528), .Y(n68234) );
  NAND2X1 U71558 ( .A(n68232), .B(n68231), .Y(n68233) );
  OR2X1 U71559 ( .A(n68234), .B(n68233), .Y(n68876) );
  NAND2X1 U71560 ( .A(n68823), .B(n68876), .Y(n68830) );
  NAND2X1 U71561 ( .A(n39679), .B(n68235), .Y(n68238) );
  NAND2X1 U71562 ( .A(n68238), .B(n68237), .Y(n68240) );
  NAND2X1 U71563 ( .A(n68240), .B(n68239), .Y(n68244) );
  XNOR2X1 U71564 ( .A(n43666), .B(n39470), .Y(n68243) );
  NAND2X1 U71565 ( .A(n68245), .B(n39301), .Y(n68895) );
  NAND2X1 U71566 ( .A(n68244), .B(n68895), .Y(n69247) );
  INVX1 U71567 ( .A(n68245), .Y(n68246) );
  NAND2X1 U71568 ( .A(n43642), .B(n68246), .Y(n69251) );
  NOR2X1 U71569 ( .A(n39870), .B(n38946), .Y(n68251) );
  NAND2X1 U71570 ( .A(n68249), .B(n43670), .Y(n68250) );
  NAND2X1 U71571 ( .A(n68250), .B(n68251), .Y(n68558) );
  NOR2X1 U71572 ( .A(n68567), .B(n43639), .Y(n68252) );
  INVX1 U71573 ( .A(n68567), .Y(n68254) );
  INVX1 U71574 ( .A(n68560), .Y(n68555) );
  NAND2X1 U71575 ( .A(n43545), .B(n68254), .Y(n68259) );
  NAND2X1 U71576 ( .A(n38913), .B(n67976), .Y(n68257) );
  NAND2X1 U71577 ( .A(n68257), .B(n68256), .Y(n68562) );
  NAND2X1 U71578 ( .A(n68259), .B(n68258), .Y(n68912) );
  XNOR2X1 U71579 ( .A(n43666), .B(n39367), .Y(n68511) );
  INVX1 U71580 ( .A(n68804), .Y(n68808) );
  NOR2X1 U71581 ( .A(n43536), .B(n68260), .Y(n68261) );
  NOR2X1 U71582 ( .A(n68264), .B(n68263), .Y(n68266) );
  NOR2X1 U71583 ( .A(n68808), .B(n40106), .Y(n68270) );
  NAND2X1 U71584 ( .A(n43535), .B(n68804), .Y(n68268) );
  NAND2X1 U71585 ( .A(n68268), .B(n68267), .Y(n68269) );
  NAND2X1 U71586 ( .A(n68273), .B(n68271), .Y(n68599) );
  NOR2X1 U71587 ( .A(n68272), .B(n68599), .Y(n68275) );
  INVX1 U71588 ( .A(n68273), .Y(n68274) );
  NAND2X1 U71589 ( .A(n43581), .B(n68276), .Y(n68600) );
  XNOR2X1 U71590 ( .A(n68793), .B(n43580), .Y(n68490) );
  NOR2X1 U71591 ( .A(n41402), .B(n41412), .Y(n68280) );
  NAND2X1 U71592 ( .A(n39512), .B(n68279), .Y(n68782) );
  NAND2X1 U71593 ( .A(n68280), .B(n68782), .Y(n68597) );
  INVX1 U71594 ( .A(n68281), .Y(n68293) );
  INVX1 U71595 ( .A(n68282), .Y(n68287) );
  INVX1 U71596 ( .A(n68283), .Y(n68285) );
  NOR2X1 U71597 ( .A(n68285), .B(n68284), .Y(n68286) );
  NOR2X1 U71598 ( .A(n68287), .B(n68286), .Y(n68291) );
  NOR2X1 U71599 ( .A(n68289), .B(n68288), .Y(n68290) );
  NOR2X1 U71600 ( .A(n68291), .B(n68290), .Y(n68292) );
  NOR2X1 U71601 ( .A(n68293), .B(n68292), .Y(n68304) );
  INVX1 U71602 ( .A(n68744), .Y(n68447) );
  XNOR2X1 U71603 ( .A(n68446), .B(n68447), .Y(n68299) );
  INVX1 U71604 ( .A(n68740), .Y(n68297) );
  NAND2X1 U71605 ( .A(n68295), .B(n68294), .Y(n68296) );
  NOR2X1 U71606 ( .A(n68297), .B(n68296), .Y(n68298) );
  XNOR2X1 U71607 ( .A(n68299), .B(n68298), .Y(n68318) );
  INVX1 U71608 ( .A(n68318), .Y(n68308) );
  INVX1 U71609 ( .A(n68314), .Y(n68319) );
  XNOR2X1 U71610 ( .A(n39128), .B(n68319), .Y(n68302) );
  XNOR2X1 U71611 ( .A(n68308), .B(n68302), .Y(n68303) );
  XNOR2X1 U71612 ( .A(n39128), .B(n68305), .Y(n68307) );
  NAND2X1 U71613 ( .A(n68307), .B(n68306), .Y(n68761) );
  NAND2X1 U71614 ( .A(n68760), .B(n68761), .Y(n68457) );
  NOR2X1 U71615 ( .A(n39566), .B(n68308), .Y(n68317) );
  NOR2X1 U71616 ( .A(n68310), .B(n68309), .Y(n68312) );
  NOR2X1 U71617 ( .A(n68312), .B(n68311), .Y(n68313) );
  NOR2X1 U71618 ( .A(n37387), .B(n68313), .Y(n68315) );
  NOR2X1 U71619 ( .A(n68315), .B(n68314), .Y(n68316) );
  NAND2X1 U71620 ( .A(n43483), .B(n44000), .Y(n68699) );
  NAND2X1 U71621 ( .A(n68683), .B(n68320), .Y(n68331) );
  NAND2X1 U71622 ( .A(n68322), .B(n68321), .Y(n68323) );
  NOR2X1 U71623 ( .A(n68324), .B(n68323), .Y(n68326) );
  NOR2X1 U71624 ( .A(n68326), .B(n68325), .Y(n68327) );
  NOR2X1 U71625 ( .A(n39332), .B(n68327), .Y(n68329) );
  INVX1 U71626 ( .A(n68683), .Y(n68328) );
  NAND2X1 U71627 ( .A(n68329), .B(n68328), .Y(n68681) );
  NAND2X1 U71628 ( .A(n41523), .B(n68681), .Y(n68330) );
  NAND2X1 U71629 ( .A(n68331), .B(n68330), .Y(n68691) );
  INVX1 U71630 ( .A(n68691), .Y(n68697) );
  XNOR2X1 U71631 ( .A(n68699), .B(n68697), .Y(n68414) );
  NAND2X1 U71632 ( .A(n43491), .B(n43983), .Y(n69041) );
  XNOR2X1 U71633 ( .A(n68379), .B(n41716), .Y(n68332) );
  XNOR2X1 U71634 ( .A(n68333), .B(n68332), .Y(n68638) );
  INVX1 U71635 ( .A(n68638), .Y(n68335) );
  NOR2X1 U71636 ( .A(n68335), .B(n68334), .Y(n68337) );
  NOR2X1 U71637 ( .A(n68335), .B(n68636), .Y(n68336) );
  NOR2X1 U71638 ( .A(n68337), .B(n68336), .Y(n68350) );
  INVX1 U71639 ( .A(n68631), .Y(n68349) );
  NOR2X1 U71640 ( .A(n38481), .B(n68638), .Y(n68348) );
  NOR2X1 U71641 ( .A(n68342), .B(n68338), .Y(n68346) );
  NAND2X1 U71642 ( .A(n68340), .B(n68339), .Y(n68344) );
  OR2X1 U71643 ( .A(n68342), .B(n68341), .Y(n68343) );
  NAND2X1 U71644 ( .A(n68344), .B(n68343), .Y(n68345) );
  NOR2X1 U71645 ( .A(n68346), .B(n68345), .Y(n68347) );
  NAND2X1 U71646 ( .A(n68348), .B(n68347), .Y(n68629) );
  NAND2X1 U71647 ( .A(n68349), .B(n68629), .Y(n69055) );
  NAND2X1 U71648 ( .A(n43942), .B(n43500), .Y(n69127) );
  NAND2X1 U71649 ( .A(n68351), .B(n68358), .Y(n68667) );
  INVX1 U71650 ( .A(n68352), .Y(n68356) );
  NOR2X1 U71651 ( .A(n68354), .B(n68353), .Y(n68355) );
  NOR2X1 U71652 ( .A(n68356), .B(n68355), .Y(n68361) );
  INVX1 U71653 ( .A(n68357), .Y(n68359) );
  NOR2X1 U71654 ( .A(n68359), .B(n68358), .Y(n68360) );
  NAND2X1 U71655 ( .A(n68361), .B(n68360), .Y(n68665) );
  NAND2X1 U71656 ( .A(n41515), .B(n68665), .Y(n68362) );
  NAND2X1 U71657 ( .A(n68667), .B(n68362), .Y(n69094) );
  NAND2X1 U71658 ( .A(n72401), .B(n41686), .Y(n68363) );
  NAND2X1 U71659 ( .A(n41510), .B(n68363), .Y(n68366) );
  NAND2X1 U71660 ( .A(n41510), .B(n68364), .Y(n68365) );
  NAND2X1 U71661 ( .A(n68366), .B(n68365), .Y(n68648) );
  NAND2X1 U71662 ( .A(n43927), .B(n43608), .Y(n68646) );
  NAND2X1 U71663 ( .A(n41510), .B(n43604), .Y(n72296) );
  XNOR2X1 U71664 ( .A(n72296), .B(n68650), .Y(n68376) );
  OR2X1 U71665 ( .A(n72302), .B(n68367), .Y(n68368) );
  NOR2X1 U71666 ( .A(n72400), .B(n68368), .Y(n68375) );
  NOR2X1 U71667 ( .A(n72303), .B(n72400), .Y(n68370) );
  NAND2X1 U71668 ( .A(n72303), .B(n72400), .Y(n68371) );
  NOR2X1 U71669 ( .A(n72310), .B(n68371), .Y(n68369) );
  NOR2X1 U71670 ( .A(n68370), .B(n68369), .Y(n68373) );
  OR2X1 U71671 ( .A(n68653), .B(n68371), .Y(n68372) );
  NAND2X1 U71672 ( .A(n68373), .B(n68372), .Y(n68374) );
  NOR2X1 U71673 ( .A(n68375), .B(n68374), .Y(n68649) );
  NAND2X1 U71674 ( .A(n72397), .B(n68377), .Y(n71857) );
  NAND2X1 U71675 ( .A(n68650), .B(n72400), .Y(n71855) );
  NAND2X1 U71676 ( .A(n71855), .B(n72396), .Y(n68378) );
  NAND2X1 U71677 ( .A(n71857), .B(n68378), .Y(n68651) );
  NAND2X1 U71678 ( .A(n43933), .B(n39844), .Y(n69096) );
  INVX1 U71679 ( .A(n68644), .Y(n69128) );
  XNOR2X1 U71680 ( .A(n69127), .B(n69128), .Y(n68392) );
  INVX1 U71681 ( .A(n68379), .Y(n68389) );
  NOR2X1 U71682 ( .A(n68382), .B(n68381), .Y(n68380) );
  NOR2X1 U71683 ( .A(n68389), .B(n68380), .Y(n68386) );
  NAND2X1 U71684 ( .A(n68382), .B(n68381), .Y(n68384) );
  NAND2X1 U71685 ( .A(n68384), .B(n68383), .Y(n68385) );
  NAND2X1 U71686 ( .A(n68386), .B(n68385), .Y(n68387) );
  NAND2X1 U71687 ( .A(n41716), .B(n68387), .Y(n68391) );
  NAND2X1 U71688 ( .A(n68389), .B(n68388), .Y(n68390) );
  NAND2X1 U71689 ( .A(n68391), .B(n68390), .Y(n68643) );
  INVX1 U71690 ( .A(n68643), .Y(n69126) );
  XNOR2X1 U71691 ( .A(n68392), .B(n69126), .Y(n69057) );
  NAND2X1 U71692 ( .A(n43972), .B(n43496), .Y(n69067) );
  INVX1 U71693 ( .A(n69067), .Y(n68634) );
  XNOR2X1 U71694 ( .A(n69057), .B(n68634), .Y(n68393) );
  XNOR2X1 U71695 ( .A(n41005), .B(n68393), .Y(n69044) );
  INVX1 U71696 ( .A(n69044), .Y(n68627) );
  XNOR2X1 U71697 ( .A(n69041), .B(n68627), .Y(n68413) );
  NAND2X1 U71698 ( .A(n43991), .B(n43487), .Y(n68682) );
  NAND2X1 U71699 ( .A(n68395), .B(n68394), .Y(n69039) );
  INVX1 U71700 ( .A(n68396), .Y(n68408) );
  NOR2X1 U71701 ( .A(n68408), .B(n68397), .Y(n68406) );
  INVX1 U71702 ( .A(n68398), .Y(n68399) );
  NAND2X1 U71703 ( .A(n68636), .B(n68399), .Y(n68400) );
  NOR2X1 U71704 ( .A(n39466), .B(n68400), .Y(n68404) );
  NAND2X1 U71705 ( .A(n68402), .B(n68401), .Y(n68403) );
  NOR2X1 U71706 ( .A(n68404), .B(n68403), .Y(n68405) );
  NOR2X1 U71707 ( .A(n68406), .B(n68405), .Y(n68411) );
  NOR2X1 U71708 ( .A(n68408), .B(n68407), .Y(n68409) );
  NOR2X1 U71709 ( .A(n41003), .B(n68409), .Y(n68410) );
  NAND2X1 U71710 ( .A(n69039), .B(n69040), .Y(n68687) );
  XNOR2X1 U71711 ( .A(n68682), .B(n68687), .Y(n68412) );
  XNOR2X1 U71712 ( .A(n68413), .B(n68412), .Y(n68696) );
  XNOR2X1 U71713 ( .A(n68414), .B(n68696), .Y(n68615) );
  NAND2X1 U71714 ( .A(n43774), .B(n44017), .Y(n68619) );
  XNOR2X1 U71715 ( .A(n68619), .B(n42026), .Y(n68415) );
  XNOR2X1 U71716 ( .A(n68615), .B(n68415), .Y(n68426) );
  NAND2X1 U71717 ( .A(n68417), .B(n68416), .Y(n68418) );
  NAND2X1 U71718 ( .A(n68418), .B(n68427), .Y(n68700) );
  NOR2X1 U71719 ( .A(n37368), .B(n68418), .Y(n68423) );
  NAND2X1 U71720 ( .A(n41207), .B(n68419), .Y(n68420) );
  NAND2X1 U71721 ( .A(n68421), .B(n68420), .Y(n68422) );
  NAND2X1 U71722 ( .A(n68423), .B(n68422), .Y(n68424) );
  NAND2X1 U71723 ( .A(n68425), .B(n68424), .Y(n68702) );
  NAND2X1 U71724 ( .A(n68700), .B(n68702), .Y(n68698) );
  XNOR2X1 U71725 ( .A(n68426), .B(n39025), .Y(n68434) );
  NAND2X1 U71726 ( .A(n68710), .B(n68429), .Y(n68707) );
  INVX1 U71727 ( .A(n68430), .Y(n68715) );
  NAND2X1 U71728 ( .A(n68712), .B(n68709), .Y(n68431) );
  OR2X1 U71729 ( .A(n68710), .B(n68431), .Y(n68432) );
  NAND2X1 U71730 ( .A(n68715), .B(n68432), .Y(n68433) );
  NAND2X1 U71731 ( .A(n68707), .B(n68433), .Y(n68706) );
  INVX1 U71732 ( .A(n68706), .Y(n68617) );
  XNOR2X1 U71733 ( .A(n68434), .B(n68617), .Y(n68439) );
  NAND2X1 U71734 ( .A(n38954), .B(n68436), .Y(n68437) );
  NAND2X1 U71735 ( .A(n42034), .B(n68437), .Y(n68438) );
  NAND2X1 U71736 ( .A(n68621), .B(n68622), .Y(n68620) );
  NAND2X1 U71737 ( .A(n68438), .B(n68620), .Y(n68618) );
  INVX1 U71738 ( .A(n68726), .Y(n68978) );
  NAND2X1 U71739 ( .A(n43795), .B(n44025), .Y(n68725) );
  INVX1 U71740 ( .A(n68725), .Y(n68970) );
  NAND2X1 U71741 ( .A(n68441), .B(n68440), .Y(n68719) );
  NAND2X1 U71742 ( .A(n68719), .B(n68720), .Y(n68977) );
  XNOR2X1 U71743 ( .A(n41118), .B(n38986), .Y(n68753) );
  NAND2X1 U71744 ( .A(n68445), .B(n68743), .Y(n68751) );
  NAND2X1 U71745 ( .A(n42712), .B(n44048), .Y(n68448) );
  NAND2X1 U71746 ( .A(n40308), .B(n68446), .Y(n68449) );
  NAND2X1 U71747 ( .A(n68447), .B(n68449), .Y(n68750) );
  INVX1 U71748 ( .A(n68751), .Y(n68747) );
  INVX1 U71749 ( .A(n68448), .Y(n68749) );
  NOR2X1 U71750 ( .A(n68744), .B(n68448), .Y(n68450) );
  NAND2X1 U71751 ( .A(n68450), .B(n68449), .Y(n68451) );
  NAND2X1 U71752 ( .A(n68452), .B(n68451), .Y(n68453) );
  NAND2X1 U71753 ( .A(n42657), .B(n44055), .Y(n68758) );
  XNOR2X1 U71754 ( .A(n43598), .B(n68758), .Y(n68455) );
  XOR2X1 U71755 ( .A(n68457), .B(n68456), .Y(n69150) );
  NAND2X1 U71756 ( .A(n68461), .B(n68460), .Y(n68462) );
  XNOR2X1 U71757 ( .A(n68462), .B(n43618), .Y(n68463) );
  XNOR2X1 U71758 ( .A(n69150), .B(n68463), .Y(n68476) );
  NOR2X1 U71759 ( .A(n43617), .B(n68465), .Y(n68466) );
  NOR2X1 U71760 ( .A(n68467), .B(n68466), .Y(n68470) );
  NAND2X1 U71761 ( .A(n40027), .B(n68468), .Y(n68469) );
  NAND2X1 U71762 ( .A(n68470), .B(n68469), .Y(n68471) );
  NOR2X1 U71763 ( .A(n68482), .B(n68471), .Y(n68475) );
  NOR2X1 U71764 ( .A(n42996), .B(n68471), .Y(n68473) );
  NOR2X1 U71765 ( .A(n68482), .B(n42997), .Y(n68472) );
  OR2X1 U71766 ( .A(n68473), .B(n68472), .Y(n68474) );
  NOR2X1 U71767 ( .A(n68475), .B(n68474), .Y(n68780) );
  XNOR2X1 U71768 ( .A(n68780), .B(n68476), .Y(n68932) );
  INVX1 U71769 ( .A(n68477), .Y(n68478) );
  NAND2X1 U71770 ( .A(n43593), .B(n68478), .Y(n68486) );
  INVX1 U71771 ( .A(n68486), .Y(n68480) );
  NOR2X1 U71772 ( .A(n68480), .B(n68025), .Y(n68481) );
  NOR2X1 U71773 ( .A(n68481), .B(n42994), .Y(n68485) );
  NOR2X1 U71774 ( .A(n41620), .B(n42993), .Y(n68484) );
  NOR2X1 U71775 ( .A(n68485), .B(n68484), .Y(n68489) );
  NOR2X1 U71776 ( .A(n41622), .B(n41620), .Y(n68488) );
  NAND2X1 U71777 ( .A(n68487), .B(n68486), .Y(n68605) );
  NAND2X1 U71778 ( .A(n68488), .B(n68605), .Y(n68607) );
  NAND2X1 U71779 ( .A(n68489), .B(n68607), .Y(n68934) );
  XNOR2X1 U71780 ( .A(n43583), .B(n43569), .Y(n70272) );
  XNOR2X1 U71781 ( .A(n68490), .B(n68794), .Y(n68802) );
  NAND2X1 U71782 ( .A(n43580), .B(n68491), .Y(n69173) );
  NAND2X1 U71783 ( .A(n39646), .B(n69174), .Y(n68492) );
  NAND2X1 U71784 ( .A(n69173), .B(n68492), .Y(n68792) );
  XNOR2X1 U71785 ( .A(n68792), .B(n43537), .Y(n68493) );
  XNOR2X1 U71786 ( .A(n68802), .B(n68493), .Y(n68494) );
  INVX1 U71787 ( .A(n68590), .Y(n68593) );
  NOR2X1 U71788 ( .A(n39629), .B(n68495), .Y(n68499) );
  NOR2X1 U71789 ( .A(n68497), .B(n68496), .Y(n68498) );
  NAND2X1 U71790 ( .A(n68499), .B(n68498), .Y(n68500) );
  NOR2X1 U71791 ( .A(n68588), .B(n68500), .Y(n68503) );
  NAND2X1 U71792 ( .A(n68583), .B(n68501), .Y(n68505) );
  NOR2X1 U71793 ( .A(n68503), .B(n68502), .Y(n68504) );
  XNOR2X1 U71794 ( .A(n68593), .B(n68504), .Y(n68921) );
  XNOR2X1 U71795 ( .A(n68921), .B(n72587), .Y(n68510) );
  XNOR2X1 U71796 ( .A(n40093), .B(n43564), .Y(n68506) );
  NOR2X1 U71797 ( .A(n68570), .B(n43627), .Y(n68508) );
  INVX1 U71798 ( .A(n68570), .Y(n68575) );
  NOR2X1 U71799 ( .A(n43620), .B(n68575), .Y(n68509) );
  XNOR2X1 U71800 ( .A(n41025), .B(n68510), .Y(n68553) );
  XNOR2X1 U71801 ( .A(n68555), .B(n68512), .Y(n68549) );
  XNOR2X1 U71802 ( .A(n68549), .B(n43643), .Y(n68513) );
  XNOR2X1 U71803 ( .A(n41072), .B(n68513), .Y(n68819) );
  XNOR2X1 U71804 ( .A(n43661), .B(n68819), .Y(n68514) );
  XOR2X1 U71805 ( .A(n68818), .B(n68514), .Y(n68826) );
  XNOR2X1 U71806 ( .A(n41036), .B(n68516), .Y(n68517) );
  XNOR2X1 U71807 ( .A(n68825), .B(n43523), .Y(n68518) );
  XNOR2X1 U71808 ( .A(n68826), .B(n68518), .Y(n68829) );
  XNOR2X1 U71809 ( .A(n68829), .B(n43679), .Y(n68519) );
  XNOR2X1 U71810 ( .A(n39841), .B(n68519), .Y(n68520) );
  XNOR2X1 U71811 ( .A(n36445), .B(n43508), .Y(n68526) );
  XNOR2X1 U71812 ( .A(n68521), .B(n43523), .Y(n68522) );
  XNOR2X1 U71813 ( .A(n38047), .B(n68522), .Y(n68523) );
  XNOR2X1 U71814 ( .A(n68523), .B(n39973), .Y(n68524) );
  XNOR2X1 U71815 ( .A(n41095), .B(n68524), .Y(n68838) );
  NOR2X1 U71816 ( .A(n38055), .B(n41431), .Y(n68525) );
  XNOR2X1 U71817 ( .A(n68526), .B(n68525), .Y(n68545) );
  XNOR2X1 U71818 ( .A(n43697), .B(n68545), .Y(n68527) );
  XNOR2X1 U71819 ( .A(n68528), .B(n68527), .Y(n68537) );
  XNOR2X1 U71820 ( .A(n68533), .B(n68532), .Y(n68534) );
  XNOR2X1 U71821 ( .A(n42049), .B(n68534), .Y(n68535) );
  MX2X1 U71822 ( .A(n68536), .B(n68535), .S0(n43719), .Y(u_muldiv_result_r[19]) );
  NAND2X1 U71823 ( .A(u_muldiv_mult_result_q[19]), .B(n44632), .Y(n13959) );
  NAND2X1 U71824 ( .A(n37955), .B(n40456), .Y(n68855) );
  NAND2X1 U71825 ( .A(n68855), .B(n37967), .Y(n68538) );
  NAND2X1 U71826 ( .A(n43705), .B(n68537), .Y(n68854) );
  NAND2X1 U71827 ( .A(n68538), .B(n68854), .Y(n68848) );
  NAND2X1 U71828 ( .A(n68540), .B(n68539), .Y(n69225) );
  NAND2X1 U71829 ( .A(n67919), .B(n43697), .Y(n68542) );
  NAND2X1 U71830 ( .A(n68542), .B(n68541), .Y(n68543) );
  NOR2X1 U71831 ( .A(n41415), .B(n68543), .Y(n68548) );
  NAND2X1 U71832 ( .A(n68547), .B(n68546), .Y(n69231) );
  NAND2X1 U71833 ( .A(n69251), .B(n69247), .Y(n68818) );
  NAND2X1 U71834 ( .A(n38694), .B(n43647), .Y(n68550) );
  NAND2X1 U71835 ( .A(n68550), .B(n68818), .Y(n68552) );
  NAND2X1 U71836 ( .A(n43642), .B(n68551), .Y(n69250) );
  AND2X1 U71837 ( .A(n68552), .B(n69250), .Y(n68881) );
  XNOR2X1 U71838 ( .A(n68553), .B(n39367), .Y(n68554) );
  INVX1 U71839 ( .A(n68557), .Y(n68556) );
  NAND2X1 U71840 ( .A(n43665), .B(n68556), .Y(n69529) );
  NAND2X1 U71841 ( .A(n68559), .B(n68558), .Y(n68892) );
  NAND2X1 U71842 ( .A(n68892), .B(n38365), .Y(n69528) );
  INVX1 U71843 ( .A(n68921), .Y(n69268) );
  XNOR2X1 U71844 ( .A(n41025), .B(n69268), .Y(n68563) );
  NAND2X1 U71845 ( .A(n68563), .B(n43636), .Y(n68561) );
  NAND2X1 U71846 ( .A(n68561), .B(n68560), .Y(n69515) );
  NAND2X1 U71847 ( .A(n69516), .B(n69515), .Y(n69209) );
  XNOR2X1 U71848 ( .A(n39919), .B(n43643), .Y(n68815) );
  NOR2X1 U71849 ( .A(n43545), .B(n39391), .Y(n68565) );
  NOR2X1 U71850 ( .A(n68563), .B(n68562), .Y(n68564) );
  NOR2X1 U71851 ( .A(n36735), .B(n43552), .Y(n68569) );
  NAND2X1 U71852 ( .A(n68567), .B(n68566), .Y(n68568) );
  NAND2X1 U71853 ( .A(n43544), .B(n68568), .Y(n68910) );
  NAND2X1 U71854 ( .A(n43619), .B(n68570), .Y(n68914) );
  NOR2X1 U71855 ( .A(n68572), .B(n43627), .Y(n68574) );
  NAND2X1 U71856 ( .A(n68575), .B(n43626), .Y(n68576) );
  NAND2X1 U71857 ( .A(n68916), .B(n68576), .Y(n68920) );
  NAND2X1 U71858 ( .A(n68914), .B(n68920), .Y(n68578) );
  NAND2X1 U71859 ( .A(n43619), .B(n36678), .Y(n68577) );
  NOR2X1 U71860 ( .A(n68578), .B(n68577), .Y(n68581) );
  NAND2X1 U71861 ( .A(n68921), .B(n43625), .Y(n68579) );
  NOR2X1 U71862 ( .A(n39004), .B(n68579), .Y(n68580) );
  NOR2X1 U71863 ( .A(n68585), .B(n68584), .Y(n68586) );
  NOR2X1 U71864 ( .A(n43563), .B(n68586), .Y(n68587) );
  NOR2X1 U71865 ( .A(n36674), .B(n68587), .Y(n68589) );
  NOR2X1 U71866 ( .A(n68590), .B(n43560), .Y(n68591) );
  NOR2X1 U71867 ( .A(n68592), .B(n68591), .Y(n68596) );
  NAND2X1 U71868 ( .A(n68594), .B(n68593), .Y(n68595) );
  NAND2X1 U71869 ( .A(n68595), .B(n38424), .Y(n69191) );
  XNOR2X1 U71870 ( .A(n69191), .B(n43565), .Y(n68813) );
  XNOR2X1 U71871 ( .A(n68785), .B(n43569), .Y(n68598) );
  NAND2X1 U71872 ( .A(n68599), .B(n68600), .Y(n68601) );
  NAND2X1 U71873 ( .A(n43581), .B(n68601), .Y(n69163) );
  NAND2X1 U71874 ( .A(n68602), .B(n68793), .Y(n69165) );
  NAND2X1 U71875 ( .A(n69163), .B(n69165), .Y(n68603) );
  NOR2X1 U71876 ( .A(n38144), .B(n68603), .Y(n68791) );
  NAND2X1 U71877 ( .A(n41620), .B(n43593), .Y(n68604) );
  NOR2X1 U71878 ( .A(n68605), .B(n68604), .Y(n68606) );
  INVX1 U71879 ( .A(n68932), .Y(n68933) );
  NAND2X1 U71880 ( .A(n68606), .B(n68933), .Y(n68609) );
  NAND2X1 U71881 ( .A(n68609), .B(n68608), .Y(n68610) );
  XNOR2X1 U71882 ( .A(n68610), .B(n43569), .Y(n68781) );
  NOR2X1 U71883 ( .A(n39570), .B(n68758), .Y(n68612) );
  NOR2X1 U71884 ( .A(n40191), .B(n68758), .Y(n68611) );
  NOR2X1 U71885 ( .A(n68612), .B(n68611), .Y(n68614) );
  NAND2X1 U71886 ( .A(n68759), .B(n39159), .Y(n68613) );
  NAND2X1 U71887 ( .A(n68614), .B(n68613), .Y(n68961) );
  XNOR2X1 U71888 ( .A(n68705), .B(n42026), .Y(n68616) );
  XNOR2X1 U71889 ( .A(n68617), .B(n68616), .Y(n68624) );
  NAND2X1 U71890 ( .A(n68624), .B(n68618), .Y(n69449) );
  NOR2X1 U71891 ( .A(n68622), .B(n68621), .Y(n68623) );
  INVX1 U71892 ( .A(n68624), .Y(n68625) );
  NAND2X1 U71893 ( .A(n69449), .B(n69448), .Y(n68986) );
  NAND2X1 U71894 ( .A(n69044), .B(n39237), .Y(n69015) );
  INVX1 U71895 ( .A(n69041), .Y(n69045) );
  INVX1 U71896 ( .A(n39237), .Y(n68628) );
  NAND2X1 U71897 ( .A(n68628), .B(n68627), .Y(n69017) );
  NAND2X1 U71898 ( .A(n69045), .B(n69017), .Y(n69012) );
  NAND2X1 U71899 ( .A(n69015), .B(n69012), .Y(n69037) );
  NAND2X1 U71900 ( .A(n68634), .B(n68629), .Y(n68630) );
  NOR2X1 U71901 ( .A(n68631), .B(n68630), .Y(n68633) );
  NOR2X1 U71902 ( .A(n41005), .B(n69057), .Y(n68632) );
  NOR2X1 U71903 ( .A(n68633), .B(n68632), .Y(n68642) );
  NAND2X1 U71904 ( .A(n68635), .B(n43934), .Y(n68637) );
  NAND2X1 U71905 ( .A(n68637), .B(n68636), .Y(n68639) );
  NAND2X1 U71906 ( .A(n68639), .B(n68638), .Y(n69056) );
  NOR2X1 U71907 ( .A(n69067), .B(n69056), .Y(n68640) );
  NOR2X1 U71908 ( .A(n41250), .B(n68640), .Y(n68641) );
  NAND2X1 U71909 ( .A(n68642), .B(n68641), .Y(n69053) );
  NAND2X1 U71910 ( .A(n68644), .B(n68643), .Y(n69125) );
  NAND2X1 U71911 ( .A(n69125), .B(n68645), .Y(n69124) );
  INVX1 U71912 ( .A(n68646), .Y(n68657) );
  NAND2X1 U71913 ( .A(n68657), .B(n68647), .Y(n69084) );
  NAND2X1 U71914 ( .A(n68657), .B(n68648), .Y(n69087) );
  NAND2X1 U71915 ( .A(n69084), .B(n69087), .Y(n69082) );
  INVX1 U71916 ( .A(n72296), .Y(n72327) );
  XNOR2X1 U71917 ( .A(n68650), .B(n68649), .Y(n69343) );
  INVX1 U71918 ( .A(n69343), .Y(n69339) );
  XNOR2X1 U71919 ( .A(n72327), .B(n69339), .Y(n69080) );
  NAND2X1 U71920 ( .A(n72327), .B(n69339), .Y(n69107) );
  NAND2X1 U71921 ( .A(n69343), .B(n72296), .Y(n69109) );
  NAND2X1 U71922 ( .A(n69109), .B(n68651), .Y(n68652) );
  NAND2X1 U71923 ( .A(n69107), .B(n68652), .Y(n69118) );
  INVX1 U71924 ( .A(n69118), .Y(n69078) );
  XNOR2X1 U71925 ( .A(n69080), .B(n69078), .Y(n68659) );
  NAND2X1 U71926 ( .A(n68654), .B(n68653), .Y(n68655) );
  NAND2X1 U71927 ( .A(n72303), .B(n68655), .Y(n69105) );
  NAND2X1 U71928 ( .A(n69105), .B(n71857), .Y(n68656) );
  NAND2X1 U71929 ( .A(n68656), .B(n71855), .Y(n69108) );
  NAND2X1 U71930 ( .A(n43933), .B(n43608), .Y(n69120) );
  INVX1 U71931 ( .A(n69120), .Y(n69106) );
  NAND2X1 U71932 ( .A(n68657), .B(n43604), .Y(n72288) );
  INVX1 U71933 ( .A(n72288), .Y(n72291) );
  XNOR2X1 U71934 ( .A(n69106), .B(n72291), .Y(n69079) );
  XNOR2X1 U71935 ( .A(n69108), .B(n69079), .Y(n68658) );
  XNOR2X1 U71936 ( .A(n68659), .B(n68658), .Y(n68660) );
  INVX1 U71937 ( .A(n69093), .Y(n68661) );
  NAND2X1 U71938 ( .A(n68661), .B(n69094), .Y(n69074) );
  INVX1 U71939 ( .A(n69074), .Y(n69092) );
  NAND2X1 U71940 ( .A(n43942), .B(n43518), .Y(n68671) );
  INVX1 U71941 ( .A(n68671), .Y(n69102) );
  NOR2X1 U71942 ( .A(n69102), .B(n43936), .Y(n68662) );
  NOR2X1 U71943 ( .A(n69092), .B(n68662), .Y(n68664) );
  NOR2X1 U71944 ( .A(n69102), .B(n69074), .Y(n68663) );
  NOR2X1 U71945 ( .A(n68664), .B(n68663), .Y(n68670) );
  NAND2X1 U71946 ( .A(n68665), .B(n43928), .Y(n68666) );
  NOR2X1 U71947 ( .A(n36706), .B(n68668), .Y(n69073) );
  NOR2X1 U71948 ( .A(n69102), .B(n69073), .Y(n68669) );
  NOR2X1 U71949 ( .A(n68670), .B(n68669), .Y(n68674) );
  NOR2X1 U71950 ( .A(n43938), .B(n68671), .Y(n68672) );
  NAND2X1 U71951 ( .A(n69073), .B(n68672), .Y(n68673) );
  NAND2X1 U71952 ( .A(n68674), .B(n68673), .Y(n69062) );
  XNOR2X1 U71953 ( .A(n69124), .B(n41683), .Y(n68675) );
  NAND2X1 U71954 ( .A(n43972), .B(n43500), .Y(n69060) );
  INVX1 U71955 ( .A(n69060), .Y(n69133) );
  XNOR2X1 U71956 ( .A(n68675), .B(n69133), .Y(n69054) );
  INVX1 U71957 ( .A(n69054), .Y(n68678) );
  NAND2X1 U71958 ( .A(n43491), .B(n43992), .Y(n69016) );
  NAND2X1 U71959 ( .A(n43982), .B(n43497), .Y(n69380) );
  INVX1 U71960 ( .A(n69380), .Y(n69071) );
  XNOR2X1 U71961 ( .A(n69016), .B(n69071), .Y(n68676) );
  XNOR2X1 U71962 ( .A(n69400), .B(n68676), .Y(n68677) );
  XNOR2X1 U71963 ( .A(n68678), .B(n68677), .Y(n68679) );
  XNOR2X1 U71964 ( .A(n69053), .B(n68679), .Y(n68680) );
  NAND2X1 U71965 ( .A(n43482), .B(n44008), .Y(n69424) );
  INVX1 U71966 ( .A(n69424), .Y(n69421) );
  XNOR2X1 U71967 ( .A(n41724), .B(n69421), .Y(n68694) );
  INVX1 U71968 ( .A(n68682), .Y(n68688) );
  NAND2X1 U71969 ( .A(n68688), .B(n68683), .Y(n68684) );
  NOR2X1 U71970 ( .A(n39396), .B(n68684), .Y(n68685) );
  NOR2X1 U71971 ( .A(n68686), .B(n68685), .Y(n68690) );
  NAND2X1 U71972 ( .A(n68688), .B(n68692), .Y(n68689) );
  NAND2X1 U71973 ( .A(n68690), .B(n68689), .Y(n69026) );
  INVX1 U71974 ( .A(n69026), .Y(n68693) );
  NAND2X1 U71975 ( .A(n68692), .B(n68691), .Y(n69024) );
  XNOR2X1 U71976 ( .A(n68694), .B(n37370), .Y(n68695) );
  XNOR2X1 U71977 ( .A(n69003), .B(n68695), .Y(n68704) );
  XNOR2X1 U71978 ( .A(n68697), .B(n68696), .Y(n68701) );
  NAND2X1 U71979 ( .A(n68701), .B(n68698), .Y(n69006) );
  NOR2X1 U71980 ( .A(n38951), .B(n68701), .Y(n68703) );
  NAND2X1 U71981 ( .A(n69006), .B(n69005), .Y(n69004) );
  INVX1 U71982 ( .A(n69004), .Y(n68995) );
  XNOR2X1 U71983 ( .A(n68704), .B(n68995), .Y(n68718) );
  INVX1 U71984 ( .A(n68705), .Y(n68708) );
  NAND2X1 U71985 ( .A(n68708), .B(n68706), .Y(n68999) );
  NOR2X1 U71986 ( .A(n38131), .B(n68708), .Y(n68717) );
  INVX1 U71987 ( .A(n68709), .Y(n68711) );
  NOR2X1 U71988 ( .A(n68711), .B(n68710), .Y(n68713) );
  NAND2X1 U71989 ( .A(n68713), .B(n68712), .Y(n68714) );
  NAND2X1 U71990 ( .A(n68715), .B(n68714), .Y(n68716) );
  NAND2X1 U71991 ( .A(n68717), .B(n68716), .Y(n68997) );
  NAND2X1 U71992 ( .A(n43774), .B(n44025), .Y(n69453) );
  INVX1 U71993 ( .A(n69453), .Y(n68991) );
  XNOR2X1 U71994 ( .A(n68964), .B(n41729), .Y(n68735) );
  NAND2X1 U71995 ( .A(n68720), .B(n68719), .Y(n68722) );
  NAND2X1 U71996 ( .A(n68970), .B(n68978), .Y(n68969) );
  NAND2X1 U71997 ( .A(n43796), .B(n44048), .Y(n68968) );
  NAND2X1 U71998 ( .A(n68969), .B(n68968), .Y(n68721) );
  NOR2X1 U71999 ( .A(n68722), .B(n68721), .Y(n68734) );
  INVX1 U72000 ( .A(n68968), .Y(n68979) );
  NAND2X1 U72001 ( .A(n68726), .B(n68725), .Y(n68723) );
  NAND2X1 U72002 ( .A(n68979), .B(n68723), .Y(n68724) );
  OR2X1 U72003 ( .A(n38986), .B(n68724), .Y(n68732) );
  OR2X1 U72004 ( .A(n68979), .B(n68725), .Y(n68730) );
  NAND2X1 U72005 ( .A(n68726), .B(n68968), .Y(n68728) );
  OR2X1 U72006 ( .A(n68726), .B(n68725), .Y(n68727) );
  NAND2X1 U72007 ( .A(n68728), .B(n68727), .Y(n68729) );
  NAND2X1 U72008 ( .A(n68730), .B(n68729), .Y(n68731) );
  NAND2X1 U72009 ( .A(n68732), .B(n68731), .Y(n68733) );
  NOR2X1 U72010 ( .A(n68734), .B(n68733), .Y(n68965) );
  XNOR2X1 U72011 ( .A(n68735), .B(n68965), .Y(n68959) );
  NOR2X1 U72012 ( .A(n68737), .B(n68736), .Y(n68741) );
  NAND2X1 U72013 ( .A(n68739), .B(n68738), .Y(n68740) );
  NAND2X1 U72014 ( .A(n68741), .B(n68740), .Y(n68742) );
  NOR2X1 U72015 ( .A(n68743), .B(n68742), .Y(n68745) );
  NOR2X1 U72016 ( .A(n68745), .B(n68744), .Y(n68746) );
  NAND2X1 U72017 ( .A(n68749), .B(n68748), .Y(n68755) );
  NAND2X1 U72018 ( .A(n40166), .B(n68750), .Y(n68752) );
  NAND2X1 U72019 ( .A(n68753), .B(n68752), .Y(n68754) );
  XNOR2X1 U72020 ( .A(n39521), .B(n42187), .Y(n68756) );
  XNOR2X1 U72021 ( .A(n68959), .B(n68756), .Y(n68757) );
  INVX1 U72022 ( .A(n69318), .Y(n69315) );
  NAND2X1 U72023 ( .A(n68761), .B(n68760), .Y(n69312) );
  NOR2X1 U72024 ( .A(n39342), .B(n39930), .Y(n68765) );
  NAND2X1 U72025 ( .A(n39930), .B(n43598), .Y(n68763) );
  NAND2X1 U72026 ( .A(n43599), .B(n69313), .Y(n68762) );
  NAND2X1 U72027 ( .A(n68763), .B(n68762), .Y(n68764) );
  NOR2X1 U72028 ( .A(n68765), .B(n68764), .Y(n68766) );
  XNOR2X1 U72029 ( .A(n69304), .B(n43618), .Y(n68778) );
  INVX1 U72030 ( .A(n68768), .Y(n68767) );
  NAND2X1 U72031 ( .A(n40683), .B(n68767), .Y(n68771) );
  NAND2X1 U72032 ( .A(n43615), .B(n68768), .Y(n68769) );
  NAND2X1 U72033 ( .A(n39731), .B(n68769), .Y(n68770) );
  NAND2X1 U72034 ( .A(n68771), .B(n68770), .Y(n69151) );
  INVX1 U72035 ( .A(n69151), .Y(n68773) );
  INVX1 U72036 ( .A(n69150), .Y(n69149) );
  NAND2X1 U72037 ( .A(n43615), .B(n69149), .Y(n68772) );
  NOR2X1 U72038 ( .A(n68773), .B(n68772), .Y(n68776) );
  NAND2X1 U72039 ( .A(n69150), .B(n40683), .Y(n68774) );
  NOR2X1 U72040 ( .A(n68774), .B(n69151), .Y(n68775) );
  NOR2X1 U72041 ( .A(n68776), .B(n68775), .Y(n68777) );
  XNOR2X1 U72042 ( .A(n68778), .B(n68777), .Y(n68939) );
  NAND2X1 U72043 ( .A(n69149), .B(n42997), .Y(n68945) );
  NAND2X1 U72044 ( .A(n43617), .B(n69150), .Y(n68779) );
  NAND2X1 U72045 ( .A(n68780), .B(n68779), .Y(n68947) );
  NAND2X1 U72046 ( .A(n68945), .B(n68947), .Y(n69305) );
  INVX1 U72047 ( .A(n69498), .Y(n69499) );
  XNOR2X1 U72048 ( .A(n68781), .B(n69499), .Y(n69164) );
  NOR2X1 U72049 ( .A(n41147), .B(n40670), .Y(n68784) );
  NOR2X1 U72050 ( .A(n68785), .B(n41147), .Y(n68783) );
  NOR2X1 U72051 ( .A(n68784), .B(n68783), .Y(n68788) );
  INVX1 U72052 ( .A(n68785), .Y(n68786) );
  NAND2X1 U72053 ( .A(n43567), .B(n68786), .Y(n68787) );
  NAND2X1 U72054 ( .A(n68788), .B(n68787), .Y(n69158) );
  XNOR2X1 U72055 ( .A(n69158), .B(n43583), .Y(n68789) );
  XNOR2X1 U72056 ( .A(n69164), .B(n68789), .Y(n68790) );
  XNOR2X1 U72057 ( .A(n68791), .B(n68790), .Y(n69288) );
  INVX1 U72058 ( .A(n69288), .Y(n69850) );
  INVX1 U72059 ( .A(n68792), .Y(n68803) );
  INVX1 U72060 ( .A(n69178), .Y(n69181) );
  NAND2X1 U72061 ( .A(n69181), .B(n39958), .Y(n68795) );
  NOR2X1 U72062 ( .A(n68803), .B(n68795), .Y(n68800) );
  NAND2X1 U72063 ( .A(n43576), .B(n69178), .Y(n68798) );
  NAND2X1 U72064 ( .A(n68796), .B(n69173), .Y(n68797) );
  NOR2X1 U72065 ( .A(n68798), .B(n68797), .Y(n68799) );
  NOR2X1 U72066 ( .A(n68800), .B(n68799), .Y(n68801) );
  XNOR2X1 U72067 ( .A(n69850), .B(n68801), .Y(n68927) );
  NOR2X1 U72068 ( .A(n40493), .B(n40093), .Y(n68805) );
  NOR2X1 U72069 ( .A(n68805), .B(n43542), .Y(n68806) );
  NOR2X1 U72070 ( .A(n68807), .B(n68806), .Y(n68812) );
  NOR2X1 U72071 ( .A(n68808), .B(n40106), .Y(n68810) );
  NAND2X1 U72072 ( .A(n68810), .B(n68809), .Y(n68811) );
  NAND2X1 U72073 ( .A(n68811), .B(n68812), .Y(n68928) );
  XNOR2X1 U72074 ( .A(n39187), .B(n68813), .Y(n68924) );
  INVX1 U72075 ( .A(n68924), .Y(n69276) );
  XNOR2X1 U72076 ( .A(n69207), .B(n69861), .Y(n68814) );
  XOR2X1 U72077 ( .A(n68905), .B(n68814), .Y(n68893) );
  XNOR2X1 U72078 ( .A(n40959), .B(n68816), .Y(n68880) );
  XNOR2X1 U72079 ( .A(n68880), .B(n43654), .Y(n68817) );
  XNOR2X1 U72080 ( .A(n68881), .B(n68817), .Y(n68872) );
  INVX1 U72081 ( .A(n68820), .Y(n68821) );
  XNOR2X1 U72082 ( .A(n43532), .B(n68871), .Y(n68822) );
  XOR2X1 U72083 ( .A(n68872), .B(n68822), .Y(n68858) );
  NOR2X1 U72084 ( .A(n43523), .B(n41060), .Y(n68828) );
  NOR2X1 U72085 ( .A(n43523), .B(n68873), .Y(n68827) );
  INVX1 U72086 ( .A(n68873), .Y(n68877) );
  XNOR2X1 U72087 ( .A(n43509), .B(n41124), .Y(n68836) );
  INVX1 U72088 ( .A(n68864), .Y(n69547) );
  NAND2X1 U72089 ( .A(n68861), .B(n68860), .Y(n68831) );
  NOR2X1 U72090 ( .A(n36523), .B(n68831), .Y(n68832) );
  NOR2X1 U72091 ( .A(n43678), .B(n68832), .Y(n68833) );
  INVX1 U72092 ( .A(n68868), .Y(n69218) );
  XNOR2X1 U72093 ( .A(n68836), .B(n69218), .Y(n68845) );
  NOR2X1 U72094 ( .A(n36445), .B(n41431), .Y(n68837) );
  NAND2X1 U72095 ( .A(n69220), .B(n68837), .Y(n69579) );
  NOR2X1 U72096 ( .A(n41204), .B(n68838), .Y(n68840) );
  NAND2X1 U72097 ( .A(n68840), .B(n68839), .Y(n68841) );
  NOR2X1 U72098 ( .A(n38061), .B(n68843), .Y(n68844) );
  XNOR2X1 U72099 ( .A(n68844), .B(n68845), .Y(n70187) );
  XNOR2X1 U72100 ( .A(n70187), .B(n43692), .Y(n68846) );
  XNOR2X1 U72101 ( .A(n41164), .B(n68846), .Y(n68856) );
  XNOR2X1 U72102 ( .A(n68856), .B(n43708), .Y(n68847) );
  XNOR2X1 U72103 ( .A(n68848), .B(n68847), .Y(n68853) );
  XNOR2X1 U72104 ( .A(n68850), .B(n68849), .Y(n68851) );
  XNOR2X1 U72105 ( .A(n42059), .B(n68851), .Y(n68852) );
  MX2X1 U72106 ( .A(n68853), .B(n68852), .S0(n43719), .Y(u_muldiv_result_r[20]) );
  NAND2X1 U72107 ( .A(u_muldiv_mult_result_q[20]), .B(n44632), .Y(n13951) );
  INVX1 U72108 ( .A(n68854), .Y(n69239) );
  INVX1 U72109 ( .A(n69546), .Y(n68859) );
  NOR2X1 U72110 ( .A(n43678), .B(n68859), .Y(n68867) );
  INVX1 U72111 ( .A(n68860), .Y(n68863) );
  INVX1 U72112 ( .A(n68861), .Y(n68862) );
  NAND2X1 U72113 ( .A(n69548), .B(n43682), .Y(n68865) );
  NAND2X1 U72114 ( .A(n68865), .B(n68864), .Y(n68866) );
  NOR2X1 U72115 ( .A(n68867), .B(n68866), .Y(n68870) );
  NAND2X1 U72116 ( .A(n69546), .B(n68868), .Y(n68869) );
  XNOR2X1 U72117 ( .A(n43509), .B(n41138), .Y(n69217) );
  NOR2X1 U72118 ( .A(n68877), .B(n43532), .Y(n68878) );
  INVX1 U72119 ( .A(n68891), .Y(n68882) );
  NAND2X1 U72120 ( .A(n68882), .B(n43658), .Y(n69243) );
  INVX1 U72121 ( .A(n68884), .Y(n68888) );
  NAND2X1 U72122 ( .A(n68886), .B(n68885), .Y(n68887) );
  NOR2X1 U72123 ( .A(n68888), .B(n68887), .Y(n68889) );
  NOR2X1 U72124 ( .A(n38945), .B(n68889), .Y(n68890) );
  NAND2X1 U72125 ( .A(n69243), .B(n36625), .Y(n69591) );
  XNOR2X1 U72126 ( .A(n43524), .B(n38605), .Y(n69215) );
  XNOR2X1 U72127 ( .A(n68893), .B(n39919), .Y(n68894) );
  NOR2X1 U72128 ( .A(n69255), .B(n43646), .Y(n68898) );
  NAND2X1 U72129 ( .A(n41036), .B(n68895), .Y(n69252) );
  NAND2X1 U72130 ( .A(n69252), .B(n43647), .Y(n68896) );
  NAND2X1 U72131 ( .A(n68550), .B(n68896), .Y(n68897) );
  NOR2X1 U72132 ( .A(n68898), .B(n68897), .Y(n68902) );
  INVX1 U72133 ( .A(n68818), .Y(n68899) );
  NAND2X1 U72134 ( .A(n68899), .B(n38694), .Y(n68900) );
  NAND2X1 U72135 ( .A(n69255), .B(n68900), .Y(n68901) );
  NAND2X1 U72136 ( .A(n68902), .B(n68901), .Y(n69536) );
  INVX1 U72137 ( .A(n68903), .Y(n68905) );
  XNOR2X1 U72138 ( .A(n69207), .B(n43633), .Y(n68904) );
  NAND2X1 U72139 ( .A(n68905), .B(n68904), .Y(n68906) );
  NAND2X1 U72140 ( .A(n68907), .B(n69527), .Y(n69865) );
  NAND2X1 U72141 ( .A(n68908), .B(n69863), .Y(n68909) );
  NOR2X1 U72142 ( .A(n39357), .B(n68909), .Y(n69213) );
  NAND2X1 U72143 ( .A(n43544), .B(n36735), .Y(n68911) );
  NAND2X1 U72144 ( .A(n36735), .B(n68912), .Y(n68913) );
  XNOR2X1 U72145 ( .A(n69513), .B(n43666), .Y(n69206) );
  NAND2X1 U72146 ( .A(n68924), .B(n43625), .Y(n68923) );
  NOR2X1 U72147 ( .A(n69268), .B(n43628), .Y(n68919) );
  INVX1 U72148 ( .A(n68914), .Y(n68915) );
  NOR2X1 U72149 ( .A(n68916), .B(n68915), .Y(n68917) );
  NOR2X1 U72150 ( .A(n68917), .B(n43627), .Y(n68918) );
  INVX1 U72151 ( .A(n68920), .Y(n68922) );
  NAND2X1 U72152 ( .A(n40186), .B(n43624), .Y(n69261) );
  NAND2X1 U72153 ( .A(n68923), .B(n69261), .Y(n68926) );
  INVX1 U72154 ( .A(n69260), .Y(n68925) );
  NAND2X1 U72155 ( .A(n68927), .B(n43539), .Y(n68931) );
  NAND2X1 U72156 ( .A(n43535), .B(n69288), .Y(n68929) );
  NAND2X1 U72157 ( .A(n39976), .B(n68929), .Y(n68930) );
  NAND2X1 U72158 ( .A(n68931), .B(n68930), .Y(n69620) );
  XNOR2X1 U72159 ( .A(n43621), .B(n72149), .Y(n69162) );
  NAND2X1 U72160 ( .A(n43593), .B(n68932), .Y(n68937) );
  NAND2X1 U72161 ( .A(n68933), .B(n42992), .Y(n68935) );
  NAND2X1 U72162 ( .A(n68935), .B(n68934), .Y(n68936) );
  NAND2X1 U72163 ( .A(n68937), .B(n68936), .Y(n68940) );
  INVX1 U72164 ( .A(n68940), .Y(n69500) );
  NOR2X1 U72165 ( .A(n69499), .B(n42994), .Y(n68938) );
  NAND2X1 U72166 ( .A(n69500), .B(n68938), .Y(n68943) );
  NOR2X1 U72167 ( .A(n43593), .B(n68939), .Y(n68941) );
  NAND2X1 U72168 ( .A(n68941), .B(n68940), .Y(n68942) );
  NAND2X1 U72169 ( .A(n68943), .B(n68942), .Y(n69157) );
  INVX1 U72170 ( .A(n69304), .Y(n69148) );
  NAND2X1 U72171 ( .A(n43617), .B(n69148), .Y(n68944) );
  NOR2X1 U72172 ( .A(n68944), .B(n68947), .Y(n68952) );
  NAND2X1 U72173 ( .A(n69148), .B(n42995), .Y(n69307) );
  INVX1 U72174 ( .A(n69307), .Y(n68950) );
  INVX1 U72175 ( .A(n68945), .Y(n68946) );
  NOR2X1 U72176 ( .A(n43617), .B(n68946), .Y(n68948) );
  NAND2X1 U72177 ( .A(n68948), .B(n68947), .Y(n68949) );
  NOR2X1 U72178 ( .A(n68950), .B(n68949), .Y(n68951) );
  NAND2X1 U72179 ( .A(n39930), .B(n68762), .Y(n69317) );
  INVX1 U72180 ( .A(n69317), .Y(n68955) );
  NAND2X1 U72181 ( .A(n39342), .B(n43598), .Y(n68953) );
  NOR2X1 U72182 ( .A(n68955), .B(n68953), .Y(n68954) );
  NAND2X1 U72183 ( .A(n68954), .B(n69318), .Y(n68958) );
  NOR2X1 U72184 ( .A(n69318), .B(n43598), .Y(n68956) );
  NAND2X1 U72185 ( .A(n68956), .B(n68955), .Y(n68957) );
  NAND2X1 U72186 ( .A(n68958), .B(n68957), .Y(n69147) );
  NAND2X1 U72187 ( .A(n68960), .B(n42999), .Y(n68963) );
  NOR2X1 U72188 ( .A(n68960), .B(n42998), .Y(n68962) );
  OR2X1 U72189 ( .A(n68962), .B(n68961), .Y(n69655) );
  INVX1 U72190 ( .A(n68964), .Y(n68973) );
  XNOR2X1 U72191 ( .A(n68973), .B(n68965), .Y(n68966) );
  NOR2X1 U72192 ( .A(n41418), .B(n41383), .Y(n68967) );
  NAND2X1 U72193 ( .A(n68966), .B(n39521), .Y(n69477) );
  NOR2X1 U72194 ( .A(n68973), .B(n68968), .Y(n68975) );
  NOR2X1 U72195 ( .A(n68970), .B(n68978), .Y(n68971) );
  NOR2X1 U72196 ( .A(n68973), .B(n68972), .Y(n68974) );
  NOR2X1 U72197 ( .A(n68975), .B(n68974), .Y(n68985) );
  NAND2X1 U72198 ( .A(n68979), .B(n68978), .Y(n68976) );
  NOR2X1 U72199 ( .A(n38986), .B(n68976), .Y(n68983) );
  NOR2X1 U72200 ( .A(n68978), .B(n68977), .Y(n68981) );
  NAND2X1 U72201 ( .A(n68979), .B(n44025), .Y(n68980) );
  NOR2X1 U72202 ( .A(n68981), .B(n68980), .Y(n68982) );
  NOR2X1 U72203 ( .A(n68983), .B(n68982), .Y(n68984) );
  NAND2X1 U72204 ( .A(n68985), .B(n68984), .Y(n69470) );
  INVX1 U72205 ( .A(n43001), .Y(n72515) );
  XNOR2X1 U72206 ( .A(n42187), .B(n72515), .Y(n71832) );
  INVX1 U72207 ( .A(n69450), .Y(n68987) );
  NAND2X1 U72208 ( .A(n68987), .B(n68986), .Y(n69447) );
  INVX1 U72209 ( .A(n69449), .Y(n68988) );
  NOR2X1 U72210 ( .A(n68988), .B(n68987), .Y(n68989) );
  NAND2X1 U72211 ( .A(n68989), .B(n69448), .Y(n68990) );
  NAND2X1 U72212 ( .A(n68991), .B(n68990), .Y(n68992) );
  NAND2X1 U72213 ( .A(n69447), .B(n68992), .Y(n69445) );
  INVX1 U72214 ( .A(n69445), .Y(n69468) );
  XNOR2X1 U72215 ( .A(n37370), .B(n69421), .Y(n68993) );
  XNOR2X1 U72216 ( .A(n68993), .B(n69003), .Y(n68994) );
  XNOR2X1 U72217 ( .A(n68995), .B(n68994), .Y(n69001) );
  NAND2X1 U72218 ( .A(n69001), .B(n68996), .Y(n69436) );
  NAND2X1 U72219 ( .A(n68997), .B(n44007), .Y(n68998) );
  NAND2X1 U72220 ( .A(n68999), .B(n68998), .Y(n69000) );
  OR2X1 U72221 ( .A(n69001), .B(n69000), .Y(n69002) );
  NAND2X1 U72222 ( .A(n41724), .B(n69002), .Y(n69439) );
  NAND2X1 U72223 ( .A(n69436), .B(n69439), .Y(n69444) );
  NAND2X1 U72224 ( .A(n43774), .B(n44048), .Y(n69462) );
  INVX1 U72225 ( .A(n69462), .Y(n69458) );
  XNOR2X1 U72226 ( .A(n41727), .B(n69458), .Y(n69141) );
  XNOR2X1 U72227 ( .A(n69003), .B(n37370), .Y(n69425) );
  INVX1 U72228 ( .A(n69425), .Y(n69420) );
  NAND2X1 U72229 ( .A(n69420), .B(n69004), .Y(n69010) );
  INVX1 U72230 ( .A(n69005), .Y(n69419) );
  INVX1 U72231 ( .A(n69006), .Y(n69418) );
  NOR2X1 U72232 ( .A(n69419), .B(n69418), .Y(n69007) );
  NAND2X1 U72233 ( .A(n69007), .B(n69425), .Y(n69008) );
  NAND2X1 U72234 ( .A(n69421), .B(n69008), .Y(n69009) );
  NAND2X1 U72235 ( .A(n69010), .B(n69009), .Y(n69432) );
  XNOR2X1 U72236 ( .A(n69054), .B(n69071), .Y(n69011) );
  INVX1 U72237 ( .A(n69050), .Y(n69038) );
  INVX1 U72238 ( .A(n69012), .Y(n69014) );
  NAND2X1 U72239 ( .A(n69015), .B(n69016), .Y(n69013) );
  NOR2X1 U72240 ( .A(n69014), .B(n69013), .Y(n69022) );
  INVX1 U72241 ( .A(n69015), .Y(n69049) );
  INVX1 U72242 ( .A(n69016), .Y(n69391) );
  NAND2X1 U72243 ( .A(n69049), .B(n69391), .Y(n69020) );
  NOR2X1 U72244 ( .A(n69041), .B(n69016), .Y(n69018) );
  NAND2X1 U72245 ( .A(n69018), .B(n69017), .Y(n69019) );
  NAND2X1 U72246 ( .A(n69020), .B(n69019), .Y(n69021) );
  NOR2X1 U72247 ( .A(n69022), .B(n69021), .Y(n69023) );
  XNOR2X1 U72248 ( .A(n69038), .B(n69023), .Y(n69404) );
  NAND2X1 U72249 ( .A(n69024), .B(n69404), .Y(n69025) );
  OR2X1 U72250 ( .A(n69026), .B(n69025), .Y(n69032) );
  INVX1 U72251 ( .A(n69032), .Y(n69028) );
  NAND2X1 U72252 ( .A(n38312), .B(n44017), .Y(n69029) );
  INVX1 U72253 ( .A(n69029), .Y(n69431) );
  INVX1 U72254 ( .A(n69400), .Y(n69406) );
  NAND2X1 U72255 ( .A(n69431), .B(n69406), .Y(n69027) );
  NOR2X1 U72256 ( .A(n69028), .B(n69027), .Y(n69031) );
  NOR2X1 U72257 ( .A(n69029), .B(n69407), .Y(n69030) );
  NOR2X1 U72258 ( .A(n69031), .B(n69030), .Y(n69036) );
  NOR2X1 U72259 ( .A(n69431), .B(n39500), .Y(n69034) );
  NAND2X1 U72260 ( .A(n69406), .B(n69032), .Y(n69033) );
  NAND2X1 U72261 ( .A(n69034), .B(n69033), .Y(n69035) );
  NAND2X1 U72262 ( .A(n69036), .B(n69035), .Y(n69139) );
  NAND2X1 U72263 ( .A(n69038), .B(n69037), .Y(n69388) );
  NOR2X1 U72264 ( .A(n69041), .B(n69039), .Y(n69043) );
  NOR2X1 U72265 ( .A(n69041), .B(n69040), .Y(n69042) );
  NOR2X1 U72266 ( .A(n69043), .B(n69042), .Y(n69047) );
  NAND2X1 U72267 ( .A(n69045), .B(n69044), .Y(n69046) );
  NAND2X1 U72268 ( .A(n69047), .B(n69046), .Y(n69048) );
  NOR2X1 U72269 ( .A(n69049), .B(n69048), .Y(n69051) );
  NAND2X1 U72270 ( .A(n69051), .B(n69050), .Y(n69390) );
  NAND2X1 U72271 ( .A(n69391), .B(n69390), .Y(n69052) );
  NAND2X1 U72272 ( .A(n69054), .B(n69053), .Y(n69376) );
  NOR2X1 U72273 ( .A(n69057), .B(n69055), .Y(n69059) );
  NOR2X1 U72274 ( .A(n69057), .B(n69056), .Y(n69058) );
  OR2X1 U72275 ( .A(n69059), .B(n69058), .Y(n69066) );
  INVX1 U72276 ( .A(n69124), .Y(n69064) );
  XNOR2X1 U72277 ( .A(n69060), .B(n69076), .Y(n69061) );
  XOR2X1 U72278 ( .A(n69062), .B(n69061), .Y(n69063) );
  XOR2X1 U72279 ( .A(n69064), .B(n69063), .Y(n69065) );
  NOR2X1 U72280 ( .A(n69066), .B(n69065), .Y(n69070) );
  NOR2X1 U72281 ( .A(n41005), .B(n69067), .Y(n69068) );
  NOR2X1 U72282 ( .A(n41250), .B(n69068), .Y(n69069) );
  NAND2X1 U72283 ( .A(n69070), .B(n69069), .Y(n69378) );
  NAND2X1 U72284 ( .A(n69071), .B(n69378), .Y(n69072) );
  NAND2X1 U72285 ( .A(n69376), .B(n69072), .Y(n69698) );
  NAND2X1 U72286 ( .A(n43991), .B(n43496), .Y(n69375) );
  INVX1 U72287 ( .A(n69375), .Y(n69699) );
  NAND2X1 U72288 ( .A(n43491), .B(n44000), .Y(n69389) );
  INVX1 U72289 ( .A(n69389), .Y(n69392) );
  XNOR2X1 U72290 ( .A(n69699), .B(n69392), .Y(n69136) );
  NAND2X1 U72291 ( .A(n69073), .B(n43934), .Y(n69075) );
  NAND2X1 U72292 ( .A(n69075), .B(n69074), .Y(n69077) );
  NAND2X1 U72293 ( .A(n69077), .B(n69076), .Y(n69104) );
  XNOR2X1 U72294 ( .A(n69079), .B(n69078), .Y(n69081) );
  NAND2X1 U72295 ( .A(n69081), .B(n69117), .Y(n69088) );
  INVX1 U72296 ( .A(n69088), .Y(n69083) );
  NOR2X1 U72297 ( .A(n69083), .B(n69082), .Y(n69086) );
  INVX1 U72298 ( .A(n69084), .Y(n69085) );
  NOR2X1 U72299 ( .A(n69086), .B(n69085), .Y(n69090) );
  OR2X1 U72300 ( .A(n69088), .B(n69087), .Y(n69089) );
  NAND2X1 U72301 ( .A(n69090), .B(n69089), .Y(n69091) );
  NOR2X1 U72302 ( .A(n69092), .B(n69091), .Y(n69100) );
  NOR2X1 U72303 ( .A(n69093), .B(n69096), .Y(n69098) );
  INVX1 U72304 ( .A(n69094), .Y(n69095) );
  NOR2X1 U72305 ( .A(n69096), .B(n69095), .Y(n69097) );
  NOR2X1 U72306 ( .A(n69098), .B(n69097), .Y(n69099) );
  NAND2X1 U72307 ( .A(n69100), .B(n69099), .Y(n69101) );
  NAND2X1 U72308 ( .A(n69102), .B(n69101), .Y(n69103) );
  NAND2X1 U72309 ( .A(n69104), .B(n69103), .Y(n69743) );
  INVX1 U72310 ( .A(n69743), .Y(n69331) );
  INVX1 U72311 ( .A(n69105), .Y(n71856) );
  NAND2X1 U72312 ( .A(n71856), .B(n72397), .Y(n69338) );
  NAND2X1 U72313 ( .A(n69338), .B(n71857), .Y(n71861) );
  INVX1 U72314 ( .A(n71861), .Y(n71523) );
  XNOR2X1 U72315 ( .A(n41862), .B(n71523), .Y(n69757) );
  INVX1 U72316 ( .A(n69757), .Y(n69358) );
  NAND2X1 U72317 ( .A(n69106), .B(n43604), .Y(n72280) );
  INVX1 U72318 ( .A(n72280), .Y(n72283) );
  XNOR2X1 U72319 ( .A(n41517), .B(n72283), .Y(n69111) );
  NAND2X1 U72320 ( .A(n69108), .B(n69107), .Y(n69110) );
  NAND2X1 U72321 ( .A(n69110), .B(n69109), .Y(n69352) );
  INVX1 U72322 ( .A(n69352), .Y(n69356) );
  XNOR2X1 U72323 ( .A(n69111), .B(n69356), .Y(n69112) );
  XNOR2X1 U72324 ( .A(n41690), .B(n69112), .Y(n69116) );
  INVX1 U72325 ( .A(n69117), .Y(n69113) );
  NAND2X1 U72326 ( .A(n72291), .B(n69113), .Y(n69115) );
  NAND2X1 U72327 ( .A(n72291), .B(n69118), .Y(n69114) );
  NAND2X1 U72328 ( .A(n69115), .B(n69114), .Y(n69335) );
  INVX1 U72329 ( .A(n69335), .Y(n69359) );
  XNOR2X1 U72330 ( .A(n69116), .B(n69359), .Y(n69122) );
  NAND2X1 U72331 ( .A(n69117), .B(n72288), .Y(n69119) );
  NOR2X1 U72332 ( .A(n69119), .B(n69118), .Y(n69121) );
  NOR2X1 U72333 ( .A(n69121), .B(n69120), .Y(n69362) );
  XNOR2X1 U72334 ( .A(n69122), .B(n69362), .Y(n69330) );
  XNOR2X1 U72335 ( .A(n69330), .B(n41526), .Y(n69123) );
  XNOR2X1 U72336 ( .A(n69331), .B(n69123), .Y(n69715) );
  NAND2X1 U72337 ( .A(n43982), .B(n43500), .Y(n69367) );
  NAND2X1 U72338 ( .A(n41683), .B(n69124), .Y(n69135) );
  NOR2X1 U72339 ( .A(n69128), .B(n69127), .Y(n69129) );
  NOR2X1 U72340 ( .A(n41683), .B(n69129), .Y(n69130) );
  NAND2X1 U72341 ( .A(n69131), .B(n69130), .Y(n69132) );
  NAND2X1 U72342 ( .A(n69133), .B(n69132), .Y(n69134) );
  NAND2X1 U72343 ( .A(n69135), .B(n69134), .Y(n69716) );
  XNOR2X1 U72344 ( .A(n69136), .B(n69385), .Y(n69137) );
  XNOR2X1 U72345 ( .A(n69698), .B(n69137), .Y(n69138) );
  NAND2X1 U72346 ( .A(n38310), .B(n44007), .Y(n69408) );
  INVX1 U72347 ( .A(n69408), .Y(n69688) );
  XNOR2X1 U72348 ( .A(n69139), .B(n41485), .Y(n69140) );
  INVX1 U72349 ( .A(n69438), .Y(n69464) );
  XNOR2X1 U72350 ( .A(n69141), .B(n41448), .Y(n69142) );
  XNOR2X1 U72351 ( .A(n71832), .B(n41442), .Y(n69143) );
  XNOR2X1 U72352 ( .A(n69470), .B(n69143), .Y(n69144) );
  XNOR2X1 U72353 ( .A(n41117), .B(n69144), .Y(n69316) );
  XNOR2X1 U72354 ( .A(n69316), .B(n43616), .Y(n69145) );
  XNOR2X1 U72355 ( .A(n40491), .B(n69145), .Y(n69146) );
  XNOR2X1 U72356 ( .A(n69147), .B(n69146), .Y(n69155) );
  NAND2X1 U72357 ( .A(n43615), .B(n69304), .Y(n69488) );
  NAND2X1 U72358 ( .A(n69149), .B(n40683), .Y(n69154) );
  NAND2X1 U72359 ( .A(n43615), .B(n69150), .Y(n69152) );
  NAND2X1 U72360 ( .A(n69152), .B(n69151), .Y(n69153) );
  NAND2X1 U72361 ( .A(n69154), .B(n69153), .Y(n69487) );
  XNOR2X1 U72362 ( .A(n69155), .B(n41637), .Y(n69311) );
  XNOR2X1 U72363 ( .A(n69627), .B(n43568), .Y(n69156) );
  NAND2X1 U72364 ( .A(n69498), .B(n40670), .Y(n69161) );
  NAND2X1 U72365 ( .A(n43567), .B(n69499), .Y(n69159) );
  NAND2X1 U72366 ( .A(n38179), .B(n69159), .Y(n69160) );
  NAND2X1 U72367 ( .A(n69161), .B(n69160), .Y(n69300) );
  INVX1 U72368 ( .A(n69293), .Y(n69294) );
  XNOR2X1 U72369 ( .A(n69162), .B(n69294), .Y(n69172) );
  INVX1 U72370 ( .A(n69163), .Y(n69166) );
  INVX1 U72371 ( .A(n69295), .Y(n69297) );
  NOR2X1 U72372 ( .A(n43582), .B(n69295), .Y(n69169) );
  NOR2X1 U72373 ( .A(n38151), .B(n69166), .Y(n69168) );
  NAND2X1 U72374 ( .A(n69168), .B(n69167), .Y(n69296) );
  NAND2X1 U72375 ( .A(n69169), .B(n69296), .Y(n69170) );
  XNOR2X1 U72376 ( .A(n69172), .B(n41134), .Y(n69189) );
  INVX1 U72377 ( .A(n69173), .Y(n69175) );
  NOR2X1 U72378 ( .A(n69175), .B(n69174), .Y(n69177) );
  NOR2X1 U72379 ( .A(n69177), .B(n69176), .Y(n69180) );
  NAND2X1 U72380 ( .A(n69178), .B(n39958), .Y(n69179) );
  NAND2X1 U72381 ( .A(n69180), .B(n69179), .Y(n69183) );
  NAND2X1 U72382 ( .A(n43577), .B(n69181), .Y(n69182) );
  NAND2X1 U72383 ( .A(n69183), .B(n69182), .Y(n69185) );
  INVX1 U72384 ( .A(n69185), .Y(n69287) );
  NOR2X1 U72385 ( .A(n69287), .B(n69289), .Y(n69187) );
  NAND2X1 U72386 ( .A(n69850), .B(n43579), .Y(n69184) );
  NOR2X1 U72387 ( .A(n69185), .B(n69184), .Y(n69186) );
  NOR2X1 U72388 ( .A(n69187), .B(n69186), .Y(n69188) );
  XNOR2X1 U72389 ( .A(n69189), .B(n69188), .Y(n69190) );
  XNOR2X1 U72390 ( .A(n40518), .B(n69190), .Y(n69198) );
  NAND2X1 U72391 ( .A(n40235), .B(n39187), .Y(n69196) );
  NAND2X1 U72392 ( .A(n39187), .B(n43559), .Y(n69195) );
  NAND2X1 U72393 ( .A(n69196), .B(n69195), .Y(n69192) );
  INVX1 U72394 ( .A(n69259), .Y(n69193) );
  NOR2X1 U72395 ( .A(n40954), .B(n69193), .Y(n69194) );
  NOR2X1 U72396 ( .A(n69194), .B(n43551), .Y(n69204) );
  NAND2X1 U72397 ( .A(n69197), .B(n69196), .Y(n69282) );
  OR2X1 U72398 ( .A(n43549), .B(n69258), .Y(n69202) );
  NAND2X1 U72399 ( .A(n69259), .B(n43549), .Y(n69199) );
  NOR2X1 U72400 ( .A(n40954), .B(n69199), .Y(n69200) );
  NAND2X1 U72401 ( .A(n69258), .B(n69200), .Y(n69201) );
  NAND2X1 U72402 ( .A(n69202), .B(n69201), .Y(n69203) );
  NOR2X1 U72403 ( .A(n69204), .B(n69203), .Y(n69205) );
  XNOR2X1 U72404 ( .A(n69206), .B(n69514), .Y(n69211) );
  INVX1 U72405 ( .A(n69517), .Y(n69523) );
  NAND2X1 U72406 ( .A(n43631), .B(n69516), .Y(n69208) );
  NOR2X1 U72407 ( .A(n43632), .B(n69517), .Y(n69210) );
  XNOR2X1 U72408 ( .A(n69211), .B(n41023), .Y(n69212) );
  XNOR2X1 U72409 ( .A(n69213), .B(n69212), .Y(n69872) );
  XNOR2X1 U72410 ( .A(n43661), .B(n69872), .Y(n69214) );
  INVX1 U72411 ( .A(n69551), .Y(n69550) );
  XNOR2X1 U72412 ( .A(n69217), .B(n41152), .Y(n69224) );
  XNOR2X1 U72413 ( .A(n41124), .B(n69218), .Y(n69580) );
  NOR2X1 U72414 ( .A(n69580), .B(n43514), .Y(n69219) );
  NAND2X1 U72415 ( .A(n43505), .B(n69220), .Y(n69221) );
  NOR2X1 U72416 ( .A(n36433), .B(n69222), .Y(n69223) );
  XNOR2X1 U72417 ( .A(n69224), .B(n69223), .Y(n69562) );
  XNOR2X1 U72418 ( .A(n69562), .B(n43692), .Y(n69232) );
  NOR2X1 U72419 ( .A(n69226), .B(n69225), .Y(n69227) );
  NOR2X1 U72420 ( .A(n43692), .B(n69227), .Y(n69228) );
  NOR2X1 U72421 ( .A(n41415), .B(n69228), .Y(n69230) );
  NAND2X1 U72422 ( .A(n69230), .B(n69229), .Y(n69560) );
  XNOR2X1 U72423 ( .A(n69241), .B(n43707), .Y(n69233) );
  XNOR2X1 U72424 ( .A(n69571), .B(n69233), .Y(n69238) );
  XNOR2X1 U72425 ( .A(n69235), .B(n69234), .Y(n69236) );
  XNOR2X1 U72426 ( .A(n69236), .B(n42070), .Y(n69237) );
  MX2X1 U72427 ( .A(n69238), .B(n69237), .S0(n43719), .Y(u_muldiv_result_r[21]) );
  NAND2X1 U72428 ( .A(u_muldiv_mult_result_q[21]), .B(n44632), .Y(n13940) );
  NAND2X1 U72429 ( .A(n69243), .B(n69242), .Y(n69537) );
  NAND2X1 U72430 ( .A(n43523), .B(n69244), .Y(n69890) );
  NAND2X1 U72431 ( .A(n69246), .B(n69245), .Y(n69889) );
  NAND2X1 U72432 ( .A(n69251), .B(n69247), .Y(n69248) );
  NAND2X1 U72433 ( .A(n69248), .B(n68550), .Y(n69249) );
  INVX1 U72434 ( .A(n69250), .Y(n69254) );
  NAND2X1 U72435 ( .A(n69252), .B(n69251), .Y(n69253) );
  NOR2X1 U72436 ( .A(n69254), .B(n69253), .Y(n69256) );
  NAND2X1 U72437 ( .A(n69256), .B(n69255), .Y(n69257) );
  INVX1 U72438 ( .A(n69872), .Y(n69875) );
  NAND2X1 U72439 ( .A(n40418), .B(n69258), .Y(n69263) );
  NAND2X1 U72440 ( .A(n69261), .B(n69260), .Y(n69262) );
  XNOR2X1 U72441 ( .A(n69263), .B(n69262), .Y(n69264) );
  NOR2X1 U72442 ( .A(n43545), .B(n69264), .Y(n69266) );
  NOR2X1 U72443 ( .A(n36678), .B(n39004), .Y(n69269) );
  NOR2X1 U72444 ( .A(n43620), .B(n69269), .Y(n69271) );
  NOR2X1 U72445 ( .A(n43620), .B(n69276), .Y(n69270) );
  NOR2X1 U72446 ( .A(n69271), .B(n69270), .Y(n69275) );
  XNOR2X1 U72447 ( .A(n69294), .B(n41134), .Y(n69849) );
  XNOR2X1 U72448 ( .A(n72149), .B(n39985), .Y(n69272) );
  XNOR2X1 U72449 ( .A(n69272), .B(n40518), .Y(n69273) );
  XNOR2X1 U72450 ( .A(n41013), .B(n69273), .Y(n69277) );
  NAND2X1 U72451 ( .A(n69277), .B(n43624), .Y(n69274) );
  NAND2X1 U72452 ( .A(n69275), .B(n69274), .Y(n69598) );
  NOR2X1 U72453 ( .A(n69276), .B(n38190), .Y(n69278) );
  XNOR2X1 U72454 ( .A(n69293), .B(n43537), .Y(n69279) );
  XNOR2X1 U72455 ( .A(n40518), .B(n69279), .Y(n69280) );
  NAND2X1 U72456 ( .A(n69280), .B(n43559), .Y(n69284) );
  INVX1 U72457 ( .A(n69280), .Y(n69281) );
  NAND2X1 U72458 ( .A(n43561), .B(n69281), .Y(n69283) );
  NAND2X1 U72459 ( .A(n39985), .B(n43539), .Y(n70124) );
  NAND2X1 U72460 ( .A(n43535), .B(n69849), .Y(n69285) );
  NAND2X1 U72461 ( .A(n69285), .B(n69620), .Y(n70123) );
  NAND2X1 U72462 ( .A(n70124), .B(n70123), .Y(n69608) );
  NAND2X1 U72463 ( .A(n43580), .B(n69288), .Y(n69286) );
  NAND2X1 U72464 ( .A(n69288), .B(n39958), .Y(n69289) );
  NOR2X1 U72465 ( .A(n41426), .B(n69289), .Y(n69290) );
  NAND2X1 U72466 ( .A(n69290), .B(n69849), .Y(n69292) );
  NAND2X1 U72467 ( .A(n43582), .B(n69297), .Y(n69298) );
  NAND2X1 U72468 ( .A(n69299), .B(n69840), .Y(n70115) );
  NAND2X1 U72469 ( .A(n38962), .B(n40670), .Y(n69303) );
  NAND2X1 U72470 ( .A(n43568), .B(n69627), .Y(n69301) );
  NAND2X1 U72471 ( .A(n69303), .B(n69302), .Y(n69842) );
  XNOR2X1 U72472 ( .A(n69842), .B(n43582), .Y(n69507) );
  NAND2X1 U72473 ( .A(n43617), .B(n69304), .Y(n69306) );
  NAND2X1 U72474 ( .A(n69306), .B(n69305), .Y(n69308) );
  NAND2X1 U72475 ( .A(n69308), .B(n69307), .Y(n69309) );
  NAND2X1 U72476 ( .A(n69310), .B(n69309), .Y(n69819) );
  NAND2X1 U72477 ( .A(n69311), .B(n42996), .Y(n69820) );
  NAND2X1 U72478 ( .A(n69820), .B(n69819), .Y(n69497) );
  NAND2X1 U72479 ( .A(n69313), .B(n69312), .Y(n69314) );
  NAND2X1 U72480 ( .A(n69314), .B(n43598), .Y(n69641) );
  NAND2X1 U72481 ( .A(n69315), .B(n43598), .Y(n69642) );
  NAND2X1 U72482 ( .A(n69641), .B(n69642), .Y(n69322) );
  NAND2X1 U72483 ( .A(n38222), .B(n43598), .Y(n69320) );
  NOR2X1 U72484 ( .A(n69318), .B(n69317), .Y(n69319) );
  NAND2X1 U72485 ( .A(n69319), .B(n38222), .Y(n69643) );
  NAND2X1 U72486 ( .A(n69320), .B(n69643), .Y(n69321) );
  NOR2X1 U72487 ( .A(n69322), .B(n69321), .Y(n69486) );
  NOR2X1 U72488 ( .A(n43597), .B(n69655), .Y(n69325) );
  XNOR2X1 U72489 ( .A(n41442), .B(n72515), .Y(n69323) );
  XNOR2X1 U72490 ( .A(n69323), .B(n38544), .Y(n69324) );
  XNOR2X1 U72491 ( .A(n41117), .B(n69324), .Y(n69656) );
  NAND2X1 U72492 ( .A(n39556), .B(n69656), .Y(n69645) );
  NAND2X1 U72493 ( .A(n69325), .B(n69645), .Y(n69329) );
  NOR2X1 U72494 ( .A(n43601), .B(n39555), .Y(n69327) );
  NAND2X1 U72495 ( .A(n69645), .B(n40491), .Y(n69326) );
  NAND2X1 U72496 ( .A(n69327), .B(n69326), .Y(n69328) );
  NAND2X1 U72497 ( .A(n69329), .B(n69328), .Y(n69484) );
  NAND2X1 U72498 ( .A(n43774), .B(n44055), .Y(n69804) );
  NAND2X1 U72499 ( .A(n38313), .B(n44025), .Y(n69796) );
  INVX1 U72500 ( .A(n69330), .Y(n69742) );
  NAND2X1 U72501 ( .A(n69742), .B(n69743), .Y(n69741) );
  NAND2X1 U72502 ( .A(n69331), .B(n69330), .Y(n69332) );
  NAND2X1 U72503 ( .A(n41526), .B(n69332), .Y(n69333) );
  NAND2X1 U72504 ( .A(n69741), .B(n69333), .Y(n69753) );
  NAND2X1 U72505 ( .A(n43982), .B(n39960), .Y(n69722) );
  NAND2X1 U72506 ( .A(n41690), .B(n69352), .Y(n69334) );
  NAND2X1 U72507 ( .A(n72283), .B(n69334), .Y(n69337) );
  NAND2X1 U72508 ( .A(n72283), .B(n69335), .Y(n69336) );
  NAND2X1 U72509 ( .A(n69337), .B(n69336), .Y(n69775) );
  INVX1 U72510 ( .A(n71862), .Y(n69341) );
  NAND2X1 U72511 ( .A(n69338), .B(n72296), .Y(n69342) );
  NAND2X1 U72512 ( .A(n69342), .B(n69339), .Y(n69756) );
  NAND2X1 U72513 ( .A(n69756), .B(n72288), .Y(n69340) );
  NOR2X1 U72514 ( .A(n69341), .B(n69340), .Y(n69350) );
  INVX1 U72515 ( .A(n69342), .Y(n69344) );
  NOR2X1 U72516 ( .A(n69344), .B(n69343), .Y(n69345) );
  NAND2X1 U72517 ( .A(n69345), .B(n72291), .Y(n69348) );
  NOR2X1 U72518 ( .A(n72296), .B(n72288), .Y(n69346) );
  NAND2X1 U72519 ( .A(n69346), .B(n71861), .Y(n69347) );
  NAND2X1 U72520 ( .A(n69348), .B(n69347), .Y(n69349) );
  NOR2X1 U72521 ( .A(n69350), .B(n69349), .Y(n69351) );
  XNOR2X1 U72522 ( .A(n69358), .B(n69351), .Y(n69989) );
  INVX1 U72523 ( .A(n69989), .Y(n69763) );
  XNOR2X1 U72524 ( .A(n72283), .B(n69763), .Y(n69767) );
  NAND2X1 U72525 ( .A(n69352), .B(n69358), .Y(n69353) );
  NAND2X1 U72526 ( .A(n72291), .B(n69353), .Y(n69762) );
  INVX1 U72527 ( .A(n69762), .Y(n69768) );
  NAND2X1 U72528 ( .A(n43972), .B(n43607), .Y(n69777) );
  NAND2X1 U72529 ( .A(n41517), .B(n43604), .Y(n72274) );
  XNOR2X1 U72530 ( .A(n69777), .B(n72274), .Y(n69354) );
  XOR2X1 U72531 ( .A(n69768), .B(n69354), .Y(n69355) );
  XNOR2X1 U72532 ( .A(n72291), .B(n72283), .Y(n72354) );
  XNOR2X1 U72533 ( .A(n72354), .B(n69356), .Y(n69357) );
  XNOR2X1 U72534 ( .A(n69358), .B(n69357), .Y(n69360) );
  XNOR2X1 U72535 ( .A(n69360), .B(n69359), .Y(n69361) );
  NAND2X1 U72536 ( .A(n41517), .B(n69361), .Y(n69724) );
  NAND2X1 U72537 ( .A(n69362), .B(n41517), .Y(n69725) );
  NAND2X1 U72538 ( .A(n69724), .B(n69725), .Y(n69727) );
  XNOR2X1 U72539 ( .A(n69722), .B(n69752), .Y(n69363) );
  XOR2X1 U72540 ( .A(n69753), .B(n69363), .Y(n69714) );
  INVX1 U72541 ( .A(n69367), .Y(n69717) );
  NAND2X1 U72542 ( .A(n69717), .B(n69368), .Y(n69711) );
  INVX1 U72543 ( .A(n69711), .Y(n69365) );
  NAND2X1 U72544 ( .A(n69716), .B(n69715), .Y(n69712) );
  NAND2X1 U72545 ( .A(n43991), .B(n43500), .Y(n69366) );
  NAND2X1 U72546 ( .A(n69712), .B(n69366), .Y(n69364) );
  NOR2X1 U72547 ( .A(n69365), .B(n69364), .Y(n69373) );
  INVX1 U72548 ( .A(n69712), .Y(n69721) );
  INVX1 U72549 ( .A(n69366), .Y(n69738) );
  NAND2X1 U72550 ( .A(n69721), .B(n69738), .Y(n69371) );
  NOR2X1 U72551 ( .A(n69367), .B(n69366), .Y(n69369) );
  NAND2X1 U72552 ( .A(n69369), .B(n69368), .Y(n69370) );
  NAND2X1 U72553 ( .A(n69371), .B(n69370), .Y(n69372) );
  NOR2X1 U72554 ( .A(n69373), .B(n69372), .Y(n69374) );
  XNOR2X1 U72555 ( .A(n69714), .B(n69374), .Y(n69706) );
  NAND2X1 U72556 ( .A(n43999), .B(n43497), .Y(n69697) );
  NOR2X1 U72557 ( .A(n69376), .B(n69375), .Y(n69377) );
  NOR2X1 U72558 ( .A(n41245), .B(n69377), .Y(n69384) );
  NAND2X1 U72559 ( .A(n69699), .B(n69378), .Y(n69379) );
  NOR2X1 U72560 ( .A(n69380), .B(n69379), .Y(n69382) );
  NAND2X1 U72561 ( .A(n69699), .B(n69385), .Y(n69700) );
  INVX1 U72562 ( .A(n69700), .Y(n69381) );
  NOR2X1 U72563 ( .A(n69382), .B(n69381), .Y(n69383) );
  NAND2X1 U72564 ( .A(n69384), .B(n69383), .Y(n69707) );
  XNOR2X1 U72565 ( .A(n69786), .B(n69790), .Y(n69399) );
  NOR2X1 U72566 ( .A(n41004), .B(n41246), .Y(n69387) );
  NOR2X1 U72567 ( .A(n41246), .B(n69389), .Y(n69386) );
  NOR2X1 U72568 ( .A(n69387), .B(n69386), .Y(n69398) );
  NOR2X1 U72569 ( .A(n69389), .B(n69388), .Y(n69396) );
  INVX1 U72570 ( .A(n69390), .Y(n69394) );
  NAND2X1 U72571 ( .A(n69392), .B(n69391), .Y(n69393) );
  NOR2X1 U72572 ( .A(n69394), .B(n69393), .Y(n69395) );
  NOR2X1 U72573 ( .A(n69396), .B(n69395), .Y(n69397) );
  NAND2X1 U72574 ( .A(n69398), .B(n69397), .Y(n69785) );
  INVX1 U72575 ( .A(n69785), .Y(n69788) );
  XNOR2X1 U72576 ( .A(n69399), .B(n69788), .Y(n69693) );
  INVX1 U72577 ( .A(n69693), .Y(n69691) );
  NAND2X1 U72578 ( .A(n38311), .B(n44016), .Y(n69409) );
  INVX1 U72579 ( .A(n69409), .Y(n69696) );
  NOR2X1 U72580 ( .A(n69404), .B(n69400), .Y(n69402) );
  NOR2X1 U72581 ( .A(n37370), .B(n69400), .Y(n69401) );
  NOR2X1 U72582 ( .A(n69696), .B(n69687), .Y(n69415) );
  NOR2X1 U72583 ( .A(n69409), .B(n69408), .Y(n69403) );
  NAND2X1 U72584 ( .A(n69403), .B(n69687), .Y(n69413) );
  NAND2X1 U72585 ( .A(n37370), .B(n69404), .Y(n69405) );
  NAND2X1 U72586 ( .A(n41239), .B(n69417), .Y(n69689) );
  NAND2X1 U72587 ( .A(n39520), .B(n69409), .Y(n69411) );
  NAND2X1 U72588 ( .A(n69411), .B(n69410), .Y(n69412) );
  NAND2X1 U72589 ( .A(n69413), .B(n69412), .Y(n69414) );
  NOR2X1 U72590 ( .A(n69415), .B(n69414), .Y(n69416) );
  XNOR2X1 U72591 ( .A(n69691), .B(n69416), .Y(n69797) );
  INVX1 U72592 ( .A(n69797), .Y(n69795) );
  INVX1 U72593 ( .A(n69433), .Y(n69429) );
  NOR2X1 U72594 ( .A(n69419), .B(n69418), .Y(n69423) );
  NAND2X1 U72595 ( .A(n69421), .B(n69420), .Y(n69422) );
  NAND2X1 U72596 ( .A(n69423), .B(n69422), .Y(n69427) );
  NAND2X1 U72597 ( .A(n69425), .B(n69424), .Y(n69426) );
  NAND2X1 U72598 ( .A(n69427), .B(n69426), .Y(n69428) );
  NAND2X1 U72599 ( .A(n69429), .B(n69428), .Y(n69430) );
  NAND2X1 U72600 ( .A(n69431), .B(n69430), .Y(n69435) );
  NAND2X1 U72601 ( .A(n69433), .B(n69432), .Y(n69434) );
  NAND2X1 U72602 ( .A(n69435), .B(n69434), .Y(n69794) );
  INVX1 U72603 ( .A(n69794), .Y(n69798) );
  NAND2X1 U72604 ( .A(n69438), .B(n69444), .Y(n69443) );
  INVX1 U72605 ( .A(n69436), .Y(n69437) );
  NOR2X1 U72606 ( .A(n69438), .B(n69437), .Y(n69440) );
  NAND2X1 U72607 ( .A(n69440), .B(n69439), .Y(n69441) );
  NAND2X1 U72608 ( .A(n41726), .B(n69441), .Y(n69442) );
  NAND2X1 U72609 ( .A(n69443), .B(n69442), .Y(n69684) );
  NAND2X1 U72610 ( .A(n43477), .B(n44048), .Y(n69681) );
  INVX1 U72611 ( .A(n69805), .Y(n69803) );
  XNOR2X1 U72612 ( .A(n69804), .B(n69803), .Y(n69461) );
  INVX1 U72613 ( .A(n69444), .Y(n69465) );
  XNOR2X1 U72614 ( .A(n41448), .B(n69465), .Y(n69455) );
  INVX1 U72615 ( .A(n69455), .Y(n69446) );
  NAND2X1 U72616 ( .A(n69446), .B(n69445), .Y(n69460) );
  INVX1 U72617 ( .A(n69448), .Y(n69452) );
  NAND2X1 U72618 ( .A(n69450), .B(n69449), .Y(n69451) );
  NOR2X1 U72619 ( .A(n69452), .B(n69451), .Y(n69454) );
  NAND2X1 U72620 ( .A(n69456), .B(n69455), .Y(n69457) );
  NAND2X1 U72621 ( .A(n69458), .B(n69457), .Y(n69459) );
  NAND2X1 U72622 ( .A(n69460), .B(n69459), .Y(n69802) );
  INVX1 U72623 ( .A(n69802), .Y(n69806) );
  XNOR2X1 U72624 ( .A(n69461), .B(n69806), .Y(n69974) );
  INVX1 U72625 ( .A(n69974), .Y(n69810) );
  NAND2X1 U72626 ( .A(n43613), .B(n43795), .Y(n72196) );
  INVX1 U72627 ( .A(n72196), .Y(n72510) );
  XNOR2X1 U72628 ( .A(n69462), .B(n41726), .Y(n69463) );
  XNOR2X1 U72629 ( .A(n69464), .B(n69463), .Y(n69466) );
  XNOR2X1 U72630 ( .A(n69466), .B(n69465), .Y(n69467) );
  XNOR2X1 U72631 ( .A(n69468), .B(n69467), .Y(n69471) );
  INVX1 U72632 ( .A(n69471), .Y(n69469) );
  NAND2X1 U72633 ( .A(n38544), .B(n69469), .Y(n69473) );
  NAND2X1 U72634 ( .A(n72510), .B(n69473), .Y(n69476) );
  NAND2X1 U72635 ( .A(n69471), .B(n69470), .Y(n69809) );
  INVX1 U72636 ( .A(n69809), .Y(n69472) );
  NOR2X1 U72637 ( .A(n72510), .B(n69472), .Y(n69474) );
  NAND2X1 U72638 ( .A(n41727), .B(n69473), .Y(n69808) );
  NAND2X1 U72639 ( .A(n69474), .B(n69808), .Y(n69475) );
  NAND2X1 U72640 ( .A(n69476), .B(n69475), .Y(n69965) );
  XNOR2X1 U72641 ( .A(n41442), .B(n38544), .Y(n69670) );
  NOR2X1 U72642 ( .A(n72515), .B(n69670), .Y(n69478) );
  NAND2X1 U72643 ( .A(n68967), .B(n69477), .Y(n69479) );
  NAND2X1 U72644 ( .A(n69478), .B(n69479), .Y(n69482) );
  INVX1 U72645 ( .A(n69670), .Y(n69668) );
  NOR2X1 U72646 ( .A(n69668), .B(n43001), .Y(n69480) );
  NAND2X1 U72647 ( .A(n69480), .B(n41117), .Y(n69481) );
  NAND2X1 U72648 ( .A(n69482), .B(n69481), .Y(n69653) );
  XNOR2X1 U72649 ( .A(n42999), .B(n69653), .Y(n69483) );
  XOR2X1 U72650 ( .A(n69675), .B(n69483), .Y(n69647) );
  XNOR2X1 U72651 ( .A(n69484), .B(n69647), .Y(n69485) );
  XNOR2X1 U72652 ( .A(n69486), .B(n69485), .Y(n70096) );
  XNOR2X1 U72653 ( .A(n43618), .B(n39306), .Y(n69493) );
  NAND2X1 U72654 ( .A(n69488), .B(n69487), .Y(n69634) );
  NAND2X1 U72655 ( .A(n69489), .B(n69639), .Y(n69492) );
  NOR2X1 U72656 ( .A(n69639), .B(n69634), .Y(n69490) );
  NAND2X1 U72657 ( .A(n69490), .B(n43616), .Y(n69491) );
  NOR2X1 U72658 ( .A(n69493), .B(n37372), .Y(n69495) );
  NOR2X1 U72659 ( .A(n69495), .B(n69494), .Y(n69496) );
  XOR2X1 U72660 ( .A(n69497), .B(n69496), .Y(n69830) );
  XNOR2X1 U72661 ( .A(n40670), .B(n69830), .Y(n69506) );
  NAND2X1 U72662 ( .A(n69498), .B(n42992), .Y(n69501) );
  NAND2X1 U72663 ( .A(n69627), .B(n42992), .Y(n69502) );
  NOR2X1 U72664 ( .A(n69502), .B(n39746), .Y(n69503) );
  NOR2X1 U72665 ( .A(n69504), .B(n69503), .Y(n69505) );
  XNOR2X1 U72666 ( .A(n69506), .B(n69505), .Y(n69843) );
  XNOR2X1 U72667 ( .A(n69507), .B(n69843), .Y(n69617) );
  XNOR2X1 U72668 ( .A(n69617), .B(n43537), .Y(n69508) );
  XNOR2X1 U72669 ( .A(n69846), .B(n69508), .Y(n69509) );
  XNOR2X1 U72670 ( .A(n41182), .B(n69509), .Y(n69607) );
  XNOR2X1 U72671 ( .A(n69607), .B(n71794), .Y(n69510) );
  XNOR2X1 U72672 ( .A(n69608), .B(n69510), .Y(n69511) );
  XNOR2X1 U72673 ( .A(n38826), .B(n69511), .Y(n69600) );
  XNOR2X1 U72674 ( .A(n71810), .B(n69600), .Y(n69512) );
  INVX1 U72675 ( .A(n69524), .Y(n69531) );
  INVX1 U72676 ( .A(n69522), .Y(n69518) );
  NOR2X1 U72677 ( .A(n69517), .B(n69518), .Y(n69519) );
  NOR2X1 U72678 ( .A(n43632), .B(n69519), .Y(n69520) );
  NOR2X1 U72679 ( .A(n69523), .B(n69522), .Y(n69525) );
  XNOR2X1 U72680 ( .A(n69601), .B(n43643), .Y(n69526) );
  XNOR2X1 U72681 ( .A(n69597), .B(n69526), .Y(n69588) );
  NAND2X1 U72682 ( .A(n69529), .B(n69528), .Y(n69530) );
  XNOR2X1 U72683 ( .A(n41023), .B(n69531), .Y(n69867) );
  NAND2X1 U72684 ( .A(n38283), .B(n43669), .Y(n69532) );
  NOR2X1 U72685 ( .A(n40959), .B(n69532), .Y(n69533) );
  XNOR2X1 U72686 ( .A(n69587), .B(n43655), .Y(n69534) );
  XOR2X1 U72687 ( .A(n40481), .B(n69535), .Y(n69885) );
  NAND2X1 U72688 ( .A(n43653), .B(n69538), .Y(n69592) );
  NAND2X1 U72689 ( .A(n69537), .B(n39495), .Y(n69886) );
  INVX1 U72690 ( .A(n69538), .Y(n69539) );
  NAND2X1 U72691 ( .A(n69539), .B(n43657), .Y(n69887) );
  NAND2X1 U72692 ( .A(n69887), .B(n69886), .Y(n69540) );
  XNOR2X1 U72693 ( .A(n41033), .B(n69574), .Y(n70479) );
  XNOR2X1 U72694 ( .A(n70479), .B(n43679), .Y(n69541) );
  XNOR2X1 U72695 ( .A(n43509), .B(n69541), .Y(n69552) );
  NOR2X1 U72696 ( .A(n69543), .B(n69542), .Y(n69544) );
  NAND2X1 U72697 ( .A(n69544), .B(n69548), .Y(n69545) );
  NOR2X1 U72698 ( .A(n69547), .B(n69546), .Y(n69549) );
  INVX1 U72699 ( .A(n70480), .Y(n69894) );
  XNOR2X1 U72700 ( .A(n69552), .B(n69894), .Y(n69559) );
  XNOR2X1 U72701 ( .A(n41138), .B(n41152), .Y(n69583) );
  NOR2X1 U72702 ( .A(n69583), .B(n69553), .Y(n69557) );
  NAND2X1 U72703 ( .A(n43505), .B(n69554), .Y(n69582) );
  NAND2X1 U72704 ( .A(n69555), .B(n69582), .Y(n69556) );
  NOR2X1 U72705 ( .A(n69557), .B(n69556), .Y(n69558) );
  XNOR2X1 U72706 ( .A(n69559), .B(n69558), .Y(n70184) );
  XNOR2X1 U72707 ( .A(n70184), .B(n43692), .Y(n69564) );
  NAND2X1 U72708 ( .A(n39157), .B(n36434), .Y(n69561) );
  OR2X1 U72709 ( .A(n69560), .B(n69561), .Y(n70185) );
  NAND2X1 U72710 ( .A(n43691), .B(n39157), .Y(n69563) );
  XNOR2X1 U72711 ( .A(n40456), .B(n69572), .Y(n69565) );
  XNOR2X1 U72712 ( .A(n69567), .B(n69566), .Y(n69568) );
  XOR2X1 U72713 ( .A(n42079), .B(n69568), .Y(n69569) );
  MX2X1 U72714 ( .A(n69570), .B(n69569), .S0(n43718), .Y(u_muldiv_result_r[22]) );
  NAND2X1 U72715 ( .A(u_muldiv_mult_result_q[22]), .B(n44632), .Y(n13932) );
  NOR2X1 U72716 ( .A(n39012), .B(n39906), .Y(n69577) );
  XNOR2X1 U72717 ( .A(n38047), .B(n41033), .Y(n69575) );
  XNOR2X1 U72718 ( .A(n69574), .B(n69575), .Y(n69576) );
  XNOR2X1 U72719 ( .A(n69577), .B(n69576), .Y(n69578) );
  NAND2X1 U72720 ( .A(n43505), .B(n69578), .Y(n70205) );
  NOR2X1 U72721 ( .A(n69580), .B(n69579), .Y(n69581) );
  NAND2X1 U72722 ( .A(n69584), .B(n43646), .Y(n69586) );
  NAND2X1 U72723 ( .A(n69586), .B(n69585), .Y(n69918) );
  XNOR2X1 U72724 ( .A(n69588), .B(n39655), .Y(n69589) );
  INVX1 U72725 ( .A(n69596), .Y(n69590) );
  NAND2X1 U72726 ( .A(n43653), .B(n69590), .Y(n69595) );
  NAND2X1 U72727 ( .A(n69592), .B(n69591), .Y(n69593) );
  NAND2X1 U72728 ( .A(n69593), .B(n69887), .Y(n69594) );
  INVX1 U72729 ( .A(n69916), .Y(n69917) );
  NOR2X1 U72730 ( .A(n69598), .B(n36775), .Y(n69599) );
  XOR2X1 U72731 ( .A(n69600), .B(n69599), .Y(n69604) );
  INVX1 U72732 ( .A(n69604), .Y(n69603) );
  NAND2X1 U72733 ( .A(n43631), .B(n69604), .Y(n69602) );
  NAND2X1 U72734 ( .A(n69603), .B(n43550), .Y(n70152) );
  NAND2X1 U72735 ( .A(n43544), .B(n69604), .Y(n69606) );
  NAND2X1 U72736 ( .A(n69606), .B(n69605), .Y(n70151) );
  INVX1 U72737 ( .A(n69607), .Y(n69614) );
  XNOR2X1 U72738 ( .A(n43566), .B(n69614), .Y(n69609) );
  INVX1 U72739 ( .A(n69608), .Y(n69613) );
  XNOR2X1 U72740 ( .A(n69609), .B(n69613), .Y(n69610) );
  XNOR2X1 U72741 ( .A(n38826), .B(n69610), .Y(n69611) );
  NAND2X1 U72742 ( .A(n43619), .B(n69611), .Y(n69941) );
  NAND2X1 U72743 ( .A(n69940), .B(n39030), .Y(n69612) );
  NAND2X1 U72744 ( .A(n70147), .B(n69612), .Y(n69860) );
  XNOR2X1 U72745 ( .A(n69614), .B(n69613), .Y(n69616) );
  INVX1 U72746 ( .A(n69616), .Y(n69615) );
  NAND2X1 U72747 ( .A(n69615), .B(n39629), .Y(n70138) );
  INVX1 U72748 ( .A(n69854), .Y(n70125) );
  NAND2X1 U72749 ( .A(n41182), .B(n70125), .Y(n70129) );
  INVX1 U72750 ( .A(n70124), .Y(n69618) );
  NOR2X1 U72751 ( .A(n38982), .B(n69619), .Y(n69624) );
  NAND2X1 U72752 ( .A(n43535), .B(n70129), .Y(n69622) );
  NAND2X1 U72753 ( .A(n39985), .B(n69620), .Y(n69621) );
  NOR2X1 U72754 ( .A(n69622), .B(n69621), .Y(n69623) );
  NOR2X1 U72755 ( .A(n43593), .B(n69625), .Y(n69630) );
  OR2X1 U72756 ( .A(n69627), .B(n69626), .Y(n69628) );
  NOR2X1 U72757 ( .A(n69830), .B(n69628), .Y(n69629) );
  NOR2X1 U72758 ( .A(n69630), .B(n69629), .Y(n69632) );
  INVX1 U72759 ( .A(n69830), .Y(n69832) );
  NAND2X1 U72760 ( .A(n69832), .B(n42992), .Y(n69631) );
  NAND2X1 U72761 ( .A(n69631), .B(n69632), .Y(n69945) );
  NAND2X1 U72762 ( .A(n69633), .B(n69634), .Y(n69635) );
  NOR2X1 U72763 ( .A(n38222), .B(n69635), .Y(n69636) );
  NOR2X1 U72764 ( .A(n43615), .B(n69636), .Y(n69638) );
  NOR2X1 U72765 ( .A(n43616), .B(n70096), .Y(n69637) );
  NOR2X1 U72766 ( .A(n41637), .B(n69639), .Y(n69640) );
  XNOR2X1 U72767 ( .A(n69947), .B(n43593), .Y(n69818) );
  NAND2X1 U72768 ( .A(n69644), .B(n69643), .Y(n70082) );
  INVX1 U72769 ( .A(n70082), .Y(n70085) );
  NAND2X1 U72770 ( .A(n69645), .B(n40491), .Y(n69659) );
  NAND2X1 U72771 ( .A(n69659), .B(n69646), .Y(n69952) );
  NAND2X1 U72772 ( .A(n43600), .B(n70087), .Y(n69648) );
  NOR2X1 U72773 ( .A(n70085), .B(n69648), .Y(n69652) );
  INVX1 U72774 ( .A(n70087), .Y(n69649) );
  NAND2X1 U72775 ( .A(n69649), .B(n43598), .Y(n69650) );
  NOR2X1 U72776 ( .A(n69650), .B(n70082), .Y(n69651) );
  INVX1 U72777 ( .A(n69675), .Y(n69677) );
  INVX1 U72778 ( .A(n69953), .Y(n69654) );
  NOR2X1 U72779 ( .A(n69654), .B(n40683), .Y(n69658) );
  OR2X1 U72780 ( .A(n69656), .B(n69655), .Y(n69657) );
  NOR2X1 U72781 ( .A(n42998), .B(n69657), .Y(n69663) );
  NAND2X1 U72782 ( .A(n69658), .B(n69663), .Y(n69667) );
  NOR2X1 U72783 ( .A(n39556), .B(n39555), .Y(n69660) );
  NAND2X1 U72784 ( .A(n69660), .B(n69659), .Y(n69661) );
  NOR2X1 U72785 ( .A(n69953), .B(n69661), .Y(n69662) );
  NOR2X1 U72786 ( .A(n43616), .B(n69662), .Y(n69665) );
  NAND2X1 U72787 ( .A(n69663), .B(n69953), .Y(n69664) );
  NAND2X1 U72788 ( .A(n69665), .B(n69664), .Y(n69666) );
  NAND2X1 U72789 ( .A(n69667), .B(n69666), .Y(n69816) );
  NAND2X1 U72790 ( .A(n72515), .B(n69668), .Y(n69669) );
  NAND2X1 U72791 ( .A(n41117), .B(n69669), .Y(n69672) );
  NAND2X1 U72792 ( .A(n69670), .B(n43000), .Y(n69671) );
  NAND2X1 U72793 ( .A(n69672), .B(n69671), .Y(n69673) );
  INVX1 U72794 ( .A(n69673), .Y(n69674) );
  NOR2X1 U72795 ( .A(n69675), .B(n69674), .Y(n69676) );
  NOR2X1 U72796 ( .A(n39274), .B(n69676), .Y(n69679) );
  NAND2X1 U72797 ( .A(n69677), .B(n43001), .Y(n69678) );
  NAND2X1 U72798 ( .A(n43613), .B(n43774), .Y(n72202) );
  INVX1 U72799 ( .A(n72202), .Y(n72200) );
  XNOR2X1 U72800 ( .A(n41731), .B(n72200), .Y(n69686) );
  INVX1 U72801 ( .A(n69685), .Y(n69680) );
  NOR2X1 U72802 ( .A(n69680), .B(n69681), .Y(n69683) );
  NOR2X1 U72803 ( .A(n39260), .B(n69681), .Y(n69682) );
  XNOR2X1 U72804 ( .A(n69686), .B(n39047), .Y(n69801) );
  NAND2X1 U72805 ( .A(n43487), .B(n44025), .Y(n70042) );
  NAND2X1 U72806 ( .A(n69688), .B(n69687), .Y(n69690) );
  NAND2X1 U72807 ( .A(n69690), .B(n69689), .Y(n69692) );
  INVX1 U72808 ( .A(n69692), .Y(n69694) );
  NAND2X1 U72809 ( .A(n69694), .B(n69693), .Y(n69695) );
  XNOR2X1 U72810 ( .A(n70042), .B(n38264), .Y(n69793) );
  INVX1 U72811 ( .A(n69697), .Y(n69705) );
  NAND2X1 U72812 ( .A(n69699), .B(n69698), .Y(n69701) );
  NAND2X1 U72813 ( .A(n69701), .B(n69700), .Y(n69702) );
  NOR2X1 U72814 ( .A(n41245), .B(n69702), .Y(n69703) );
  NAND2X1 U72815 ( .A(n69703), .B(n69706), .Y(n69704) );
  NAND2X1 U72816 ( .A(n69705), .B(n69704), .Y(n69710) );
  INVX1 U72817 ( .A(n69706), .Y(n69708) );
  NAND2X1 U72818 ( .A(n69708), .B(n69707), .Y(n69709) );
  NAND2X1 U72819 ( .A(n69710), .B(n69709), .Y(n70023) );
  NAND2X1 U72820 ( .A(n69712), .B(n69711), .Y(n69713) );
  NAND2X1 U72821 ( .A(n69714), .B(n69713), .Y(n69740) );
  NAND2X1 U72822 ( .A(n69717), .B(n69715), .Y(n69719) );
  NAND2X1 U72823 ( .A(n69717), .B(n69716), .Y(n69718) );
  NAND2X1 U72824 ( .A(n69719), .B(n69718), .Y(n69720) );
  NOR2X1 U72825 ( .A(n69721), .B(n69720), .Y(n69736) );
  INVX1 U72826 ( .A(n69753), .Y(n69734) );
  INVX1 U72827 ( .A(n69722), .Y(n69751) );
  XNOR2X1 U72828 ( .A(n69751), .B(n69723), .Y(n69726) );
  NOR2X1 U72829 ( .A(n69726), .B(n69724), .Y(n69732) );
  NOR2X1 U72830 ( .A(n69726), .B(n69725), .Y(n69730) );
  INVX1 U72831 ( .A(n69726), .Y(n69728) );
  NOR2X1 U72832 ( .A(n69728), .B(n69727), .Y(n69729) );
  OR2X1 U72833 ( .A(n69730), .B(n69729), .Y(n69731) );
  NOR2X1 U72834 ( .A(n69732), .B(n69731), .Y(n69733) );
  XOR2X1 U72835 ( .A(n69734), .B(n69733), .Y(n69735) );
  NAND2X1 U72836 ( .A(n69736), .B(n69735), .Y(n69737) );
  NAND2X1 U72837 ( .A(n69738), .B(n69737), .Y(n69739) );
  NAND2X1 U72838 ( .A(n69740), .B(n69739), .Y(n70323) );
  INVX1 U72839 ( .A(n70323), .Y(n70020) );
  NAND2X1 U72840 ( .A(n43991), .B(n39961), .Y(n70010) );
  INVX1 U72841 ( .A(n69741), .Y(n69747) );
  NAND2X1 U72842 ( .A(n69742), .B(n41526), .Y(n69745) );
  NAND2X1 U72843 ( .A(n41526), .B(n69743), .Y(n69744) );
  NAND2X1 U72844 ( .A(n69745), .B(n69744), .Y(n69746) );
  NOR2X1 U72845 ( .A(n69747), .B(n69746), .Y(n69749) );
  INVX1 U72846 ( .A(n69752), .Y(n69748) );
  NAND2X1 U72847 ( .A(n69749), .B(n69748), .Y(n69750) );
  NAND2X1 U72848 ( .A(n69751), .B(n69750), .Y(n69755) );
  NAND2X1 U72849 ( .A(n69753), .B(n69752), .Y(n69754) );
  NAND2X1 U72850 ( .A(n69755), .B(n69754), .Y(n70286) );
  INVX1 U72851 ( .A(n70286), .Y(n70012) );
  XNOR2X1 U72852 ( .A(n70010), .B(n70012), .Y(n69781) );
  INVX1 U72853 ( .A(n72274), .Y(n72326) );
  XNOR2X1 U72854 ( .A(n69989), .B(n72283), .Y(n69760) );
  NAND2X1 U72855 ( .A(n71862), .B(n69756), .Y(n71865) );
  NAND2X1 U72856 ( .A(n72291), .B(n71865), .Y(n69759) );
  NAND2X1 U72857 ( .A(n72291), .B(n69757), .Y(n69758) );
  NAND2X1 U72858 ( .A(n69759), .B(n69758), .Y(n71872) );
  INVX1 U72859 ( .A(n69992), .Y(n70299) );
  NAND2X1 U72860 ( .A(n43982), .B(n43607), .Y(n70006) );
  INVX1 U72861 ( .A(n70006), .Y(n69991) );
  INVX1 U72862 ( .A(n69777), .Y(n69761) );
  NAND2X1 U72863 ( .A(n69761), .B(n43604), .Y(n72268) );
  INVX1 U72864 ( .A(n72268), .Y(n72355) );
  XNOR2X1 U72865 ( .A(n69991), .B(n72355), .Y(n69765) );
  NAND2X1 U72866 ( .A(n69763), .B(n69762), .Y(n69764) );
  NAND2X1 U72867 ( .A(n72283), .B(n69764), .Y(n69993) );
  INVX1 U72868 ( .A(n69993), .Y(n69997) );
  XNOR2X1 U72869 ( .A(n69765), .B(n69997), .Y(n69766) );
  XNOR2X1 U72870 ( .A(n41692), .B(n69766), .Y(n69772) );
  NAND2X1 U72871 ( .A(n72326), .B(n69773), .Y(n69770) );
  NAND2X1 U72872 ( .A(n72326), .B(n69775), .Y(n69769) );
  NAND2X1 U72873 ( .A(n69770), .B(n69769), .Y(n70004) );
  INVX1 U72874 ( .A(n70004), .Y(n69771) );
  XNOR2X1 U72875 ( .A(n69772), .B(n69771), .Y(n69780) );
  INVX1 U72876 ( .A(n69773), .Y(n69774) );
  NAND2X1 U72877 ( .A(n69774), .B(n72274), .Y(n69776) );
  NOR2X1 U72878 ( .A(n69776), .B(n69775), .Y(n69778) );
  NOR2X1 U72879 ( .A(n69778), .B(n69777), .Y(n69779) );
  XNOR2X1 U72880 ( .A(n69780), .B(n69779), .Y(n70285) );
  INVX1 U72881 ( .A(n70285), .Y(n70011) );
  XNOR2X1 U72882 ( .A(n69781), .B(n70011), .Y(n70021) );
  NAND2X1 U72883 ( .A(n43999), .B(n43500), .Y(n70016) );
  XNOR2X1 U72884 ( .A(n70016), .B(n42033), .Y(n69782) );
  XNOR2X1 U72885 ( .A(n70021), .B(n69782), .Y(n69783) );
  XNOR2X1 U72886 ( .A(n70020), .B(n69783), .Y(n70030) );
  XNOR2X1 U72887 ( .A(n70030), .B(n41529), .Y(n69784) );
  NAND2X1 U72888 ( .A(n69786), .B(n69785), .Y(n69792) );
  INVX1 U72889 ( .A(n69786), .Y(n69787) );
  NAND2X1 U72890 ( .A(n69788), .B(n69787), .Y(n69789) );
  NAND2X1 U72891 ( .A(n69790), .B(n69789), .Y(n69791) );
  NAND2X1 U72892 ( .A(n69792), .B(n69791), .Y(n70033) );
  INVX1 U72893 ( .A(n70047), .Y(n70043) );
  XNOR2X1 U72894 ( .A(n69793), .B(n70043), .Y(n70055) );
  NAND2X1 U72895 ( .A(n43484), .B(n44048), .Y(n70054) );
  NAND2X1 U72896 ( .A(n69795), .B(n69794), .Y(n70058) );
  INVX1 U72897 ( .A(n69796), .Y(n69799) );
  NAND2X1 U72898 ( .A(n69798), .B(n69797), .Y(n70056) );
  NAND2X1 U72899 ( .A(n69799), .B(n70056), .Y(n69800) );
  NAND2X1 U72900 ( .A(n70058), .B(n69800), .Y(n70052) );
  INVX1 U72901 ( .A(n70065), .Y(n69985) );
  XNOR2X1 U72902 ( .A(n69801), .B(n69985), .Y(n69959) );
  XNOR2X1 U72903 ( .A(n72515), .B(n72510), .Y(n70077) );
  INVX1 U72904 ( .A(n70077), .Y(n71582) );
  XNOR2X1 U72905 ( .A(n69959), .B(n71582), .Y(n69807) );
  NAND2X1 U72906 ( .A(n69803), .B(n69802), .Y(n70069) );
  NAND2X1 U72907 ( .A(n70069), .B(n70068), .Y(n70393) );
  INVX1 U72908 ( .A(n70393), .Y(n69977) );
  XNOR2X1 U72909 ( .A(n69807), .B(n69977), .Y(n69814) );
  NAND2X1 U72910 ( .A(n69809), .B(n69808), .Y(n69973) );
  NOR2X1 U72911 ( .A(n69974), .B(n69973), .Y(n69813) );
  NAND2X1 U72912 ( .A(n69810), .B(n72196), .Y(n69975) );
  OR2X1 U72913 ( .A(n72510), .B(n69973), .Y(n69811) );
  NAND2X1 U72914 ( .A(n69975), .B(n69811), .Y(n69812) );
  NOR2X1 U72915 ( .A(n69813), .B(n69812), .Y(n69962) );
  XNOR2X1 U72916 ( .A(n69814), .B(n69962), .Y(n69815) );
  XNOR2X1 U72917 ( .A(n41647), .B(n69815), .Y(n70084) );
  INVX1 U72918 ( .A(n70084), .Y(n70086) );
  XNOR2X1 U72919 ( .A(n69816), .B(n70086), .Y(n69817) );
  XNOR2X1 U72920 ( .A(n69818), .B(n41638), .Y(n69825) );
  NOR2X1 U72921 ( .A(n70096), .B(n42995), .Y(n69821) );
  NAND2X1 U72922 ( .A(n69820), .B(n69819), .Y(n70097) );
  NAND2X1 U72923 ( .A(n69821), .B(n70097), .Y(n69823) );
  NOR2X1 U72924 ( .A(n38899), .B(n69823), .Y(n69829) );
  NOR2X1 U72925 ( .A(n69822), .B(n38899), .Y(n69827) );
  NAND2X1 U72926 ( .A(n69823), .B(n69822), .Y(n69824) );
  NOR2X1 U72927 ( .A(n69825), .B(n69824), .Y(n69826) );
  OR2X1 U72928 ( .A(n69827), .B(n69826), .Y(n69828) );
  NOR2X1 U72929 ( .A(n69829), .B(n69828), .Y(n69943) );
  XNOR2X1 U72930 ( .A(n38191), .B(n69943), .Y(n70109) );
  XNOR2X1 U72931 ( .A(n70109), .B(n43568), .Y(n69838) );
  INVX1 U72932 ( .A(n70726), .Y(n72152) );
  NAND2X1 U72933 ( .A(n43568), .B(n69830), .Y(n69831) );
  NAND2X1 U72934 ( .A(n69831), .B(n69842), .Y(n70111) );
  NOR2X1 U72935 ( .A(n72152), .B(n70111), .Y(n69836) );
  NAND2X1 U72936 ( .A(n70111), .B(n72152), .Y(n69834) );
  NAND2X1 U72937 ( .A(n69832), .B(n40670), .Y(n70110) );
  NAND2X1 U72938 ( .A(n69834), .B(n69833), .Y(n69835) );
  NOR2X1 U72939 ( .A(n69836), .B(n69835), .Y(n69837) );
  XNOR2X1 U72940 ( .A(n69838), .B(n69837), .Y(n69848) );
  NOR2X1 U72941 ( .A(n39284), .B(n69840), .Y(n69841) );
  NOR2X1 U72942 ( .A(n43582), .B(n69841), .Y(n69845) );
  NOR2X1 U72943 ( .A(n43582), .B(n39983), .Y(n69844) );
  XNOR2X1 U72944 ( .A(n39372), .B(n69848), .Y(n69858) );
  NOR2X1 U72945 ( .A(n43578), .B(n69849), .Y(n69853) );
  NOR2X1 U72946 ( .A(n69850), .B(n41426), .Y(n69851) );
  NOR2X1 U72947 ( .A(n43579), .B(n69851), .Y(n69852) );
  NOR2X1 U72948 ( .A(n69853), .B(n69852), .Y(n69857) );
  NAND2X1 U72949 ( .A(n69855), .B(n69854), .Y(n69856) );
  NAND2X1 U72950 ( .A(n69857), .B(n69856), .Y(n70118) );
  XNOR2X1 U72951 ( .A(n43553), .B(n70144), .Y(n69859) );
  XNOR2X1 U72952 ( .A(n69922), .B(n69861), .Y(n69862) );
  NAND2X1 U72953 ( .A(n43665), .B(n70453), .Y(n69870) );
  NOR2X1 U72954 ( .A(n43665), .B(n38283), .Y(n69864) );
  NOR2X1 U72955 ( .A(n40167), .B(n69864), .Y(n69866) );
  INVX1 U72956 ( .A(n38388), .Y(n69868) );
  NAND2X1 U72957 ( .A(n69868), .B(n43669), .Y(n69927) );
  NAND2X1 U72958 ( .A(n69928), .B(n69927), .Y(n69869) );
  NAND2X1 U72959 ( .A(n69870), .B(n69869), .Y(n69871) );
  NAND2X1 U72960 ( .A(n41358), .B(n69872), .Y(n69873) );
  OR2X1 U72961 ( .A(n38154), .B(n69873), .Y(n69874) );
  NOR2X1 U72962 ( .A(n69878), .B(n69874), .Y(n70158) );
  NOR2X1 U72963 ( .A(n69875), .B(n69916), .Y(n69876) );
  NAND2X1 U72964 ( .A(n69876), .B(n41358), .Y(n70159) );
  INVX1 U72965 ( .A(n70159), .Y(n69879) );
  XNOR2X1 U72966 ( .A(n69877), .B(n41017), .Y(n69878) );
  NOR2X1 U72967 ( .A(n69879), .B(n39511), .Y(n69883) );
  NOR2X1 U72968 ( .A(n69917), .B(n39301), .Y(n69881) );
  NAND2X1 U72969 ( .A(n69881), .B(n69880), .Y(n69882) );
  INVX1 U72970 ( .A(n38174), .Y(n69888) );
  NAND2X1 U72971 ( .A(n43522), .B(n69888), .Y(n70165) );
  NAND2X1 U72972 ( .A(n70167), .B(n43528), .Y(n69892) );
  NAND2X1 U72973 ( .A(n69890), .B(n69889), .Y(n69891) );
  NAND2X1 U72974 ( .A(n69892), .B(n69891), .Y(n70164) );
  NOR2X1 U72975 ( .A(n36544), .B(n43687), .Y(n69893) );
  NOR2X1 U72976 ( .A(n69894), .B(n69893), .Y(n69895) );
  NOR2X1 U72977 ( .A(n38046), .B(n69895), .Y(n69896) );
  XOR2X1 U72978 ( .A(n70178), .B(n69896), .Y(n70181) );
  XNOR2X1 U72979 ( .A(n70181), .B(n43508), .Y(n69897) );
  XNOR2X1 U72980 ( .A(n70190), .B(n43692), .Y(n69905) );
  NAND2X1 U72981 ( .A(n69898), .B(n70186), .Y(n69899) );
  NOR2X1 U72982 ( .A(n36543), .B(n69899), .Y(n69903) );
  NAND2X1 U72983 ( .A(n70185), .B(n43697), .Y(n69901) );
  NAND2X1 U72984 ( .A(n70184), .B(n43697), .Y(n69900) );
  NAND2X1 U72985 ( .A(n69901), .B(n69900), .Y(n69902) );
  NOR2X1 U72986 ( .A(n69903), .B(n69902), .Y(n69904) );
  XNOR2X1 U72987 ( .A(n69905), .B(n69904), .Y(n69914) );
  XNOR2X1 U72988 ( .A(n69907), .B(n69906), .Y(n69908) );
  XNOR2X1 U72989 ( .A(n42089), .B(n69908), .Y(n69909) );
  MX2X1 U72990 ( .A(n69910), .B(n69909), .S0(n43718), .Y(u_muldiv_result_r[23]) );
  NAND2X1 U72991 ( .A(u_muldiv_mult_result_q[23]), .B(n44632), .Y(n13921) );
  NOR2X1 U72992 ( .A(n69914), .B(n43710), .Y(n69912) );
  NOR2X1 U72993 ( .A(n69912), .B(n69913), .Y(n69915) );
  NAND2X1 U72994 ( .A(n69878), .B(n39301), .Y(n70467) );
  NAND2X1 U72995 ( .A(n69920), .B(n70470), .Y(n69921) );
  XNOR2X1 U72996 ( .A(n43655), .B(n41046), .Y(n70157) );
  INVX1 U72997 ( .A(n69922), .Y(n69932) );
  XNOR2X1 U72998 ( .A(n43633), .B(n69932), .Y(n69923) );
  XNOR2X1 U72999 ( .A(n69923), .B(n39858), .Y(n69924) );
  INVX1 U73000 ( .A(n70452), .Y(n69925) );
  NOR2X1 U73001 ( .A(n41017), .B(n69925), .Y(n69931) );
  NAND2X1 U73002 ( .A(n70452), .B(n43669), .Y(n69929) );
  NAND2X1 U73003 ( .A(n39842), .B(n69929), .Y(n69930) );
  NOR2X1 U73004 ( .A(n69930), .B(n69931), .Y(n70465) );
  XNOR2X1 U73005 ( .A(n69932), .B(n39858), .Y(n69933) );
  XNOR2X1 U73006 ( .A(n70136), .B(n43565), .Y(n69937) );
  XNOR2X1 U73007 ( .A(n39153), .B(n69937), .Y(n69939) );
  INVX1 U73008 ( .A(n69939), .Y(n69938) );
  NAND2X1 U73009 ( .A(n69938), .B(n43623), .Y(n70445) );
  NAND2X1 U73010 ( .A(n69940), .B(n69941), .Y(n69942) );
  XNOR2X1 U73011 ( .A(n43569), .B(n38191), .Y(n69944) );
  NAND2X1 U73012 ( .A(n70116), .B(n43586), .Y(n70239) );
  NAND2X1 U73013 ( .A(n70238), .B(n70239), .Y(n70114) );
  NAND2X1 U73014 ( .A(n70270), .B(n42993), .Y(n70428) );
  INVX1 U73015 ( .A(n70270), .Y(n70265) );
  NAND2X1 U73016 ( .A(n43592), .B(n70265), .Y(n69946) );
  NAND2X1 U73017 ( .A(n69946), .B(n69945), .Y(n70429) );
  NAND2X1 U73018 ( .A(n70086), .B(n40683), .Y(n69950) );
  NAND2X1 U73019 ( .A(n43615), .B(n70084), .Y(n69948) );
  NAND2X1 U73020 ( .A(n69948), .B(n69947), .Y(n69949) );
  NAND2X1 U73021 ( .A(n69950), .B(n69949), .Y(n70262) );
  INVX1 U73022 ( .A(n70262), .Y(n70258) );
  NOR2X1 U73023 ( .A(n69953), .B(n69952), .Y(n69951) );
  NOR2X1 U73024 ( .A(n39556), .B(n69951), .Y(n69956) );
  NAND2X1 U73025 ( .A(n69953), .B(n69952), .Y(n69954) );
  NOR2X1 U73026 ( .A(n70084), .B(n69954), .Y(n69955) );
  NOR2X1 U73027 ( .A(n69956), .B(n69955), .Y(n69958) );
  NAND2X1 U73028 ( .A(n70086), .B(n42998), .Y(n69957) );
  NAND2X1 U73029 ( .A(n69958), .B(n69957), .Y(n70415) );
  INVX1 U73030 ( .A(n70415), .Y(n70412) );
  INVX1 U73031 ( .A(n43000), .Y(n69963) );
  INVX1 U73032 ( .A(n69959), .Y(n69978) );
  XNOR2X1 U73033 ( .A(n72510), .B(n69978), .Y(n69960) );
  XNOR2X1 U73034 ( .A(n69960), .B(n69977), .Y(n69961) );
  XNOR2X1 U73035 ( .A(n69962), .B(n69961), .Y(n69964) );
  NOR2X1 U73036 ( .A(n69963), .B(n69964), .Y(n69972) );
  OR2X1 U73037 ( .A(n41647), .B(n69964), .Y(n69970) );
  XNOR2X1 U73038 ( .A(n69974), .B(n69965), .Y(n69967) );
  NAND2X1 U73039 ( .A(n69967), .B(n69966), .Y(n69968) );
  NAND2X1 U73040 ( .A(n69968), .B(n43000), .Y(n69969) );
  NAND2X1 U73041 ( .A(n69970), .B(n69969), .Y(n69971) );
  NOR2X1 U73042 ( .A(n69972), .B(n69971), .Y(n70407) );
  NAND2X1 U73043 ( .A(n69976), .B(n69975), .Y(n69980) );
  XNOR2X1 U73044 ( .A(n69978), .B(n69977), .Y(n69981) );
  NAND2X1 U73045 ( .A(n72510), .B(n69981), .Y(n69979) );
  NAND2X1 U73046 ( .A(n69980), .B(n69979), .Y(n69984) );
  INVX1 U73047 ( .A(n69981), .Y(n69982) );
  NAND2X1 U73048 ( .A(n69982), .B(n72196), .Y(n69983) );
  NAND2X1 U73049 ( .A(n69984), .B(n69983), .Y(n70273) );
  NAND2X1 U73050 ( .A(n70065), .B(n38950), .Y(n69988) );
  NAND2X1 U73051 ( .A(n39047), .B(n69985), .Y(n69986) );
  NAND2X1 U73052 ( .A(n41731), .B(n69986), .Y(n69987) );
  NAND2X1 U73053 ( .A(n69988), .B(n69987), .Y(n70387) );
  INVX1 U73054 ( .A(n70387), .Y(n70681) );
  NAND2X1 U73055 ( .A(n43486), .B(n44048), .Y(n70381) );
  NAND2X1 U73056 ( .A(n72283), .B(n69989), .Y(n69990) );
  NAND2X1 U73057 ( .A(n71873), .B(n69990), .Y(n71877) );
  XNOR2X1 U73058 ( .A(n70299), .B(n41694), .Y(n70623) );
  INVX1 U73059 ( .A(n70623), .Y(n70303) );
  NAND2X1 U73060 ( .A(n43991), .B(n43607), .Y(n70316) );
  INVX1 U73061 ( .A(n70316), .Y(n70301) );
  NAND2X1 U73062 ( .A(n69991), .B(n43604), .Y(n72328) );
  INVX1 U73063 ( .A(n72328), .Y(n72263) );
  XNOR2X1 U73064 ( .A(n70301), .B(n72263), .Y(n69995) );
  NAND2X1 U73065 ( .A(n69993), .B(n69992), .Y(n69994) );
  NAND2X1 U73066 ( .A(n72326), .B(n69994), .Y(n70302) );
  INVX1 U73067 ( .A(n70302), .Y(n70307) );
  XNOR2X1 U73068 ( .A(n69995), .B(n70307), .Y(n69996) );
  XNOR2X1 U73069 ( .A(n41695), .B(n69996), .Y(n70002) );
  XNOR2X1 U73070 ( .A(n41692), .B(n69997), .Y(n70003) );
  INVX1 U73071 ( .A(n70003), .Y(n69998) );
  NAND2X1 U73072 ( .A(n72355), .B(n69998), .Y(n70000) );
  NAND2X1 U73073 ( .A(n72355), .B(n70004), .Y(n69999) );
  NAND2X1 U73074 ( .A(n70000), .B(n69999), .Y(n70314) );
  INVX1 U73075 ( .A(n70314), .Y(n70001) );
  XNOR2X1 U73076 ( .A(n70002), .B(n70001), .Y(n70009) );
  NAND2X1 U73077 ( .A(n70003), .B(n72268), .Y(n70005) );
  NOR2X1 U73078 ( .A(n70005), .B(n70004), .Y(n70007) );
  NOR2X1 U73079 ( .A(n70007), .B(n70006), .Y(n70008) );
  XNOR2X1 U73080 ( .A(n70009), .B(n70008), .Y(n70294) );
  XNOR2X1 U73081 ( .A(n70294), .B(n41528), .Y(n70015) );
  INVX1 U73082 ( .A(n70010), .Y(n70287) );
  NAND2X1 U73083 ( .A(n70012), .B(n70011), .Y(n70013) );
  NAND2X1 U73084 ( .A(n70287), .B(n70013), .Y(n70014) );
  NAND2X1 U73085 ( .A(n70285), .B(n70286), .Y(n70284) );
  NAND2X1 U73086 ( .A(n70014), .B(n70284), .Y(n70296) );
  INVX1 U73087 ( .A(n70331), .Y(n70327) );
  INVX1 U73088 ( .A(n70021), .Y(n70322) );
  NAND2X1 U73089 ( .A(n70322), .B(n70323), .Y(n70321) );
  INVX1 U73090 ( .A(n70016), .Y(n70324) );
  NAND2X1 U73091 ( .A(n70020), .B(n70021), .Y(n70017) );
  NAND2X1 U73092 ( .A(n70324), .B(n70017), .Y(n70018) );
  NAND2X1 U73093 ( .A(n70321), .B(n70018), .Y(n70330) );
  NAND2X1 U73094 ( .A(n44007), .B(n43500), .Y(n70320) );
  INVX1 U73095 ( .A(n70345), .Y(n70342) );
  XNOR2X1 U73096 ( .A(n70320), .B(n70342), .Y(n70019) );
  XNOR2X1 U73097 ( .A(n70336), .B(n70019), .Y(n70029) );
  XNOR2X1 U73098 ( .A(n70021), .B(n70020), .Y(n70022) );
  XNOR2X1 U73099 ( .A(n70324), .B(n70022), .Y(n70024) );
  NAND2X1 U73100 ( .A(n70024), .B(n70023), .Y(n70028) );
  INVX1 U73101 ( .A(n70023), .Y(n70031) );
  INVX1 U73102 ( .A(n70024), .Y(n70025) );
  NAND2X1 U73103 ( .A(n70031), .B(n70025), .Y(n70026) );
  NAND2X1 U73104 ( .A(n42033), .B(n70026), .Y(n70027) );
  NAND2X1 U73105 ( .A(n70028), .B(n70027), .Y(n70338) );
  INVX1 U73106 ( .A(n70338), .Y(n70341) );
  XNOR2X1 U73107 ( .A(n70029), .B(n70341), .Y(n70355) );
  NAND2X1 U73108 ( .A(n41492), .B(n70033), .Y(n70034) );
  NAND2X1 U73109 ( .A(n41529), .B(n41492), .Y(n70032) );
  NAND2X1 U73110 ( .A(n43491), .B(n44025), .Y(n70360) );
  NOR2X1 U73111 ( .A(n36780), .B(n70360), .Y(n70038) );
  NAND2X1 U73112 ( .A(n70032), .B(n70360), .Y(n70036) );
  NAND2X1 U73113 ( .A(n41529), .B(n70033), .Y(n70353) );
  NAND2X1 U73114 ( .A(n70034), .B(n70353), .Y(n70035) );
  NOR2X1 U73115 ( .A(n70036), .B(n70035), .Y(n70037) );
  NOR2X1 U73116 ( .A(n70038), .B(n70037), .Y(n70040) );
  OR2X1 U73117 ( .A(n70360), .B(n70353), .Y(n70039) );
  NAND2X1 U73118 ( .A(n70040), .B(n70039), .Y(n70041) );
  XNOR2X1 U73119 ( .A(n70355), .B(n70041), .Y(n70280) );
  INVX1 U73120 ( .A(n70280), .Y(n70380) );
  XNOR2X1 U73121 ( .A(n70381), .B(n70380), .Y(n70050) );
  INVX1 U73122 ( .A(n70042), .Y(n70045) );
  NAND2X1 U73123 ( .A(n38264), .B(n70043), .Y(n70044) );
  NAND2X1 U73124 ( .A(n70045), .B(n70044), .Y(n70049) );
  NAND2X1 U73125 ( .A(n70047), .B(n70046), .Y(n70048) );
  NAND2X1 U73126 ( .A(n70049), .B(n70048), .Y(n70281) );
  INVX1 U73127 ( .A(n70281), .Y(n70379) );
  XNOR2X1 U73128 ( .A(n70050), .B(n70379), .Y(n70368) );
  NAND2X1 U73129 ( .A(n43614), .B(n43477), .Y(n72208) );
  INVX1 U73130 ( .A(n72208), .Y(n72212) );
  XNOR2X1 U73131 ( .A(n41730), .B(n72212), .Y(n70063) );
  INVX1 U73132 ( .A(n70055), .Y(n70053) );
  NAND2X1 U73133 ( .A(n70053), .B(n70052), .Y(n70062) );
  INVX1 U73134 ( .A(n70054), .Y(n70060) );
  NAND2X1 U73135 ( .A(n70056), .B(n44024), .Y(n70057) );
  NAND2X1 U73136 ( .A(n70060), .B(n70059), .Y(n70061) );
  NAND2X1 U73137 ( .A(n70062), .B(n70061), .Y(n70369) );
  INVX1 U73138 ( .A(n70369), .Y(n70385) );
  XNOR2X1 U73139 ( .A(n70063), .B(n70385), .Y(n70064) );
  XNOR2X1 U73140 ( .A(n70065), .B(n41731), .Y(n70066) );
  XNOR2X1 U73141 ( .A(n39047), .B(n70066), .Y(n70395) );
  INVX1 U73142 ( .A(n70395), .Y(n70070) );
  NAND2X1 U73143 ( .A(n72200), .B(n70068), .Y(n70067) );
  NOR2X1 U73144 ( .A(n70070), .B(n70067), .Y(n70075) );
  NOR2X1 U73145 ( .A(n72200), .B(n70069), .Y(n70071) );
  NAND2X1 U73146 ( .A(n70071), .B(n70070), .Y(n70072) );
  NAND2X1 U73147 ( .A(n70073), .B(n70072), .Y(n70074) );
  NOR2X1 U73148 ( .A(n70075), .B(n70074), .Y(n70076) );
  XNOR2X1 U73149 ( .A(n41468), .B(n70076), .Y(n70404) );
  XNOR2X1 U73150 ( .A(n70077), .B(n70404), .Y(n70078) );
  XOR2X1 U73151 ( .A(n70273), .B(n70078), .Y(n70259) );
  XNOR2X1 U73152 ( .A(n70407), .B(n70259), .Y(n70409) );
  XNOR2X1 U73153 ( .A(n43602), .B(n39556), .Y(n70079) );
  XNOR2X1 U73154 ( .A(n70079), .B(n43616), .Y(n70080) );
  XNOR2X1 U73155 ( .A(n70409), .B(n70080), .Y(n70081) );
  XNOR2X1 U73156 ( .A(n70412), .B(n70081), .Y(n70094) );
  NAND2X1 U73157 ( .A(n70082), .B(n70087), .Y(n70083) );
  NOR2X1 U73158 ( .A(n70084), .B(n70083), .Y(n70093) );
  NOR2X1 U73159 ( .A(n43601), .B(n70085), .Y(n70091) );
  NAND2X1 U73160 ( .A(n70086), .B(n43598), .Y(n70089) );
  NAND2X1 U73161 ( .A(n70087), .B(n43598), .Y(n70088) );
  NAND2X1 U73162 ( .A(n70089), .B(n70088), .Y(n70090) );
  OR2X1 U73163 ( .A(n70091), .B(n70090), .Y(n70092) );
  NOR2X1 U73164 ( .A(n70093), .B(n70092), .Y(n70423) );
  XNOR2X1 U73165 ( .A(n70094), .B(n70423), .Y(n70095) );
  NAND2X1 U73166 ( .A(n39306), .B(n42997), .Y(n70100) );
  NAND2X1 U73167 ( .A(n43617), .B(n70096), .Y(n70098) );
  NAND2X1 U73168 ( .A(n70098), .B(n70097), .Y(n70099) );
  NAND2X1 U73169 ( .A(n70100), .B(n70099), .Y(n70269) );
  INVX1 U73170 ( .A(n70269), .Y(n70264) );
  NOR2X1 U73171 ( .A(n43618), .B(n70270), .Y(n70101) );
  NAND2X1 U73172 ( .A(n70264), .B(n70101), .Y(n70104) );
  NOR2X1 U73173 ( .A(n70265), .B(n42996), .Y(n70102) );
  NAND2X1 U73174 ( .A(n70102), .B(n70269), .Y(n70103) );
  NAND2X1 U73175 ( .A(n70104), .B(n70103), .Y(n70105) );
  INVX1 U73176 ( .A(n71079), .Y(n72353) );
  XNOR2X1 U73177 ( .A(n70105), .B(n72353), .Y(n70106) );
  XNOR2X1 U73178 ( .A(n70578), .B(n70106), .Y(n70107) );
  XNOR2X1 U73179 ( .A(n41419), .B(n70107), .Y(n70242) );
  XNOR2X1 U73180 ( .A(n70242), .B(n43582), .Y(n70112) );
  INVX1 U73181 ( .A(n70109), .Y(n70108) );
  NAND2X1 U73182 ( .A(n43568), .B(n70109), .Y(n70255) );
  NAND2X1 U73183 ( .A(n70111), .B(n70110), .Y(n70254) );
  XNOR2X1 U73184 ( .A(n70112), .B(n39886), .Y(n70237) );
  XNOR2X1 U73185 ( .A(n43574), .B(n70237), .Y(n70113) );
  XNOR2X1 U73186 ( .A(n70114), .B(n70113), .Y(n70219) );
  AND2X1 U73187 ( .A(n70117), .B(n70116), .Y(n70119) );
  NOR2X1 U73188 ( .A(n41143), .B(n41149), .Y(n70120) );
  NAND2X1 U73189 ( .A(n70119), .B(n39958), .Y(n70220) );
  NAND2X1 U73190 ( .A(n70120), .B(n70220), .Y(n70121) );
  XNOR2X1 U73191 ( .A(n70121), .B(n43537), .Y(n70122) );
  XNOR2X1 U73192 ( .A(n70219), .B(n70122), .Y(n70134) );
  INVX1 U73193 ( .A(n70136), .Y(n70135) );
  NAND2X1 U73194 ( .A(n70124), .B(n70123), .Y(n70130) );
  INVX1 U73195 ( .A(n70130), .Y(n70126) );
  NAND2X1 U73196 ( .A(n70128), .B(n70127), .Y(n70218) );
  NAND2X1 U73197 ( .A(n70130), .B(n70129), .Y(n70132) );
  NAND2X1 U73198 ( .A(n70132), .B(n70131), .Y(n70133) );
  INVX1 U73199 ( .A(n70233), .Y(n70539) );
  XNOR2X1 U73200 ( .A(n70134), .B(n70539), .Y(n70230) );
  XNOR2X1 U73201 ( .A(n71794), .B(n43546), .Y(n70439) );
  NAND2X1 U73202 ( .A(n70135), .B(n39629), .Y(n70141) );
  NAND2X1 U73203 ( .A(n43562), .B(n70136), .Y(n70140) );
  NAND2X1 U73204 ( .A(n70138), .B(n70137), .Y(n70139) );
  NAND2X1 U73205 ( .A(n70140), .B(n70139), .Y(n70223) );
  XNOR2X1 U73206 ( .A(n70439), .B(n41104), .Y(n70142) );
  XNOR2X1 U73207 ( .A(n70230), .B(n70142), .Y(n70143) );
  XNOR2X1 U73208 ( .A(n41101), .B(n70143), .Y(n70215) );
  NAND2X1 U73209 ( .A(n70145), .B(n43548), .Y(n70155) );
  INVX1 U73210 ( .A(n70145), .Y(n70148) );
  NOR2X1 U73211 ( .A(n70148), .B(n70147), .Y(n70146) );
  NOR2X1 U73212 ( .A(n70146), .B(n43552), .Y(n70150) );
  NAND2X1 U73213 ( .A(n70148), .B(n70147), .Y(n70149) );
  NAND2X1 U73214 ( .A(n70150), .B(n70149), .Y(n70154) );
  NAND2X1 U73215 ( .A(n70152), .B(n70151), .Y(n70153) );
  XNOR2X1 U73216 ( .A(n70762), .B(n70458), .Y(n70156) );
  XNOR2X1 U73217 ( .A(n70157), .B(n70471), .Y(n70163) );
  NOR2X1 U73218 ( .A(n39511), .B(n41266), .Y(n70160) );
  NAND2X1 U73219 ( .A(n70209), .B(n43658), .Y(n70511) );
  NAND2X1 U73220 ( .A(n70472), .B(n70161), .Y(n70512) );
  NOR2X1 U73221 ( .A(n39331), .B(n38557), .Y(n70162) );
  XNOR2X1 U73222 ( .A(n70163), .B(n70162), .Y(n70836) );
  NAND2X1 U73223 ( .A(n70165), .B(n70164), .Y(n70477) );
  NOR2X1 U73224 ( .A(n70478), .B(n70166), .Y(n70170) );
  NAND2X1 U73225 ( .A(n70478), .B(n70210), .Y(n70168) );
  NOR2X1 U73226 ( .A(n43526), .B(n70168), .Y(n70169) );
  NOR2X1 U73227 ( .A(n70170), .B(n70169), .Y(n70171) );
  XNOR2X1 U73228 ( .A(n43509), .B(n38048), .Y(n70180) );
  NAND2X1 U73229 ( .A(n70172), .B(n43682), .Y(n70173) );
  NOR2X1 U73230 ( .A(n39906), .B(n70173), .Y(n70176) );
  NOR2X1 U73231 ( .A(n70479), .B(n70174), .Y(n70175) );
  NOR2X1 U73232 ( .A(n70176), .B(n70175), .Y(n70177) );
  NOR2X1 U73233 ( .A(n38046), .B(n70177), .Y(n70179) );
  XNOR2X1 U73234 ( .A(n70180), .B(n41089), .Y(n70183) );
  NOR2X1 U73235 ( .A(n41339), .B(n70207), .Y(n70182) );
  XNOR2X1 U73236 ( .A(n70183), .B(n70182), .Y(n70203) );
  XNOR2X1 U73237 ( .A(n70203), .B(n43692), .Y(n70192) );
  NOR2X1 U73238 ( .A(n39005), .B(n36543), .Y(n70189) );
  NOR2X1 U73239 ( .A(n70187), .B(n41164), .Y(n70188) );
  NAND2X1 U73240 ( .A(n71130), .B(n71129), .Y(n70204) );
  NOR2X1 U73241 ( .A(n36541), .B(n70204), .Y(n70191) );
  XNOR2X1 U73242 ( .A(n70192), .B(n70191), .Y(n70200) );
  XNOR2X1 U73243 ( .A(n70200), .B(n43708), .Y(n70193) );
  XNOR2X1 U73244 ( .A(n38032), .B(n70193), .Y(n70198) );
  XNOR2X1 U73245 ( .A(n70195), .B(n70194), .Y(n70196) );
  XNOR2X1 U73246 ( .A(n42097), .B(n70196), .Y(n70197) );
  NAND2X1 U73247 ( .A(u_muldiv_mult_result_q[24]), .B(n44631), .Y(n13913) );
  NAND2X1 U73248 ( .A(n70200), .B(n43710), .Y(n70199) );
  INVX1 U73249 ( .A(n70203), .Y(n70202) );
  NAND2X1 U73250 ( .A(n70202), .B(n43697), .Y(n71128) );
  NAND2X1 U73251 ( .A(n43691), .B(n70203), .Y(n71132) );
  XNOR2X1 U73252 ( .A(n38048), .B(n41089), .Y(n70208) );
  NAND2X1 U73253 ( .A(n43505), .B(n70208), .Y(n70783) );
  NAND2X1 U73254 ( .A(n70783), .B(n70785), .Y(n70790) );
  NAND2X1 U73255 ( .A(n70211), .B(n70210), .Y(n70767) );
  NAND2X1 U73256 ( .A(n70836), .B(n43528), .Y(n70213) );
  NAND2X1 U73257 ( .A(n40405), .B(n70213), .Y(n70214) );
  INVX1 U73258 ( .A(n70217), .Y(n70216) );
  NAND2X1 U73259 ( .A(n43631), .B(n70216), .Y(n70516) );
  NAND2X1 U73260 ( .A(n70516), .B(n70517), .Y(n70534) );
  XNOR2X1 U73261 ( .A(n70218), .B(n72149), .Y(n70221) );
  INVX1 U73262 ( .A(n70537), .Y(n70536) );
  XNOR2X1 U73263 ( .A(n70221), .B(n70536), .Y(n70442) );
  XNOR2X1 U73264 ( .A(n43627), .B(n70442), .Y(n70222) );
  XOR2X1 U73265 ( .A(n70223), .B(n70222), .Y(n70225) );
  NAND2X1 U73266 ( .A(n70225), .B(n43548), .Y(n70224) );
  XNOR2X1 U73267 ( .A(n41101), .B(n70225), .Y(n70226) );
  NAND2X1 U73268 ( .A(n43544), .B(n70226), .Y(n70227) );
  NAND2X1 U73269 ( .A(n70228), .B(n70227), .Y(n70546) );
  INVX1 U73270 ( .A(n70230), .Y(n70229) );
  NAND2X1 U73271 ( .A(n43562), .B(n70229), .Y(n70549) );
  NAND2X1 U73272 ( .A(n70230), .B(n39629), .Y(n70231) );
  NAND2X1 U73273 ( .A(n41104), .B(n70231), .Y(n70548) );
  NOR2X1 U73274 ( .A(n43536), .B(n70537), .Y(n70232) );
  NAND2X1 U73275 ( .A(n70539), .B(n70232), .Y(n70236) );
  NOR2X1 U73276 ( .A(n70536), .B(n43541), .Y(n70234) );
  NAND2X1 U73277 ( .A(n70234), .B(n70233), .Y(n70235) );
  NAND2X1 U73278 ( .A(n70236), .B(n70235), .Y(n70755) );
  NAND2X1 U73279 ( .A(n70239), .B(n70238), .Y(n70244) );
  INVX1 U73280 ( .A(n70901), .Y(n70241) );
  NAND2X1 U73281 ( .A(n70562), .B(n43573), .Y(n70243) );
  NOR2X1 U73282 ( .A(n36604), .B(n70243), .Y(n70246) );
  NOR2X1 U73283 ( .A(n43573), .B(n70244), .Y(n70245) );
  NOR2X1 U73284 ( .A(n70246), .B(n70245), .Y(n70253) );
  INVX1 U73285 ( .A(n70562), .Y(n70247) );
  NAND2X1 U73286 ( .A(n70247), .B(n43573), .Y(n70251) );
  NAND2X1 U73287 ( .A(n39862), .B(n43573), .Y(n70249) );
  NAND2X1 U73288 ( .A(n70249), .B(n70562), .Y(n70250) );
  NAND2X1 U73289 ( .A(n70251), .B(n70250), .Y(n70252) );
  NAND2X1 U73290 ( .A(n70253), .B(n70252), .Y(n70437) );
  NAND2X1 U73291 ( .A(n43568), .B(n70578), .Y(n70744) );
  NAND2X1 U73292 ( .A(n70255), .B(n70254), .Y(n70256) );
  NAND2X1 U73293 ( .A(n43567), .B(n70256), .Y(n70743) );
  NAND2X1 U73294 ( .A(n70572), .B(n70743), .Y(n70257) );
  NOR2X1 U73295 ( .A(n38142), .B(n70257), .Y(n70436) );
  NAND2X1 U73296 ( .A(n70258), .B(n43616), .Y(n70567) );
  XNOR2X1 U73297 ( .A(n38873), .B(n39556), .Y(n70260) );
  XNOR2X1 U73298 ( .A(n70260), .B(n70259), .Y(n70261) );
  XNOR2X1 U73299 ( .A(n70412), .B(n70261), .Y(n70420) );
  INVX1 U73300 ( .A(n70420), .Y(n70421) );
  NAND2X1 U73301 ( .A(n43615), .B(n70420), .Y(n70568) );
  NAND2X1 U73302 ( .A(n70263), .B(n70568), .Y(n70728) );
  NOR2X1 U73303 ( .A(n70265), .B(n70264), .Y(n70266) );
  NOR2X1 U73304 ( .A(n70266), .B(n42997), .Y(n70268) );
  NOR2X1 U73305 ( .A(n38302), .B(n42995), .Y(n70267) );
  NOR2X1 U73306 ( .A(n70270), .B(n70269), .Y(n70271) );
  INVX1 U73307 ( .A(n70733), .Y(n70735) );
  XNOR2X1 U73308 ( .A(n70728), .B(n70735), .Y(n70426) );
  INVX1 U73309 ( .A(n70272), .Y(n71819) );
  XNOR2X1 U73310 ( .A(n43618), .B(n43616), .Y(n70569) );
  INVX1 U73311 ( .A(n70569), .Y(n72358) );
  XNOR2X1 U73312 ( .A(n71819), .B(n72358), .Y(n70424) );
  NAND2X1 U73313 ( .A(n72510), .B(n70404), .Y(n70277) );
  INVX1 U73314 ( .A(n70273), .Y(n70275) );
  INVX1 U73315 ( .A(n70404), .Y(n70405) );
  NAND2X1 U73316 ( .A(n70405), .B(n72196), .Y(n70274) );
  NAND2X1 U73317 ( .A(n70275), .B(n70274), .Y(n70276) );
  AND2X1 U73318 ( .A(n70277), .B(n70276), .Y(n70933) );
  INVX1 U73319 ( .A(n70381), .Y(n70279) );
  NAND2X1 U73320 ( .A(n70379), .B(n70380), .Y(n70278) );
  NAND2X1 U73321 ( .A(n70279), .B(n70278), .Y(n70283) );
  NAND2X1 U73322 ( .A(n70281), .B(n70280), .Y(n70282) );
  NAND2X1 U73323 ( .A(n70283), .B(n70282), .Y(n70616) );
  INVX1 U73324 ( .A(n70284), .Y(n70291) );
  NAND2X1 U73325 ( .A(n70287), .B(n70285), .Y(n70289) );
  NAND2X1 U73326 ( .A(n70287), .B(n70286), .Y(n70288) );
  NAND2X1 U73327 ( .A(n70289), .B(n70288), .Y(n70290) );
  NOR2X1 U73328 ( .A(n70291), .B(n70290), .Y(n70292) );
  NAND2X1 U73329 ( .A(n70294), .B(n70292), .Y(n70293) );
  NAND2X1 U73330 ( .A(n41528), .B(n70293), .Y(n70298) );
  INVX1 U73331 ( .A(n70294), .Y(n70295) );
  NAND2X1 U73332 ( .A(n70296), .B(n70295), .Y(n70297) );
  NAND2X1 U73333 ( .A(n70298), .B(n70297), .Y(n71014) );
  NAND2X1 U73334 ( .A(n72326), .B(n70299), .Y(n70300) );
  NAND2X1 U73335 ( .A(n71878), .B(n70300), .Y(n71882) );
  XNOR2X1 U73336 ( .A(n70303), .B(n41696), .Y(n70627) );
  INVX1 U73337 ( .A(n70627), .Y(n70995) );
  NAND2X1 U73338 ( .A(n43999), .B(n43607), .Y(n70640) );
  INVX1 U73339 ( .A(n70640), .Y(n70626) );
  NAND2X1 U73340 ( .A(n70301), .B(n43603), .Y(n72356) );
  INVX1 U73341 ( .A(n72356), .Y(n72422) );
  XNOR2X1 U73342 ( .A(n70626), .B(n72422), .Y(n70305) );
  NAND2X1 U73343 ( .A(n70303), .B(n70302), .Y(n70304) );
  NAND2X1 U73344 ( .A(n72355), .B(n70304), .Y(n70628) );
  INVX1 U73345 ( .A(n70628), .Y(n70632) );
  XNOR2X1 U73346 ( .A(n70305), .B(n70632), .Y(n70306) );
  XNOR2X1 U73347 ( .A(n41697), .B(n70306), .Y(n70311) );
  XNOR2X1 U73348 ( .A(n41695), .B(n70307), .Y(n70312) );
  NAND2X1 U73349 ( .A(n72263), .B(n70312), .Y(n70309) );
  NAND2X1 U73350 ( .A(n72263), .B(n70314), .Y(n70308) );
  NAND2X1 U73351 ( .A(n70309), .B(n70308), .Y(n70638) );
  INVX1 U73352 ( .A(n70638), .Y(n70310) );
  XNOR2X1 U73353 ( .A(n70311), .B(n70310), .Y(n70319) );
  INVX1 U73354 ( .A(n70312), .Y(n70313) );
  NAND2X1 U73355 ( .A(n70313), .B(n72328), .Y(n70315) );
  NOR2X1 U73356 ( .A(n70315), .B(n70314), .Y(n70317) );
  NOR2X1 U73357 ( .A(n70317), .B(n70316), .Y(n70318) );
  XNOR2X1 U73358 ( .A(n70319), .B(n70318), .Y(n71013) );
  INVX1 U73359 ( .A(n70646), .Y(n70650) );
  INVX1 U73360 ( .A(n70320), .Y(n70337) );
  NAND2X1 U73361 ( .A(n70324), .B(n70322), .Y(n70326) );
  NAND2X1 U73362 ( .A(n70324), .B(n70323), .Y(n70325) );
  NAND2X1 U73363 ( .A(n70328), .B(n70327), .Y(n70329) );
  NAND2X1 U73364 ( .A(n70337), .B(n70329), .Y(n70333) );
  NAND2X1 U73365 ( .A(n70331), .B(n70330), .Y(n70332) );
  NAND2X1 U73366 ( .A(n70333), .B(n70332), .Y(n70651) );
  NOR2X1 U73367 ( .A(n43503), .B(n44022), .Y(n70334) );
  XNOR2X1 U73368 ( .A(n70651), .B(n70334), .Y(n70335) );
  XNOR2X1 U73369 ( .A(n70650), .B(n70335), .Y(n70660) );
  INVX1 U73370 ( .A(n70340), .Y(n70339) );
  NAND2X1 U73371 ( .A(n70339), .B(n70338), .Y(n70608) );
  NAND2X1 U73372 ( .A(n43496), .B(n44024), .Y(n70609) );
  NAND2X1 U73373 ( .A(n70608), .B(n70609), .Y(n70344) );
  NAND2X1 U73374 ( .A(n70341), .B(n70340), .Y(n70346) );
  NAND2X1 U73375 ( .A(n70342), .B(n70346), .Y(n70607) );
  INVX1 U73376 ( .A(n70607), .Y(n70343) );
  NOR2X1 U73377 ( .A(n70344), .B(n70343), .Y(n70351) );
  OR2X1 U73378 ( .A(n70609), .B(n70608), .Y(n70349) );
  NOR2X1 U73379 ( .A(n70345), .B(n70609), .Y(n70347) );
  NAND2X1 U73380 ( .A(n70347), .B(n70346), .Y(n70348) );
  NAND2X1 U73381 ( .A(n70349), .B(n70348), .Y(n70350) );
  NOR2X1 U73382 ( .A(n70351), .B(n70350), .Y(n70352) );
  XOR2X1 U73383 ( .A(n70660), .B(n70352), .Y(n70613) );
  NAND2X1 U73384 ( .A(n36780), .B(n70353), .Y(n70354) );
  NAND2X1 U73385 ( .A(n70355), .B(n70354), .Y(n70606) );
  NAND2X1 U73386 ( .A(n43491), .B(n44047), .Y(n70359) );
  NAND2X1 U73387 ( .A(n70606), .B(n70359), .Y(n70358) );
  INVX1 U73388 ( .A(n70360), .Y(n70356) );
  NAND2X1 U73389 ( .A(n70356), .B(n70361), .Y(n70605) );
  INVX1 U73390 ( .A(n70605), .Y(n70357) );
  NOR2X1 U73391 ( .A(n70358), .B(n70357), .Y(n70366) );
  OR2X1 U73392 ( .A(n70359), .B(n70606), .Y(n70364) );
  NOR2X1 U73393 ( .A(n70360), .B(n70359), .Y(n70362) );
  NAND2X1 U73394 ( .A(n70362), .B(n70361), .Y(n70363) );
  NAND2X1 U73395 ( .A(n70364), .B(n70363), .Y(n70365) );
  XNOR2X1 U73396 ( .A(n70367), .B(n41733), .Y(n70601) );
  INVX1 U73397 ( .A(n70601), .Y(n70598) );
  NAND2X1 U73398 ( .A(n70385), .B(n70368), .Y(n70374) );
  NAND2X1 U73399 ( .A(n41730), .B(n70374), .Y(n70596) );
  INVX1 U73400 ( .A(n70596), .Y(n70373) );
  INVX1 U73401 ( .A(n70368), .Y(n70370) );
  NAND2X1 U73402 ( .A(n70370), .B(n70369), .Y(n70597) );
  NAND2X1 U73403 ( .A(n43614), .B(n43482), .Y(n72219) );
  NAND2X1 U73404 ( .A(n70597), .B(n72219), .Y(n70372) );
  NOR2X1 U73405 ( .A(n70373), .B(n70372), .Y(n70377) );
  INVX1 U73406 ( .A(n70374), .Y(n70375) );
  NOR2X1 U73407 ( .A(n70375), .B(n72219), .Y(n70376) );
  NOR2X1 U73408 ( .A(n70377), .B(n70376), .Y(n70378) );
  XNOR2X1 U73409 ( .A(n70598), .B(n70378), .Y(n70677) );
  INVX1 U73410 ( .A(n70677), .Y(n70678) );
  XNOR2X1 U73411 ( .A(n70380), .B(n70379), .Y(n70383) );
  XNOR2X1 U73412 ( .A(n70381), .B(n41730), .Y(n70382) );
  XNOR2X1 U73413 ( .A(n70383), .B(n70382), .Y(n70384) );
  XNOR2X1 U73414 ( .A(n70385), .B(n70384), .Y(n70679) );
  INVX1 U73415 ( .A(n70679), .Y(n70386) );
  NAND2X1 U73416 ( .A(n70386), .B(n72208), .Y(n70682) );
  INVX1 U73417 ( .A(n70682), .Y(n70391) );
  NOR2X1 U73418 ( .A(n70681), .B(n72212), .Y(n70389) );
  NOR2X1 U73419 ( .A(n70679), .B(n70387), .Y(n70388) );
  NOR2X1 U73420 ( .A(n70389), .B(n70388), .Y(n70390) );
  NOR2X1 U73421 ( .A(n70391), .B(n70390), .Y(n70392) );
  XNOR2X1 U73422 ( .A(n70678), .B(n70392), .Y(n70704) );
  NOR2X1 U73423 ( .A(n70395), .B(n72202), .Y(n70394) );
  NOR2X1 U73424 ( .A(n70394), .B(n70393), .Y(n70691) );
  NAND2X1 U73425 ( .A(n70395), .B(n72202), .Y(n70692) );
  NAND2X1 U73426 ( .A(n70692), .B(n72202), .Y(n70396) );
  NOR2X1 U73427 ( .A(n70691), .B(n70396), .Y(n70397) );
  NAND2X1 U73428 ( .A(n70397), .B(n41468), .Y(n70400) );
  NOR2X1 U73429 ( .A(n37389), .B(n72202), .Y(n70398) );
  NAND2X1 U73430 ( .A(n70398), .B(n70691), .Y(n70399) );
  NAND2X1 U73431 ( .A(n70400), .B(n70399), .Y(n70401) );
  XNOR2X1 U73432 ( .A(n70401), .B(n71582), .Y(n70402) );
  XNOR2X1 U73433 ( .A(n70704), .B(n70402), .Y(n70403) );
  XNOR2X1 U73434 ( .A(n70933), .B(n70403), .Y(n70716) );
  NAND2X1 U73435 ( .A(n72515), .B(n70404), .Y(n70706) );
  NAND2X1 U73436 ( .A(n70405), .B(n43000), .Y(n70406) );
  NAND2X1 U73437 ( .A(n38873), .B(n70406), .Y(n70705) );
  XNOR2X1 U73438 ( .A(n70717), .B(n39556), .Y(n70408) );
  XNOR2X1 U73439 ( .A(n70716), .B(n70408), .Y(n70589) );
  NAND2X1 U73440 ( .A(n39556), .B(n70409), .Y(n70588) );
  NAND2X1 U73441 ( .A(n70588), .B(n43597), .Y(n70414) );
  INVX1 U73442 ( .A(n70409), .Y(n70410) );
  NAND2X1 U73443 ( .A(n70410), .B(n42999), .Y(n70411) );
  NAND2X1 U73444 ( .A(n70412), .B(n70411), .Y(n70587) );
  INVX1 U73445 ( .A(n70587), .Y(n70413) );
  NOR2X1 U73446 ( .A(n70414), .B(n70413), .Y(n70419) );
  NOR2X1 U73447 ( .A(n43597), .B(n70415), .Y(n70417) );
  NOR2X1 U73448 ( .A(n43597), .B(n70588), .Y(n70416) );
  OR2X1 U73449 ( .A(n70417), .B(n70416), .Y(n70418) );
  NAND2X1 U73450 ( .A(n70421), .B(n43597), .Y(n70422) );
  XNOR2X1 U73451 ( .A(n70729), .B(n38938), .Y(n70583) );
  INVX1 U73452 ( .A(n70583), .Y(n70582) );
  XNOR2X1 U73453 ( .A(n70424), .B(n70582), .Y(n70425) );
  XNOR2X1 U73454 ( .A(n70426), .B(n70425), .Y(n70435) );
  NAND2X1 U73455 ( .A(n43592), .B(n38302), .Y(n70427) );
  NOR2X1 U73456 ( .A(n70427), .B(n70429), .Y(n70433) );
  NAND2X1 U73457 ( .A(n70428), .B(n42994), .Y(n70431) );
  NAND2X1 U73458 ( .A(n70578), .B(n70429), .Y(n70430) );
  NOR2X1 U73459 ( .A(n70431), .B(n70430), .Y(n70432) );
  NOR2X1 U73460 ( .A(n70433), .B(n70432), .Y(n70434) );
  XNOR2X1 U73461 ( .A(n70437), .B(n41193), .Y(n70438) );
  XNOR2X1 U73462 ( .A(n70755), .B(n70440), .Y(n70441) );
  XNOR2X1 U73463 ( .A(n40986), .B(n70441), .Y(n70530) );
  INVX1 U73464 ( .A(n70446), .Y(n70443) );
  NAND2X1 U73465 ( .A(n43619), .B(n70443), .Y(n70448) );
  NAND2X1 U73466 ( .A(n70448), .B(n70447), .Y(n70555) );
  XNOR2X1 U73467 ( .A(n70555), .B(n43633), .Y(n70449) );
  XNOR2X1 U73468 ( .A(n70530), .B(n70449), .Y(n70450) );
  XNOR2X1 U73469 ( .A(n38898), .B(n70450), .Y(n70526) );
  XNOR2X1 U73470 ( .A(n70762), .B(n70526), .Y(n70451) );
  XOR2X1 U73471 ( .A(n70534), .B(n70451), .Y(n70775) );
  NOR2X1 U73472 ( .A(n70453), .B(n38208), .Y(n70454) );
  NOR2X1 U73473 ( .A(n70454), .B(n38555), .Y(n70455) );
  NOR2X1 U73474 ( .A(n69925), .B(n70455), .Y(n70456) );
  INVX1 U73475 ( .A(n70458), .Y(n70462) );
  XNOR2X1 U73476 ( .A(n70462), .B(n38422), .Y(n70460) );
  NAND2X1 U73477 ( .A(n70771), .B(n70770), .Y(n70528) );
  NAND2X1 U73478 ( .A(n69878), .B(n70470), .Y(n70461) );
  XNOR2X1 U73479 ( .A(n43667), .B(n70462), .Y(n70463) );
  XNOR2X1 U73480 ( .A(n70463), .B(n38422), .Y(n70464) );
  XNOR2X1 U73481 ( .A(n70465), .B(n70464), .Y(n70468) );
  INVX1 U73482 ( .A(n70468), .Y(n70466) );
  INVX1 U73483 ( .A(n70467), .Y(n70469) );
  NAND2X1 U73484 ( .A(n70776), .B(n41042), .Y(n70524) );
  XNOR2X1 U73485 ( .A(n41046), .B(n70471), .Y(n70475) );
  INVX1 U73486 ( .A(n70472), .Y(n70473) );
  NOR2X1 U73487 ( .A(n39362), .B(n70473), .Y(n70474) );
  NAND2X1 U73488 ( .A(n70513), .B(n70829), .Y(n70509) );
  XNOR2X1 U73489 ( .A(n72586), .B(n40162), .Y(n70476) );
  XNOR2X1 U73490 ( .A(n43509), .B(n38558), .Y(n70492) );
  NAND2X1 U73491 ( .A(n43677), .B(n70479), .Y(n70481) );
  NAND2X1 U73492 ( .A(n70481), .B(n70480), .Y(n70482) );
  NAND2X1 U73493 ( .A(n36548), .B(n70482), .Y(n71111) );
  NOR2X1 U73494 ( .A(n39887), .B(n70483), .Y(n70485) );
  NAND2X1 U73495 ( .A(n40173), .B(n70504), .Y(n70484) );
  NAND2X1 U73496 ( .A(n70485), .B(n70484), .Y(n70488) );
  NOR2X1 U73497 ( .A(n70486), .B(n43688), .Y(n70487) );
  NAND2X1 U73498 ( .A(n39580), .B(n70487), .Y(n70491) );
  NOR2X1 U73499 ( .A(n43678), .B(n36560), .Y(n70489) );
  NAND2X1 U73500 ( .A(n70488), .B(n70489), .Y(n70490) );
  XNOR2X1 U73501 ( .A(n71137), .B(n43692), .Y(n70493) );
  XNOR2X1 U73502 ( .A(n70500), .B(n43708), .Y(n70494) );
  XNOR2X1 U73503 ( .A(n38080), .B(n70494), .Y(n70499) );
  XNOR2X1 U73504 ( .A(n70496), .B(n70495), .Y(n70497) );
  XNOR2X1 U73505 ( .A(n70497), .B(n42103), .Y(n70498) );
  MX2X1 U73506 ( .A(n70499), .B(n70498), .S0(n43719), .Y(u_muldiv_result_r[25]) );
  NAND2X1 U73507 ( .A(u_muldiv_mult_result_q[25]), .B(n44631), .Y(n13902) );
  NAND2X1 U73508 ( .A(n70500), .B(n43710), .Y(n70812) );
  NAND2X1 U73509 ( .A(n70501), .B(n36560), .Y(n70502) );
  NOR2X1 U73510 ( .A(n40173), .B(n70502), .Y(n70503) );
  NOR2X1 U73511 ( .A(n70503), .B(n71110), .Y(n70506) );
  NOR2X1 U73512 ( .A(n41307), .B(n41301), .Y(n70505) );
  NAND2X1 U73513 ( .A(n70505), .B(n70506), .Y(n70507) );
  NAND2X1 U73514 ( .A(n43677), .B(n38558), .Y(n71152) );
  INVX1 U73515 ( .A(n70508), .Y(n70510) );
  NAND2X1 U73516 ( .A(n70510), .B(n70509), .Y(n71166) );
  NAND2X1 U73517 ( .A(n70512), .B(n70511), .Y(n70514) );
  NAND2X1 U73518 ( .A(n70514), .B(n70513), .Y(n70830) );
  NAND2X1 U73519 ( .A(n71105), .B(n70831), .Y(n70515) );
  NOR2X1 U73520 ( .A(n39843), .B(n70515), .Y(n70765) );
  NOR2X1 U73521 ( .A(n38555), .B(n70517), .Y(n70518) );
  NOR2X1 U73522 ( .A(n70519), .B(n70518), .Y(n70520) );
  XNOR2X1 U73523 ( .A(n70526), .B(n70520), .Y(n70521) );
  INVX1 U73524 ( .A(n70523), .Y(n70522) );
  NAND2X1 U73525 ( .A(n43642), .B(n70522), .Y(n70824) );
  NAND2X1 U73526 ( .A(n70523), .B(n39301), .Y(n70525) );
  NAND2X1 U73527 ( .A(n70525), .B(n70524), .Y(n70825) );
  NAND2X1 U73528 ( .A(n70824), .B(n70825), .Y(n71173) );
  NAND2X1 U73529 ( .A(n70527), .B(n43668), .Y(n70529) );
  NAND2X1 U73530 ( .A(n70529), .B(n70528), .Y(n70848) );
  NAND2X1 U73531 ( .A(n70849), .B(n70848), .Y(n70845) );
  XNOR2X1 U73532 ( .A(n70530), .B(n39811), .Y(n70531) );
  XNOR2X1 U73533 ( .A(n38898), .B(n70531), .Y(n70532) );
  INVX1 U73534 ( .A(n70532), .Y(n70533) );
  NAND2X1 U73535 ( .A(n70533), .B(n39186), .Y(n70535) );
  NAND2X1 U73536 ( .A(n43535), .B(n70536), .Y(n70550) );
  NAND2X1 U73537 ( .A(n70537), .B(n43539), .Y(n70538) );
  NAND2X1 U73538 ( .A(n70539), .B(n70538), .Y(n70551) );
  NAND2X1 U73539 ( .A(n70550), .B(n70551), .Y(n70888) );
  XNOR2X1 U73540 ( .A(n43541), .B(n43621), .Y(n70540) );
  XNOR2X1 U73541 ( .A(n43566), .B(n70540), .Y(n70541) );
  INVX1 U73542 ( .A(n70889), .Y(n70558) );
  XNOR2X1 U73543 ( .A(n70541), .B(n70558), .Y(n70542) );
  XNOR2X1 U73544 ( .A(n39811), .B(n70543), .Y(n70545) );
  INVX1 U73545 ( .A(n70545), .Y(n70544) );
  NAND2X1 U73546 ( .A(n70545), .B(n43549), .Y(n70547) );
  XNOR2X1 U73547 ( .A(n70856), .B(n43633), .Y(n70761) );
  NAND2X1 U73548 ( .A(n70549), .B(n70548), .Y(n70756) );
  NAND2X1 U73549 ( .A(n70551), .B(n70550), .Y(n70552) );
  XOR2X1 U73550 ( .A(n70752), .B(n70552), .Y(n70553) );
  XOR2X1 U73551 ( .A(n70889), .B(n70553), .Y(n70554) );
  NAND2X1 U73552 ( .A(n70556), .B(n70555), .Y(n70868) );
  NAND2X1 U73553 ( .A(n43619), .B(n70557), .Y(n70867) );
  NAND2X1 U73554 ( .A(n70867), .B(n70868), .Y(n70861) );
  INVX1 U73555 ( .A(n70861), .Y(n71187) );
  NAND2X1 U73556 ( .A(n43535), .B(n70889), .Y(n70893) );
  NAND2X1 U73557 ( .A(n70559), .B(n70888), .Y(n70892) );
  NAND2X1 U73558 ( .A(n70893), .B(n70892), .Y(n70857) );
  INVX1 U73559 ( .A(n70560), .Y(n72078) );
  XNOR2X1 U73560 ( .A(n70897), .B(n72078), .Y(n70754) );
  NAND2X1 U73561 ( .A(n36604), .B(n70561), .Y(n70563) );
  NAND2X1 U73562 ( .A(n70563), .B(n70562), .Y(n70576) );
  NAND2X1 U73563 ( .A(n43577), .B(n70564), .Y(n70903) );
  INVX1 U73564 ( .A(n70564), .Y(n70565) );
  NAND2X1 U73565 ( .A(n70903), .B(n70900), .Y(n70881) );
  NAND2X1 U73566 ( .A(n70568), .B(n70567), .Y(n70570) );
  XNOR2X1 U73567 ( .A(n70733), .B(n70571), .Y(n70912) );
  INVX1 U73568 ( .A(n70743), .Y(n70573) );
  NAND2X1 U73569 ( .A(n43582), .B(n70574), .Y(n71088) );
  INVX1 U73570 ( .A(n70574), .Y(n70575) );
  NAND2X1 U73571 ( .A(n70575), .B(n43586), .Y(n70577) );
  NAND2X1 U73572 ( .A(n70577), .B(n70576), .Y(n71087) );
  INVX1 U73573 ( .A(n70912), .Y(n70746) );
  NAND2X1 U73574 ( .A(n43592), .B(n70746), .Y(n71078) );
  NAND2X1 U73575 ( .A(n43592), .B(n70578), .Y(n70581) );
  NAND2X1 U73576 ( .A(n38302), .B(n42994), .Y(n70579) );
  NAND2X1 U73577 ( .A(n41419), .B(n70579), .Y(n70580) );
  NAND2X1 U73578 ( .A(n43615), .B(n70582), .Y(n70586) );
  NAND2X1 U73579 ( .A(n70583), .B(n40683), .Y(n70584) );
  NAND2X1 U73580 ( .A(n70584), .B(n70728), .Y(n70585) );
  XNOR2X1 U73581 ( .A(n70589), .B(n39704), .Y(n70591) );
  INVX1 U73582 ( .A(n70591), .Y(n70590) );
  NAND2X1 U73583 ( .A(n43599), .B(n70590), .Y(n70595) );
  NAND2X1 U73584 ( .A(n70591), .B(n43597), .Y(n70593) );
  NAND2X1 U73585 ( .A(n70593), .B(n70592), .Y(n70594) );
  NAND2X1 U73586 ( .A(n70595), .B(n70594), .Y(n71055) );
  XNOR2X1 U73587 ( .A(n43618), .B(n41531), .Y(n70723) );
  NAND2X1 U73588 ( .A(n70597), .B(n70596), .Y(n70600) );
  NOR2X1 U73589 ( .A(n72219), .B(n70600), .Y(n70599) );
  INVX1 U73590 ( .A(n72219), .Y(n72217) );
  NAND2X1 U73591 ( .A(n72217), .B(n70598), .Y(n70971) );
  NAND2X1 U73592 ( .A(n70599), .B(n70971), .Y(n70604) );
  INVX1 U73593 ( .A(n70600), .Y(n70972) );
  NOR2X1 U73594 ( .A(n72217), .B(n70972), .Y(n70602) );
  NAND2X1 U73595 ( .A(n70601), .B(n72219), .Y(n70973) );
  NAND2X1 U73596 ( .A(n70602), .B(n70973), .Y(n70603) );
  XNOR2X1 U73597 ( .A(n72200), .B(n72212), .Y(n70675) );
  NAND2X1 U73598 ( .A(n70606), .B(n70605), .Y(n70614) );
  INVX1 U73599 ( .A(n70660), .Y(n70662) );
  NAND2X1 U73600 ( .A(n70608), .B(n70607), .Y(n70661) );
  INVX1 U73601 ( .A(n70609), .Y(n70665) );
  XNOR2X1 U73602 ( .A(n70661), .B(n70665), .Y(n70610) );
  NAND2X1 U73603 ( .A(n70611), .B(n44047), .Y(n70959) );
  INVX1 U73604 ( .A(n70959), .Y(n70612) );
  NAND2X1 U73605 ( .A(n70612), .B(n43493), .Y(n70615) );
  NAND2X1 U73606 ( .A(n70614), .B(n70613), .Y(n70954) );
  NAND2X1 U73607 ( .A(n70615), .B(n70954), .Y(n70979) );
  NAND2X1 U73608 ( .A(n70617), .B(n70616), .Y(n70620) );
  OR2X1 U73609 ( .A(n70617), .B(n70616), .Y(n70618) );
  NAND2X1 U73610 ( .A(n41733), .B(n70618), .Y(n70619) );
  NAND2X1 U73611 ( .A(n70620), .B(n70619), .Y(n70965) );
  INVX1 U73612 ( .A(n70965), .Y(n71341) );
  XNOR2X1 U73613 ( .A(n70979), .B(n71341), .Y(n70674) );
  NAND2X1 U73614 ( .A(n43491), .B(n44055), .Y(n70958) );
  NAND2X1 U73615 ( .A(n71013), .B(n71014), .Y(n71012) );
  OR2X1 U73616 ( .A(n71013), .B(n71014), .Y(n70621) );
  NAND2X1 U73617 ( .A(n42061), .B(n70621), .Y(n70622) );
  NAND2X1 U73618 ( .A(n71012), .B(n70622), .Y(n71010) );
  XNOR2X1 U73619 ( .A(n71010), .B(n41530), .Y(n70644) );
  NAND2X1 U73620 ( .A(n72355), .B(n71882), .Y(n70625) );
  NAND2X1 U73621 ( .A(n72355), .B(n70623), .Y(n70624) );
  NAND2X1 U73622 ( .A(n70625), .B(n70624), .Y(n71889) );
  XNOR2X1 U73623 ( .A(n70995), .B(n41701), .Y(n71308) );
  INVX1 U73624 ( .A(n71308), .Y(n70998) );
  NAND2X1 U73625 ( .A(n70626), .B(n43603), .Y(n72428) );
  INVX1 U73626 ( .A(n72428), .Y(n72425) );
  XNOR2X1 U73627 ( .A(n42056), .B(n72425), .Y(n70630) );
  NAND2X1 U73628 ( .A(n70628), .B(n70627), .Y(n70629) );
  NAND2X1 U73629 ( .A(n72263), .B(n70629), .Y(n70993) );
  INVX1 U73630 ( .A(n70993), .Y(n71000) );
  XNOR2X1 U73631 ( .A(n70630), .B(n71000), .Y(n70631) );
  XNOR2X1 U73632 ( .A(n41702), .B(n70631), .Y(n70636) );
  XNOR2X1 U73633 ( .A(n41697), .B(n70632), .Y(n70637) );
  INVX1 U73634 ( .A(n70637), .Y(n70633) );
  NAND2X1 U73635 ( .A(n72422), .B(n70633), .Y(n70635) );
  NAND2X1 U73636 ( .A(n72422), .B(n70638), .Y(n70634) );
  NAND2X1 U73637 ( .A(n70635), .B(n70634), .Y(n71001) );
  INVX1 U73638 ( .A(n71001), .Y(n71007) );
  XNOR2X1 U73639 ( .A(n70636), .B(n71007), .Y(n70643) );
  NAND2X1 U73640 ( .A(n70637), .B(n72356), .Y(n70639) );
  NOR2X1 U73641 ( .A(n70639), .B(n70638), .Y(n70641) );
  NOR2X1 U73642 ( .A(n70641), .B(n70640), .Y(n70642) );
  XNOR2X1 U73643 ( .A(n70643), .B(n70642), .Y(n71020) );
  INVX1 U73644 ( .A(n71020), .Y(n71011) );
  XNOR2X1 U73645 ( .A(n70644), .B(n71011), .Y(n70990) );
  INVX1 U73646 ( .A(n70991), .Y(n70645) );
  NAND2X1 U73647 ( .A(n70645), .B(n44016), .Y(n70649) );
  INVX1 U73648 ( .A(n70651), .Y(n70647) );
  NAND2X1 U73649 ( .A(n70647), .B(n70646), .Y(n70648) );
  NAND2X1 U73650 ( .A(n70648), .B(n43500), .Y(n70985) );
  NOR2X1 U73651 ( .A(n70649), .B(n70985), .Y(n70659) );
  NAND2X1 U73652 ( .A(n70985), .B(n70991), .Y(n70657) );
  NAND2X1 U73653 ( .A(n70651), .B(n70650), .Y(n70987) );
  INVX1 U73654 ( .A(n70987), .Y(n70652) );
  NAND2X1 U73655 ( .A(n70652), .B(n70991), .Y(n70655) );
  NAND2X1 U73656 ( .A(n44020), .B(n70991), .Y(n70653) );
  NAND2X1 U73657 ( .A(n70653), .B(n70987), .Y(n70654) );
  NAND2X1 U73658 ( .A(n70655), .B(n70654), .Y(n70656) );
  NAND2X1 U73659 ( .A(n70657), .B(n70656), .Y(n70658) );
  NAND2X1 U73660 ( .A(n70660), .B(n70661), .Y(n70667) );
  INVX1 U73661 ( .A(n70661), .Y(n70663) );
  NAND2X1 U73662 ( .A(n70663), .B(n70662), .Y(n70664) );
  NAND2X1 U73663 ( .A(n70665), .B(n70664), .Y(n70666) );
  NAND2X1 U73664 ( .A(n70667), .B(n70666), .Y(n71027) );
  INVX1 U73665 ( .A(n71027), .Y(n70668) );
  XNOR2X1 U73666 ( .A(n71028), .B(n70668), .Y(n70670) );
  NOR2X1 U73667 ( .A(n44052), .B(n43499), .Y(n70669) );
  XNOR2X1 U73668 ( .A(n70670), .B(n70669), .Y(n70952) );
  NAND2X1 U73669 ( .A(n43614), .B(n38310), .Y(n72225) );
  INVX1 U73670 ( .A(n72225), .Y(n72318) );
  XNOR2X1 U73671 ( .A(n70952), .B(n72318), .Y(n70672) );
  XNOR2X1 U73672 ( .A(n70958), .B(n70672), .Y(n70673) );
  XNOR2X1 U73673 ( .A(n70674), .B(n70673), .Y(n70969) );
  INVX1 U73674 ( .A(n70969), .Y(n70970) );
  XNOR2X1 U73675 ( .A(n70675), .B(n70970), .Y(n70676) );
  XNOR2X1 U73676 ( .A(n41673), .B(n70676), .Y(n70689) );
  NAND2X1 U73677 ( .A(n70677), .B(n72208), .Y(n70687) );
  NAND2X1 U73678 ( .A(n72212), .B(n70678), .Y(n70685) );
  NAND2X1 U73679 ( .A(n72212), .B(n70679), .Y(n70680) );
  NAND2X1 U73680 ( .A(n70681), .B(n70680), .Y(n70683) );
  NAND2X1 U73681 ( .A(n70683), .B(n70682), .Y(n70684) );
  NAND2X1 U73682 ( .A(n70685), .B(n70684), .Y(n70686) );
  NAND2X1 U73683 ( .A(n70687), .B(n70686), .Y(n70948) );
  INVX1 U73684 ( .A(n70948), .Y(n70688) );
  XNOR2X1 U73685 ( .A(n70689), .B(n70688), .Y(n70698) );
  NOR2X1 U73686 ( .A(n72200), .B(n41468), .Y(n70690) );
  NOR2X1 U73687 ( .A(n70691), .B(n70690), .Y(n70693) );
  NOR2X1 U73688 ( .A(n72200), .B(n70696), .Y(n70695) );
  INVX1 U73689 ( .A(n70704), .Y(n70931) );
  INVX1 U73690 ( .A(n70696), .Y(n70697) );
  INVX1 U73691 ( .A(n70935), .Y(n70930) );
  NAND2X1 U73692 ( .A(n70931), .B(n72196), .Y(n70699) );
  NOR2X1 U73693 ( .A(n70933), .B(n70699), .Y(n70702) );
  NAND2X1 U73694 ( .A(n70933), .B(n72510), .Y(n70700) );
  NOR2X1 U73695 ( .A(n41668), .B(n70700), .Y(n70701) );
  NOR2X1 U73696 ( .A(n70702), .B(n70701), .Y(n70703) );
  XNOR2X1 U73697 ( .A(n70930), .B(n70703), .Y(n70926) );
  INVX1 U73698 ( .A(n70926), .Y(n71259) );
  NAND2X1 U73699 ( .A(n70704), .B(n43001), .Y(n70707) );
  NAND2X1 U73700 ( .A(n70706), .B(n70705), .Y(n70717) );
  NAND2X1 U73701 ( .A(n70707), .B(n70717), .Y(n70923) );
  NAND2X1 U73702 ( .A(n70923), .B(n43000), .Y(n70711) );
  NOR2X1 U73703 ( .A(n71259), .B(n70711), .Y(n70710) );
  NAND2X1 U73704 ( .A(n72515), .B(n70717), .Y(n70708) );
  NAND2X1 U73705 ( .A(n72515), .B(n70931), .Y(n70924) );
  NOR2X1 U73706 ( .A(n71259), .B(n41461), .Y(n70709) );
  NOR2X1 U73707 ( .A(n70710), .B(n70709), .Y(n70715) );
  INVX1 U73708 ( .A(n70711), .Y(n70712) );
  NOR2X1 U73709 ( .A(n70712), .B(n70926), .Y(n70713) );
  NAND2X1 U73710 ( .A(n70713), .B(n41461), .Y(n70714) );
  NAND2X1 U73711 ( .A(n70715), .B(n70714), .Y(n71048) );
  NAND2X1 U73712 ( .A(n39704), .B(n39556), .Y(n70718) );
  NOR2X1 U73713 ( .A(n39126), .B(n71043), .Y(n70721) );
  INVX1 U73714 ( .A(n70719), .Y(n71042) );
  NAND2X1 U73715 ( .A(n39556), .B(n70719), .Y(n71045) );
  NOR2X1 U73716 ( .A(n70721), .B(n70720), .Y(n70722) );
  XNOR2X1 U73717 ( .A(n39066), .B(n70722), .Y(n71060) );
  INVX1 U73718 ( .A(n71060), .Y(n71056) );
  XNOR2X1 U73719 ( .A(n70723), .B(n71056), .Y(n70724) );
  XNOR2X1 U73720 ( .A(n71055), .B(n70724), .Y(n70725) );
  XNOR2X1 U73721 ( .A(n70726), .B(n43593), .Y(n70727) );
  XNOR2X1 U73722 ( .A(n41453), .B(n70727), .Y(n70740) );
  XNOR2X1 U73723 ( .A(n43616), .B(n70729), .Y(n70730) );
  XNOR2X1 U73724 ( .A(n70730), .B(n38938), .Y(n70731) );
  INVX1 U73725 ( .A(n70734), .Y(n70732) );
  NOR2X1 U73726 ( .A(n70732), .B(n42996), .Y(n70739) );
  NAND2X1 U73727 ( .A(n70734), .B(n70733), .Y(n70737) );
  OR2X1 U73728 ( .A(n70735), .B(n42997), .Y(n70736) );
  NAND2X1 U73729 ( .A(n70737), .B(n70736), .Y(n70738) );
  NOR2X1 U73730 ( .A(n70739), .B(n70738), .Y(n71072) );
  XNOR2X1 U73731 ( .A(n70740), .B(n71072), .Y(n70741) );
  XNOR2X1 U73732 ( .A(n41451), .B(n70741), .Y(n70750) );
  NOR2X1 U73733 ( .A(n43568), .B(n70912), .Y(n70742) );
  NAND2X1 U73734 ( .A(n38127), .B(n70742), .Y(n70749) );
  NAND2X1 U73735 ( .A(n70744), .B(n70743), .Y(n70745) );
  NOR2X1 U73736 ( .A(n40670), .B(n70745), .Y(n70747) );
  NAND2X1 U73737 ( .A(n43567), .B(n70746), .Y(n70915) );
  NAND2X1 U73738 ( .A(n70747), .B(n70915), .Y(n70748) );
  XNOR2X1 U73739 ( .A(n70750), .B(n41656), .Y(n70751) );
  XNOR2X1 U73740 ( .A(n41129), .B(n70751), .Y(n71218) );
  XNOR2X1 U73741 ( .A(n70752), .B(n71218), .Y(n70753) );
  XOR2X1 U73742 ( .A(n70881), .B(n70753), .Y(n70858) );
  XNOR2X1 U73743 ( .A(n70754), .B(n70858), .Y(n70760) );
  NAND2X1 U73744 ( .A(n70758), .B(n39629), .Y(n70757) );
  NAND2X1 U73745 ( .A(n70757), .B(n70756), .Y(n70869) );
  INVX1 U73746 ( .A(n70758), .Y(n70759) );
  NAND2X1 U73747 ( .A(n70759), .B(n43563), .Y(n70870) );
  NAND2X1 U73748 ( .A(n70869), .B(n70870), .Y(n70860) );
  INVX1 U73749 ( .A(n70860), .Y(n70885) );
  XNOR2X1 U73750 ( .A(n70761), .B(n40976), .Y(n70850) );
  XNOR2X1 U73751 ( .A(n70762), .B(n70850), .Y(n70763) );
  XNOR2X1 U73752 ( .A(n72586), .B(n70823), .Y(n70764) );
  INVX1 U73753 ( .A(n70766), .Y(n70768) );
  NOR2X1 U73754 ( .A(n39326), .B(n70769), .Y(n70779) );
  NOR2X1 U73755 ( .A(n43656), .B(n70771), .Y(n70772) );
  NOR2X1 U73756 ( .A(n70773), .B(n70772), .Y(n70774) );
  XNOR2X1 U73757 ( .A(n70775), .B(n70774), .Y(n70777) );
  XNOR2X1 U73758 ( .A(n70777), .B(n40956), .Y(n70778) );
  XNOR2X1 U73759 ( .A(n40162), .B(n70778), .Y(n70780) );
  XNOR2X1 U73760 ( .A(n41020), .B(n41028), .Y(n70787) );
  XNOR2X1 U73761 ( .A(n71109), .B(n41281), .Y(n70789) );
  NAND2X1 U73762 ( .A(n70789), .B(n43514), .Y(n70781) );
  OR2X1 U73763 ( .A(n38538), .B(n70781), .Y(n70782) );
  NOR2X1 U73764 ( .A(n71145), .B(n70782), .Y(n70815) );
  NAND2X1 U73765 ( .A(n38538), .B(n70784), .Y(n70786) );
  NOR2X1 U73766 ( .A(n70789), .B(n70786), .Y(n70788) );
  NOR2X1 U73767 ( .A(n70815), .B(n39925), .Y(n70793) );
  XNOR2X1 U73768 ( .A(n41020), .B(n41028), .Y(n71145) );
  NOR2X1 U73769 ( .A(n36564), .B(n70788), .Y(n70792) );
  NAND2X1 U73770 ( .A(n70792), .B(n70791), .Y(n70816) );
  INVX1 U73771 ( .A(n71137), .Y(n70794) );
  NAND2X1 U73772 ( .A(n41454), .B(n70794), .Y(n70819) );
  XNOR2X1 U73773 ( .A(n71416), .B(n70795), .Y(n70803) );
  XNOR2X1 U73774 ( .A(n43715), .B(n70803), .Y(n70796) );
  XNOR2X1 U73775 ( .A(n70797), .B(n70796), .Y(n70802) );
  XNOR2X1 U73776 ( .A(n70799), .B(n70798), .Y(n70800) );
  XOR2X1 U73777 ( .A(n42109), .B(n70800), .Y(n70801) );
  MX2X1 U73778 ( .A(n70802), .B(n70801), .S0(n43718), .Y(u_muldiv_result_r[26]) );
  NAND2X1 U73779 ( .A(u_muldiv_mult_result_q[26]), .B(n44631), .Y(n13894) );
  NOR2X1 U73780 ( .A(n70803), .B(n43714), .Y(n70804) );
  NOR2X1 U73781 ( .A(n40020), .B(n70806), .Y(n70807) );
  NOR2X1 U73782 ( .A(n38069), .B(n70807), .Y(n70811) );
  NOR2X1 U73783 ( .A(n41197), .B(n36436), .Y(n70808) );
  NAND2X1 U73784 ( .A(n70808), .B(n40982), .Y(n70809) );
  NAND2X1 U73785 ( .A(n43705), .B(n70809), .Y(n70810) );
  NAND2X1 U73786 ( .A(n70811), .B(n70810), .Y(n70813) );
  NAND2X1 U73787 ( .A(n71125), .B(n38887), .Y(n71120) );
  NAND2X1 U73788 ( .A(n70793), .B(n70816), .Y(n70817) );
  NAND2X1 U73789 ( .A(n70787), .B(n43512), .Y(n71704) );
  NAND2X1 U73790 ( .A(n70821), .B(n70820), .Y(n71144) );
  NAND2X1 U73791 ( .A(n71144), .B(n70822), .Y(n71703) );
  NAND2X1 U73792 ( .A(n70824), .B(n70825), .Y(n70826) );
  XNOR2X1 U73793 ( .A(n70827), .B(n43654), .Y(n70828) );
  XNOR2X1 U73794 ( .A(n40956), .B(n70828), .Y(n70834) );
  NAND2X1 U73795 ( .A(n70829), .B(n43657), .Y(n70832) );
  NAND2X1 U73796 ( .A(n43653), .B(n70830), .Y(n70831) );
  NAND2X1 U73797 ( .A(n70831), .B(n70832), .Y(n70833) );
  NOR2X1 U73798 ( .A(n70834), .B(n70833), .Y(n70835) );
  NOR2X1 U73799 ( .A(n40562), .B(n71157), .Y(n70842) );
  NOR2X1 U73800 ( .A(n70839), .B(n70838), .Y(n70841) );
  NAND2X1 U73801 ( .A(n70841), .B(n70840), .Y(n71158) );
  NOR2X1 U73802 ( .A(n71157), .B(n43532), .Y(n70843) );
  XNOR2X1 U73803 ( .A(n43673), .B(n70851), .Y(n70844) );
  NAND2X1 U73804 ( .A(n71174), .B(n70847), .Y(n71176) );
  INVX1 U73805 ( .A(n70850), .Y(n70853) );
  XNOR2X1 U73806 ( .A(n70851), .B(n70853), .Y(n70852) );
  NAND2X1 U73807 ( .A(n70853), .B(n38555), .Y(n71170) );
  INVX1 U73808 ( .A(n39043), .Y(n70866) );
  XNOR2X1 U73809 ( .A(n70866), .B(n40976), .Y(n70854) );
  INVX1 U73810 ( .A(n70854), .Y(n70855) );
  NAND2X1 U73811 ( .A(n70855), .B(n39186), .Y(n71180) );
  NAND2X1 U73812 ( .A(n38692), .B(n71180), .Y(n71101) );
  NOR2X1 U73813 ( .A(n43546), .B(n39043), .Y(n70864) );
  INVX1 U73814 ( .A(n70857), .Y(n71217) );
  XNOR2X1 U73815 ( .A(n43628), .B(n70872), .Y(n70859) );
  INVX1 U73816 ( .A(n70865), .Y(n70862) );
  NOR2X1 U73817 ( .A(n43546), .B(n70862), .Y(n70863) );
  NAND2X1 U73818 ( .A(n70868), .B(n70867), .Y(n70874) );
  NAND2X1 U73819 ( .A(n70870), .B(n70869), .Y(n70871) );
  XNOR2X1 U73820 ( .A(n70872), .B(n70871), .Y(n70875) );
  NAND2X1 U73821 ( .A(n43619), .B(n70875), .Y(n71186) );
  NAND2X1 U73822 ( .A(n71810), .B(n71186), .Y(n70873) );
  NOR2X1 U73823 ( .A(n70874), .B(n70873), .Y(n70878) );
  INVX1 U73824 ( .A(n70875), .Y(n70876) );
  NAND2X1 U73825 ( .A(n70876), .B(n43623), .Y(n71188) );
  NOR2X1 U73826 ( .A(n72587), .B(n71188), .Y(n70877) );
  NOR2X1 U73827 ( .A(n70878), .B(n70877), .Y(n70880) );
  NAND2X1 U73828 ( .A(n71189), .B(n72587), .Y(n70879) );
  NAND2X1 U73829 ( .A(n70880), .B(n70879), .Y(n71098) );
  INVX1 U73830 ( .A(n70881), .Y(n71230) );
  XNOR2X1 U73831 ( .A(n71218), .B(n43537), .Y(n70882) );
  XNOR2X1 U73832 ( .A(n71230), .B(n70882), .Y(n70886) );
  XNOR2X1 U73833 ( .A(n70886), .B(n71217), .Y(n70883) );
  NAND2X1 U73834 ( .A(n43562), .B(n70883), .Y(n70884) );
  INVX1 U73835 ( .A(n70886), .Y(n70887) );
  XNOR2X1 U73836 ( .A(n71212), .B(n43621), .Y(n71097) );
  INVX1 U73837 ( .A(n71218), .Y(n70894) );
  NAND2X1 U73838 ( .A(n70894), .B(n43539), .Y(n70891) );
  NAND2X1 U73839 ( .A(n70889), .B(n70888), .Y(n70890) );
  NOR2X1 U73840 ( .A(n70891), .B(n70890), .Y(n70899) );
  NAND2X1 U73841 ( .A(n70893), .B(n70892), .Y(n70897) );
  XNOR2X1 U73842 ( .A(n70894), .B(n71230), .Y(n71215) );
  INVX1 U73843 ( .A(n71215), .Y(n70895) );
  NAND2X1 U73844 ( .A(n43535), .B(n70895), .Y(n70896) );
  NOR2X1 U73845 ( .A(n70897), .B(n70896), .Y(n70898) );
  NOR2X1 U73846 ( .A(n70899), .B(n70898), .Y(n71096) );
  INVX1 U73847 ( .A(n70900), .Y(n70905) );
  NAND2X1 U73848 ( .A(n43576), .B(n38889), .Y(n70902) );
  NOR2X1 U73849 ( .A(n39869), .B(n70902), .Y(n70904) );
  NOR2X1 U73850 ( .A(n70905), .B(n41462), .Y(n70910) );
  XNOR2X1 U73851 ( .A(n71072), .B(n41453), .Y(n71075) );
  INVX1 U73852 ( .A(n71075), .Y(n71077) );
  XNOR2X1 U73853 ( .A(n42993), .B(n43582), .Y(n70906) );
  XNOR2X1 U73854 ( .A(n71077), .B(n70906), .Y(n70907) );
  XNOR2X1 U73855 ( .A(n70907), .B(n41451), .Y(n70908) );
  XNOR2X1 U73856 ( .A(n41129), .B(n70908), .Y(n71227) );
  NOR2X1 U73857 ( .A(n41462), .B(n71227), .Y(n70909) );
  NOR2X1 U73858 ( .A(n70910), .B(n70909), .Y(n70911) );
  NAND2X1 U73859 ( .A(n43576), .B(n71227), .Y(n71229) );
  NAND2X1 U73860 ( .A(n70911), .B(n71229), .Y(n71211) );
  NAND2X1 U73861 ( .A(n70912), .B(n40670), .Y(n70914) );
  NAND2X1 U73862 ( .A(n70914), .B(n70913), .Y(n70916) );
  NAND2X1 U73863 ( .A(n70916), .B(n70915), .Y(n70920) );
  NOR2X1 U73864 ( .A(n43568), .B(n70920), .Y(n70919) );
  XNOR2X1 U73865 ( .A(n71075), .B(n43593), .Y(n70917) );
  XNOR2X1 U73866 ( .A(n41451), .B(n70917), .Y(n70921) );
  INVX1 U73867 ( .A(n70921), .Y(n71086) );
  NOR2X1 U73868 ( .A(n43568), .B(n71086), .Y(n70918) );
  INVX1 U73869 ( .A(n70920), .Y(n70922) );
  NAND2X1 U73870 ( .A(n70924), .B(n70923), .Y(n70927) );
  INVX1 U73871 ( .A(n70927), .Y(n71261) );
  NAND2X1 U73872 ( .A(n71261), .B(n70926), .Y(n70925) );
  NOR2X1 U73873 ( .A(n43001), .B(n70925), .Y(n70929) );
  NAND2X1 U73874 ( .A(n70926), .B(n43000), .Y(n71262) );
  NOR2X1 U73875 ( .A(n70929), .B(n70928), .Y(n71041) );
  NAND2X1 U73876 ( .A(n70930), .B(n72196), .Y(n70939) );
  NOR2X1 U73877 ( .A(n72510), .B(n70931), .Y(n70932) );
  NOR2X1 U73878 ( .A(n70933), .B(n70932), .Y(n70934) );
  NOR2X1 U73879 ( .A(n41668), .B(n70934), .Y(n70937) );
  NAND2X1 U73880 ( .A(n72510), .B(n70935), .Y(n70936) );
  NAND2X1 U73881 ( .A(n70937), .B(n70936), .Y(n70938) );
  NAND2X1 U73882 ( .A(n70939), .B(n70938), .Y(n71273) );
  INVX1 U73883 ( .A(n71273), .Y(n70945) );
  XNOR2X1 U73884 ( .A(n41673), .B(n70970), .Y(n70947) );
  INVX1 U73885 ( .A(n70947), .Y(n70946) );
  NAND2X1 U73886 ( .A(n70946), .B(n72202), .Y(n70943) );
  NAND2X1 U73887 ( .A(n72200), .B(n70947), .Y(n70941) );
  NAND2X1 U73888 ( .A(n70941), .B(n70940), .Y(n70942) );
  NAND2X1 U73889 ( .A(n70943), .B(n70942), .Y(n71280) );
  XNOR2X1 U73890 ( .A(n71280), .B(n72510), .Y(n70944) );
  XNOR2X1 U73891 ( .A(n70945), .B(n70944), .Y(n71039) );
  NAND2X1 U73892 ( .A(n70946), .B(n72208), .Y(n70951) );
  NAND2X1 U73893 ( .A(n72212), .B(n70947), .Y(n70949) );
  NAND2X1 U73894 ( .A(n70949), .B(n70948), .Y(n70950) );
  NAND2X1 U73895 ( .A(n70951), .B(n70950), .Y(n71359) );
  NOR2X1 U73896 ( .A(n71341), .B(n72318), .Y(n70963) );
  INVX1 U73897 ( .A(n70952), .Y(n70980) );
  INVX1 U73898 ( .A(n70954), .Y(n70953) );
  NOR2X1 U73899 ( .A(n70953), .B(n70958), .Y(n70957) );
  INVX1 U73900 ( .A(n70958), .Y(n70955) );
  NOR2X1 U73901 ( .A(n70955), .B(n70954), .Y(n70956) );
  NOR2X1 U73902 ( .A(n70957), .B(n70956), .Y(n70961) );
  NOR2X1 U73903 ( .A(n70959), .B(n70958), .Y(n70960) );
  NOR2X1 U73904 ( .A(n70961), .B(n70960), .Y(n70962) );
  XNOR2X1 U73905 ( .A(n70980), .B(n70962), .Y(n70964) );
  NAND2X1 U73906 ( .A(n70964), .B(n72225), .Y(n71342) );
  NAND2X1 U73907 ( .A(n70963), .B(n71342), .Y(n70968) );
  INVX1 U73908 ( .A(n70964), .Y(n71339) );
  NOR2X1 U73909 ( .A(n71339), .B(n70965), .Y(n70966) );
  NAND2X1 U73910 ( .A(n72318), .B(n70966), .Y(n70967) );
  NAND2X1 U73911 ( .A(n70968), .B(n70967), .Y(n71350) );
  NAND2X1 U73912 ( .A(n70969), .B(n72219), .Y(n70978) );
  NAND2X1 U73913 ( .A(n72217), .B(n70970), .Y(n70976) );
  NAND2X1 U73914 ( .A(n70972), .B(n70971), .Y(n70974) );
  NAND2X1 U73915 ( .A(n70974), .B(n70973), .Y(n70975) );
  NAND2X1 U73916 ( .A(n70976), .B(n70975), .Y(n70977) );
  NAND2X1 U73917 ( .A(n70978), .B(n70977), .Y(n71352) );
  XNOR2X1 U73918 ( .A(n71350), .B(n71352), .Y(n71038) );
  NAND2X1 U73919 ( .A(n70980), .B(n70979), .Y(n70984) );
  NOR2X1 U73920 ( .A(n70980), .B(n70979), .Y(n70981) );
  NOR2X1 U73921 ( .A(n44060), .B(n70981), .Y(n70982) );
  NAND2X1 U73922 ( .A(n70982), .B(n43493), .Y(n70983) );
  INVX1 U73923 ( .A(n70985), .Y(n70986) );
  NAND2X1 U73924 ( .A(n70986), .B(n44016), .Y(n70988) );
  NAND2X1 U73925 ( .A(n70988), .B(n70987), .Y(n70989) );
  NAND2X1 U73926 ( .A(n70990), .B(n70989), .Y(n71328) );
  NOR2X1 U73927 ( .A(n70990), .B(n70989), .Y(n70992) );
  OR2X1 U73928 ( .A(n70992), .B(n70991), .Y(n71331) );
  NAND2X1 U73929 ( .A(n71328), .B(n71331), .Y(n71327) );
  NAND2X1 U73930 ( .A(n44016), .B(n43607), .Y(n71299) );
  NAND2X1 U73931 ( .A(n42056), .B(n43603), .Y(n72434) );
  NAND2X1 U73932 ( .A(n70998), .B(n70993), .Y(n70994) );
  NAND2X1 U73933 ( .A(n72422), .B(n70994), .Y(n71305) );
  NAND2X1 U73934 ( .A(n72263), .B(n71889), .Y(n70997) );
  NAND2X1 U73935 ( .A(n72263), .B(n70995), .Y(n70996) );
  NAND2X1 U73936 ( .A(n70997), .B(n70996), .Y(n71886) );
  XNOR2X1 U73937 ( .A(n70998), .B(n41700), .Y(n71307) );
  XNOR2X1 U73938 ( .A(n72428), .B(n71307), .Y(n70999) );
  XNOR2X1 U73939 ( .A(n72434), .B(n71314), .Y(n71004) );
  XNOR2X1 U73940 ( .A(n41702), .B(n71000), .Y(n71005) );
  NAND2X1 U73941 ( .A(n72425), .B(n71005), .Y(n71003) );
  NAND2X1 U73942 ( .A(n72425), .B(n71001), .Y(n71002) );
  NAND2X1 U73943 ( .A(n71003), .B(n71002), .Y(n71315) );
  NOR2X1 U73944 ( .A(n72425), .B(n71005), .Y(n71006) );
  NAND2X1 U73945 ( .A(n71007), .B(n71006), .Y(n71008) );
  AND2X1 U73946 ( .A(n42056), .B(n71008), .Y(n71301) );
  XNOR2X1 U73947 ( .A(n71009), .B(n71301), .Y(n71320) );
  NAND2X1 U73948 ( .A(n44024), .B(n39960), .Y(n71024) );
  NAND2X1 U73949 ( .A(n71011), .B(n71010), .Y(n71023) );
  INVX1 U73950 ( .A(n71012), .Y(n71018) );
  NAND2X1 U73951 ( .A(n71013), .B(n42061), .Y(n71016) );
  NAND2X1 U73952 ( .A(n42061), .B(n71014), .Y(n71015) );
  NAND2X1 U73953 ( .A(n71016), .B(n71015), .Y(n71017) );
  NOR2X1 U73954 ( .A(n71018), .B(n71017), .Y(n71019) );
  NAND2X1 U73955 ( .A(n71020), .B(n71019), .Y(n71021) );
  NAND2X1 U73956 ( .A(n41530), .B(n71021), .Y(n71022) );
  NAND2X1 U73957 ( .A(n71023), .B(n71022), .Y(n71319) );
  XNOR2X1 U73958 ( .A(n71024), .B(n71319), .Y(n71025) );
  XNOR2X1 U73959 ( .A(n71327), .B(n71329), .Y(n71026) );
  XNOR2X1 U73960 ( .A(n71026), .B(n41735), .Y(n71291) );
  INVX1 U73961 ( .A(n71291), .Y(n71292) );
  NAND2X1 U73962 ( .A(n71028), .B(n71027), .Y(n71032) );
  NOR2X1 U73963 ( .A(n71028), .B(n71027), .Y(n71029) );
  NOR2X1 U73964 ( .A(n44052), .B(n71029), .Y(n71030) );
  NAND2X1 U73965 ( .A(n71030), .B(n43496), .Y(n71031) );
  NAND2X1 U73966 ( .A(n71032), .B(n71031), .Y(n71290) );
  INVX1 U73967 ( .A(n71290), .Y(n71293) );
  XNOR2X1 U73968 ( .A(n71292), .B(n71293), .Y(n71035) );
  NAND2X1 U73969 ( .A(n43614), .B(n43493), .Y(n72233) );
  XNOR2X1 U73970 ( .A(n72233), .B(n41736), .Y(n71034) );
  XNOR2X1 U73971 ( .A(n71035), .B(n71034), .Y(n71036) );
  XNOR2X1 U73972 ( .A(n41679), .B(n71036), .Y(n71338) );
  XNOR2X1 U73973 ( .A(n72212), .B(n72217), .Y(n71348) );
  XNOR2X1 U73974 ( .A(n71338), .B(n71348), .Y(n71037) );
  XNOR2X1 U73975 ( .A(n71038), .B(n71037), .Y(n71277) );
  XNOR2X1 U73976 ( .A(n71039), .B(n71265), .Y(n71040) );
  XNOR2X1 U73977 ( .A(n71041), .B(n71040), .Y(n71250) );
  INVX1 U73978 ( .A(n71250), .Y(n71249) );
  NAND2X1 U73979 ( .A(n71042), .B(n42998), .Y(n71044) );
  NAND2X1 U73980 ( .A(n71044), .B(n71043), .Y(n71046) );
  NAND2X1 U73981 ( .A(n71046), .B(n71045), .Y(n71049) );
  INVX1 U73982 ( .A(n71049), .Y(n71252) );
  NAND2X1 U73983 ( .A(n71252), .B(n39556), .Y(n71047) );
  NOR2X1 U73984 ( .A(n39066), .B(n71047), .Y(n71053) );
  NAND2X1 U73985 ( .A(n71048), .B(n42998), .Y(n71253) );
  INVX1 U73986 ( .A(n71253), .Y(n71051) );
  NAND2X1 U73987 ( .A(n71049), .B(n42999), .Y(n71050) );
  NOR2X1 U73988 ( .A(n71051), .B(n71050), .Y(n71052) );
  NOR2X1 U73989 ( .A(n71053), .B(n71052), .Y(n71054) );
  XNOR2X1 U73990 ( .A(n71249), .B(n71054), .Y(n71246) );
  INVX1 U73991 ( .A(n71246), .Y(n71243) );
  XNOR2X1 U73992 ( .A(n43602), .B(n71243), .Y(n71068) );
  NAND2X1 U73993 ( .A(n71060), .B(n43597), .Y(n71059) );
  INVX1 U73994 ( .A(n71055), .Y(n71062) );
  NAND2X1 U73995 ( .A(n43599), .B(n71056), .Y(n71057) );
  NAND2X1 U73996 ( .A(n71062), .B(n71057), .Y(n71058) );
  NAND2X1 U73997 ( .A(n71059), .B(n71058), .Y(n71244) );
  INVX1 U73998 ( .A(n71244), .Y(n71234) );
  XNOR2X1 U73999 ( .A(n72358), .B(n71234), .Y(n71066) );
  XNOR2X1 U74000 ( .A(n71060), .B(n43602), .Y(n71061) );
  XNOR2X1 U74001 ( .A(n71062), .B(n71061), .Y(n71070) );
  INVX1 U74002 ( .A(n71070), .Y(n71069) );
  NAND2X1 U74003 ( .A(n71069), .B(n40683), .Y(n71065) );
  NAND2X1 U74004 ( .A(n43615), .B(n71070), .Y(n71063) );
  NAND2X1 U74005 ( .A(n41657), .B(n71063), .Y(n71064) );
  NAND2X1 U74006 ( .A(n71065), .B(n71064), .Y(n71368) );
  NAND2X1 U74007 ( .A(n71069), .B(n42995), .Y(n71074) );
  NAND2X1 U74008 ( .A(n43617), .B(n71070), .Y(n71071) );
  NAND2X1 U74009 ( .A(n71072), .B(n71071), .Y(n71073) );
  NAND2X1 U74010 ( .A(n71074), .B(n71073), .Y(n71235) );
  NAND2X1 U74011 ( .A(n43592), .B(n71075), .Y(n71373) );
  NOR2X1 U74012 ( .A(n71079), .B(n71076), .Y(n71084) );
  NAND2X1 U74013 ( .A(n71077), .B(n42993), .Y(n71374) );
  NAND2X1 U74014 ( .A(n71079), .B(n71078), .Y(n71082) );
  NAND2X1 U74015 ( .A(n71373), .B(n71080), .Y(n71081) );
  NOR2X1 U74016 ( .A(n71084), .B(n71083), .Y(n71085) );
  INVX1 U74017 ( .A(n71386), .Y(n71387) );
  NAND2X1 U74018 ( .A(n41656), .B(n71086), .Y(n71388) );
  NAND2X1 U74019 ( .A(n71088), .B(n71087), .Y(n71091) );
  NAND2X1 U74020 ( .A(n71091), .B(n43585), .Y(n71089) );
  NOR2X1 U74021 ( .A(n71388), .B(n71089), .Y(n71093) );
  NAND2X1 U74022 ( .A(n43581), .B(n71388), .Y(n71090) );
  NOR2X1 U74023 ( .A(n71091), .B(n71090), .Y(n71092) );
  NOR2X1 U74024 ( .A(n71093), .B(n71092), .Y(n71094) );
  XNOR2X1 U74025 ( .A(n43560), .B(n71226), .Y(n71095) );
  XNOR2X1 U74026 ( .A(n71097), .B(n71204), .Y(n71190) );
  INVX1 U74027 ( .A(n71190), .Y(n71198) );
  XNOR2X1 U74028 ( .A(n39728), .B(n71099), .Y(n71178) );
  XNOR2X1 U74029 ( .A(n43672), .B(n71178), .Y(n71100) );
  XNOR2X1 U74030 ( .A(n71101), .B(n71100), .Y(n71167) );
  XNOR2X1 U74031 ( .A(n71102), .B(n71167), .Y(n71103) );
  XNOR2X1 U74032 ( .A(n71161), .B(n43523), .Y(n71107) );
  NAND2X1 U74033 ( .A(n71104), .B(n43657), .Y(n71747) );
  INVX1 U74034 ( .A(n71169), .Y(n71162) );
  XNOR2X1 U74035 ( .A(n71107), .B(n71162), .Y(n71150) );
  XNOR2X1 U74036 ( .A(n43687), .B(n71150), .Y(n71108) );
  XOR2X1 U74037 ( .A(n38145), .B(n71108), .Y(n71149) );
  NOR2X1 U74038 ( .A(n43678), .B(n71109), .Y(n71110) );
  NAND2X1 U74039 ( .A(n36559), .B(n71111), .Y(n71112) );
  NOR2X1 U74040 ( .A(n39887), .B(n71112), .Y(n71113) );
  NAND2X1 U74041 ( .A(n43676), .B(n71116), .Y(n71154) );
  NAND2X1 U74042 ( .A(n71434), .B(n71435), .Y(n71430) );
  XNOR2X1 U74043 ( .A(n43694), .B(n43508), .Y(n71404) );
  XNOR2X1 U74044 ( .A(n71430), .B(n71404), .Y(n71117) );
  XOR2X1 U74045 ( .A(n71149), .B(n71117), .Y(n71118) );
  XNOR2X1 U74046 ( .A(n71126), .B(n43707), .Y(n71119) );
  XNOR2X1 U74047 ( .A(n71120), .B(n71119), .Y(n71124) );
  XNOR2X1 U74048 ( .A(n36350), .B(n71121), .Y(n71122) );
  XNOR2X1 U74049 ( .A(n71122), .B(n42115), .Y(n71123) );
  MX2X1 U74050 ( .A(n71124), .B(n71123), .S0(n43718), .Y(u_muldiv_result_r[27]) );
  NAND2X1 U74051 ( .A(u_muldiv_mult_result_q[27]), .B(n44631), .Y(n13883) );
  NAND2X1 U74052 ( .A(n72107), .B(n72715), .Y(n71407) );
  XNOR2X1 U74053 ( .A(n43508), .B(n71430), .Y(n71127) );
  XNOR2X1 U74054 ( .A(n71149), .B(n71127), .Y(n71143) );
  INVX1 U74055 ( .A(n71143), .Y(n71418) );
  INVX1 U74056 ( .A(n71128), .Y(n71136) );
  NAND2X1 U74057 ( .A(n71130), .B(n71129), .Y(n71134) );
  NAND2X1 U74058 ( .A(n71132), .B(n71131), .Y(n71133) );
  NOR2X1 U74059 ( .A(n71134), .B(n71133), .Y(n71135) );
  NOR2X1 U74060 ( .A(n71136), .B(n71135), .Y(n71139) );
  NOR2X1 U74061 ( .A(n71137), .B(n43702), .Y(n71138) );
  NOR2X1 U74062 ( .A(n71139), .B(n71138), .Y(n71140) );
  INVX1 U74063 ( .A(n71704), .Y(n71148) );
  NOR2X1 U74064 ( .A(n70787), .B(n43512), .Y(n71146) );
  NOR2X1 U74065 ( .A(n36573), .B(n71146), .Y(n71147) );
  NAND2X1 U74066 ( .A(n43507), .B(n71706), .Y(n71724) );
  NAND2X1 U74067 ( .A(n43676), .B(n38435), .Y(n71156) );
  INVX1 U74068 ( .A(n71157), .Y(n71159) );
  NOR2X1 U74069 ( .A(n71159), .B(n40320), .Y(n71160) );
  NOR2X1 U74070 ( .A(n71160), .B(n43528), .Y(n71164) );
  INVX1 U74071 ( .A(n71161), .Y(n71163) );
  NOR2X1 U74072 ( .A(n71164), .B(n40262), .Y(n71165) );
  NAND2X1 U74073 ( .A(n41035), .B(n40955), .Y(n71697) );
  NAND2X1 U74074 ( .A(n71166), .B(n43657), .Y(n71749) );
  NAND2X1 U74075 ( .A(n71749), .B(n71747), .Y(n71426) );
  XNOR2X1 U74076 ( .A(n43644), .B(n38931), .Y(n71168) );
  INVX1 U74077 ( .A(n71167), .Y(n71172) );
  NAND2X1 U74078 ( .A(n71748), .B(n71169), .Y(n71423) );
  NAND2X1 U74079 ( .A(n71748), .B(n43656), .Y(n71424) );
  OR2X1 U74080 ( .A(n71426), .B(n71425), .Y(n71698) );
  NAND2X1 U74081 ( .A(n71171), .B(n71170), .Y(n71182) );
  NAND2X1 U74082 ( .A(n71174), .B(n71173), .Y(n71175) );
  NAND2X1 U74083 ( .A(n71177), .B(n71176), .Y(n71688) );
  NAND2X1 U74084 ( .A(n71180), .B(n71179), .Y(n71195) );
  INVX1 U74085 ( .A(n71195), .Y(n71185) );
  NAND2X1 U74086 ( .A(n71181), .B(n38555), .Y(n71184) );
  NAND2X1 U74087 ( .A(n71187), .B(n71186), .Y(n71189) );
  NAND2X1 U74088 ( .A(n71189), .B(n71188), .Y(n71206) );
  XNOR2X1 U74089 ( .A(n71190), .B(n43546), .Y(n71191) );
  XNOR2X1 U74090 ( .A(n71206), .B(n71191), .Y(n71192) );
  XNOR2X1 U74091 ( .A(n39728), .B(n71192), .Y(n71196) );
  INVX1 U74092 ( .A(n71196), .Y(n71193) );
  NOR2X1 U74093 ( .A(n43632), .B(n71193), .Y(n71194) );
  NAND2X1 U74094 ( .A(n71196), .B(n71195), .Y(n71197) );
  INVX1 U74095 ( .A(n71439), .Y(n71449) );
  NAND2X1 U74096 ( .A(n71199), .B(n43549), .Y(n71203) );
  INVX1 U74097 ( .A(n71199), .Y(n71200) );
  NAND2X1 U74098 ( .A(n43544), .B(n71200), .Y(n71202) );
  NAND2X1 U74099 ( .A(n71202), .B(n71201), .Y(n71442) );
  NAND2X1 U74100 ( .A(n71203), .B(n71442), .Y(n71660) );
  INVX1 U74101 ( .A(n71208), .Y(n71205) );
  NAND2X1 U74102 ( .A(n43619), .B(n71205), .Y(n71207) );
  NAND2X1 U74103 ( .A(n71207), .B(n71206), .Y(n71210) );
  NAND2X1 U74104 ( .A(n71208), .B(n43623), .Y(n71209) );
  NAND2X1 U74105 ( .A(n71210), .B(n71209), .Y(n71668) );
  INVX1 U74106 ( .A(n71668), .Y(n71469) );
  NAND2X1 U74107 ( .A(n39581), .B(n43563), .Y(n71213) );
  INVX1 U74108 ( .A(n71662), .Y(n71799) );
  XNOR2X1 U74109 ( .A(n43633), .B(n72078), .Y(n71461) );
  INVX1 U74110 ( .A(n71461), .Y(n71459) );
  XNOR2X1 U74111 ( .A(n71799), .B(n71459), .Y(n71397) );
  NAND2X1 U74112 ( .A(n71214), .B(n43539), .Y(n71224) );
  NAND2X1 U74113 ( .A(n39581), .B(n43536), .Y(n71222) );
  NAND2X1 U74114 ( .A(n43535), .B(n71215), .Y(n71216) );
  NAND2X1 U74115 ( .A(n71217), .B(n71216), .Y(n71220) );
  NAND2X1 U74116 ( .A(n71218), .B(n43539), .Y(n71219) );
  NAND2X1 U74117 ( .A(n71220), .B(n71219), .Y(n71221) );
  NAND2X1 U74118 ( .A(n71222), .B(n71221), .Y(n71223) );
  NAND2X1 U74119 ( .A(n71224), .B(n71223), .Y(n71654) );
  INVX1 U74120 ( .A(n71226), .Y(n71225) );
  NAND2X1 U74121 ( .A(n71225), .B(n43573), .Y(n71645) );
  NAND2X1 U74122 ( .A(n43577), .B(n71226), .Y(n71232) );
  INVX1 U74123 ( .A(n71227), .Y(n71228) );
  NAND2X1 U74124 ( .A(n71228), .B(n43573), .Y(n71642) );
  NAND2X1 U74125 ( .A(n71230), .B(n71229), .Y(n71641) );
  NAND2X1 U74126 ( .A(n71642), .B(n71641), .Y(n71231) );
  NAND2X1 U74127 ( .A(n71232), .B(n71231), .Y(n71233) );
  NAND2X1 U74128 ( .A(n39236), .B(n42996), .Y(n71238) );
  NAND2X1 U74129 ( .A(n39788), .B(n43618), .Y(n71236) );
  NAND2X1 U74130 ( .A(n71236), .B(n71235), .Y(n71237) );
  XNOR2X1 U74131 ( .A(n72353), .B(n41670), .Y(n71630) );
  NAND2X1 U74132 ( .A(n71606), .B(n40670), .Y(n71242) );
  INVX1 U74133 ( .A(n71606), .Y(n71607) );
  NAND2X1 U74134 ( .A(n43567), .B(n71607), .Y(n71240) );
  NAND2X1 U74135 ( .A(n71240), .B(n71239), .Y(n71241) );
  XNOR2X1 U74136 ( .A(n71630), .B(n41800), .Y(n71385) );
  NAND2X1 U74137 ( .A(n43602), .B(n71243), .Y(n71245) );
  NAND2X1 U74138 ( .A(n71245), .B(n71244), .Y(n71248) );
  NAND2X1 U74139 ( .A(n71246), .B(n43597), .Y(n71247) );
  NAND2X1 U74140 ( .A(n71248), .B(n71247), .Y(n71480) );
  NAND2X1 U74141 ( .A(n71249), .B(n42998), .Y(n71258) );
  NAND2X1 U74142 ( .A(n39556), .B(n71250), .Y(n71256) );
  NAND2X1 U74143 ( .A(n39066), .B(n39556), .Y(n71251) );
  NAND2X1 U74144 ( .A(n71252), .B(n71251), .Y(n71254) );
  NAND2X1 U74145 ( .A(n71254), .B(n71253), .Y(n71255) );
  NAND2X1 U74146 ( .A(n71256), .B(n71255), .Y(n71257) );
  XNOR2X1 U74147 ( .A(n41531), .B(n41667), .Y(n71366) );
  NAND2X1 U74148 ( .A(n72515), .B(n71259), .Y(n71260) );
  NAND2X1 U74149 ( .A(n71261), .B(n71260), .Y(n71263) );
  NAND2X1 U74150 ( .A(n71263), .B(n71262), .Y(n71268) );
  INVX1 U74151 ( .A(n71268), .Y(n71264) );
  NOR2X1 U74152 ( .A(n72515), .B(n71264), .Y(n71267) );
  INVX1 U74153 ( .A(n71271), .Y(n71272) );
  NOR2X1 U74154 ( .A(n72515), .B(n71272), .Y(n71266) );
  NOR2X1 U74155 ( .A(n71267), .B(n71266), .Y(n71270) );
  NAND2X1 U74156 ( .A(n71268), .B(n71271), .Y(n71269) );
  NAND2X1 U74157 ( .A(n71270), .B(n71269), .Y(n71487) );
  NAND2X1 U74158 ( .A(n71271), .B(n72196), .Y(n71276) );
  NAND2X1 U74159 ( .A(n72510), .B(n71272), .Y(n71274) );
  NAND2X1 U74160 ( .A(n71274), .B(n71273), .Y(n71275) );
  NAND2X1 U74161 ( .A(n71278), .B(n72202), .Y(n71283) );
  INVX1 U74162 ( .A(n71278), .Y(n71279) );
  NAND2X1 U74163 ( .A(n72200), .B(n71279), .Y(n71281) );
  NAND2X1 U74164 ( .A(n71281), .B(n71280), .Y(n71282) );
  XNOR2X1 U74165 ( .A(n71582), .B(n41823), .Y(n71364) );
  XNOR2X1 U74166 ( .A(n71290), .B(n41736), .Y(n71284) );
  XNOR2X1 U74167 ( .A(n71292), .B(n71284), .Y(n71285) );
  NAND2X1 U74168 ( .A(n71285), .B(n72233), .Y(n71289) );
  INVX1 U74169 ( .A(n72233), .Y(n72317) );
  INVX1 U74170 ( .A(n71285), .Y(n71286) );
  NAND2X1 U74171 ( .A(n72317), .B(n71286), .Y(n71287) );
  NAND2X1 U74172 ( .A(n41679), .B(n71287), .Y(n71288) );
  NAND2X1 U74173 ( .A(n71289), .B(n71288), .Y(n71504) );
  NAND2X1 U74174 ( .A(n71291), .B(n71290), .Y(n71296) );
  NAND2X1 U74175 ( .A(n71293), .B(n71292), .Y(n71294) );
  NAND2X1 U74176 ( .A(n41736), .B(n71294), .Y(n71295) );
  NAND2X1 U74177 ( .A(n71296), .B(n71295), .Y(n71559) );
  INVX1 U74178 ( .A(n71559), .Y(n71566) );
  NAND2X1 U74179 ( .A(n43500), .B(n44054), .Y(n71549) );
  NAND2X1 U74180 ( .A(n43614), .B(n43497), .Y(n72241) );
  INVX1 U74181 ( .A(n72241), .Y(n72347) );
  XNOR2X1 U74182 ( .A(n71549), .B(n72347), .Y(n71298) );
  XNOR2X1 U74183 ( .A(n72317), .B(n71298), .Y(n71336) );
  INVX1 U74184 ( .A(n71299), .Y(n71304) );
  NAND2X1 U74185 ( .A(n71304), .B(n71300), .Y(n71303) );
  NAND2X1 U74186 ( .A(n71301), .B(n71304), .Y(n71302) );
  NAND2X1 U74187 ( .A(n71303), .B(n71302), .Y(n71532) );
  NAND2X1 U74188 ( .A(n44024), .B(n43607), .Y(n71530) );
  NAND2X1 U74189 ( .A(n71304), .B(n43603), .Y(n72323) );
  NAND2X1 U74190 ( .A(n71305), .B(n71307), .Y(n71306) );
  NAND2X1 U74191 ( .A(n72425), .B(n71306), .Y(n71516) );
  INVX1 U74192 ( .A(n71307), .Y(n71520) );
  NAND2X1 U74193 ( .A(n72422), .B(n71886), .Y(n71310) );
  NAND2X1 U74194 ( .A(n72422), .B(n71308), .Y(n71309) );
  NAND2X1 U74195 ( .A(n71310), .B(n71309), .Y(n71312) );
  INVX1 U74196 ( .A(n71312), .Y(n71311) );
  NAND2X1 U74197 ( .A(n71311), .B(n72428), .Y(n71893) );
  NAND2X1 U74198 ( .A(n72425), .B(n71312), .Y(n71894) );
  XNOR2X1 U74199 ( .A(n71520), .B(n41703), .Y(n71517) );
  XNOR2X1 U74200 ( .A(n72434), .B(n71517), .Y(n71313) );
  XNOR2X1 U74201 ( .A(n72323), .B(n71511), .Y(n71318) );
  INVX1 U74202 ( .A(n72434), .Y(n72439) );
  NAND2X1 U74203 ( .A(n72439), .B(n71314), .Y(n71317) );
  NAND2X1 U74204 ( .A(n72439), .B(n71315), .Y(n71316) );
  NAND2X1 U74205 ( .A(n71317), .B(n71316), .Y(n71512) );
  NAND2X1 U74206 ( .A(n71320), .B(n71319), .Y(n71324) );
  NOR2X1 U74207 ( .A(n71320), .B(n71319), .Y(n71321) );
  NOR2X1 U74208 ( .A(n44028), .B(n71321), .Y(n71322) );
  NAND2X1 U74209 ( .A(n71322), .B(n39961), .Y(n71323) );
  NAND2X1 U74210 ( .A(n71324), .B(n71323), .Y(n71539) );
  NOR2X1 U74211 ( .A(n44053), .B(n36706), .Y(n71325) );
  XNOR2X1 U74212 ( .A(n71326), .B(n71325), .Y(n71548) );
  INVX1 U74213 ( .A(n71548), .Y(n71550) );
  NAND2X1 U74214 ( .A(n71327), .B(n71329), .Y(n71335) );
  INVX1 U74215 ( .A(n71328), .Y(n71330) );
  NOR2X1 U74216 ( .A(n71330), .B(n71329), .Y(n71332) );
  NAND2X1 U74217 ( .A(n71332), .B(n71331), .Y(n71333) );
  NAND2X1 U74218 ( .A(n41735), .B(n71333), .Y(n71334) );
  NAND2X1 U74219 ( .A(n71335), .B(n71334), .Y(n71547) );
  INVX1 U74220 ( .A(n71547), .Y(n71551) );
  XNOR2X1 U74221 ( .A(n71336), .B(n41254), .Y(n71337) );
  XNOR2X1 U74222 ( .A(n71566), .B(n71337), .Y(n71503) );
  INVX1 U74223 ( .A(n71338), .Y(n71351) );
  NAND2X1 U74224 ( .A(n71351), .B(n72225), .Y(n71347) );
  NAND2X1 U74225 ( .A(n72318), .B(n71338), .Y(n71345) );
  NAND2X1 U74226 ( .A(n72318), .B(n71339), .Y(n71340) );
  NAND2X1 U74227 ( .A(n71341), .B(n71340), .Y(n71343) );
  NAND2X1 U74228 ( .A(n71343), .B(n71342), .Y(n71344) );
  NAND2X1 U74229 ( .A(n71345), .B(n71344), .Y(n71346) );
  NAND2X1 U74230 ( .A(n71347), .B(n71346), .Y(n71493) );
  INVX1 U74231 ( .A(n71348), .Y(n72319) );
  XNOR2X1 U74232 ( .A(n71493), .B(n72319), .Y(n71349) );
  XNOR2X1 U74233 ( .A(n71494), .B(n71349), .Y(n71356) );
  NAND2X1 U74234 ( .A(n71357), .B(n72219), .Y(n71355) );
  INVX1 U74235 ( .A(n71357), .Y(n71358) );
  NAND2X1 U74236 ( .A(n72217), .B(n71358), .Y(n71353) );
  NAND2X1 U74237 ( .A(n71353), .B(n71352), .Y(n71354) );
  XNOR2X1 U74238 ( .A(n71356), .B(n41833), .Y(n71363) );
  NAND2X1 U74239 ( .A(n71357), .B(n72208), .Y(n71362) );
  NAND2X1 U74240 ( .A(n72212), .B(n71358), .Y(n71360) );
  NAND2X1 U74241 ( .A(n71360), .B(n71359), .Y(n71361) );
  XNOR2X1 U74242 ( .A(n71363), .B(n41832), .Y(n71577) );
  INVX1 U74243 ( .A(n71577), .Y(n71578) );
  XNOR2X1 U74244 ( .A(n71364), .B(n41676), .Y(n71365) );
  XNOR2X1 U74245 ( .A(n41821), .B(n71365), .Y(n71596) );
  XNOR2X1 U74246 ( .A(n71366), .B(n71479), .Y(n71367) );
  XNOR2X1 U74247 ( .A(n71480), .B(n71367), .Y(n71372) );
  NAND2X1 U74248 ( .A(n39236), .B(n40683), .Y(n71371) );
  NAND2X1 U74249 ( .A(n39788), .B(n43616), .Y(n71369) );
  NAND2X1 U74250 ( .A(n71369), .B(n71368), .Y(n71370) );
  XNOR2X1 U74251 ( .A(n71372), .B(n41784), .Y(n71614) );
  INVX1 U74252 ( .A(n71614), .Y(n71615) );
  XNOR2X1 U74253 ( .A(n43618), .B(n71615), .Y(n71475) );
  NAND2X1 U74254 ( .A(n41451), .B(n71373), .Y(n71375) );
  NAND2X1 U74255 ( .A(n71375), .B(n71374), .Y(n71608) );
  NAND2X1 U74256 ( .A(n43581), .B(n71608), .Y(n71377) );
  NAND2X1 U74257 ( .A(n43592), .B(n43585), .Y(n71376) );
  NOR2X1 U74258 ( .A(n71607), .B(n71377), .Y(n71381) );
  NAND2X1 U74259 ( .A(n71608), .B(n42994), .Y(n71378) );
  NAND2X1 U74260 ( .A(n71378), .B(n43585), .Y(n71379) );
  NOR2X1 U74261 ( .A(n71606), .B(n71379), .Y(n71380) );
  OR2X1 U74262 ( .A(n71381), .B(n71380), .Y(n71382) );
  NOR2X1 U74263 ( .A(n71383), .B(n71382), .Y(n71384) );
  NAND2X1 U74264 ( .A(n71386), .B(n43585), .Y(n71623) );
  NAND2X1 U74265 ( .A(n43581), .B(n71387), .Y(n71393) );
  NAND2X1 U74266 ( .A(n71388), .B(n43585), .Y(n71391) );
  OR2X1 U74267 ( .A(n43589), .B(n71388), .Y(n71389) );
  NAND2X1 U74268 ( .A(n41129), .B(n71389), .Y(n71390) );
  NAND2X1 U74269 ( .A(n71391), .B(n71390), .Y(n71392) );
  NAND2X1 U74270 ( .A(n71393), .B(n71392), .Y(n71624) );
  NAND2X1 U74271 ( .A(n71623), .B(n71624), .Y(n71452) );
  XNOR2X1 U74272 ( .A(n43537), .B(n43579), .Y(n71638) );
  XNOR2X1 U74273 ( .A(n71638), .B(n43564), .Y(n71394) );
  XNOR2X1 U74274 ( .A(n71452), .B(n71394), .Y(n71395) );
  XNOR2X1 U74275 ( .A(n71622), .B(n71395), .Y(n71665) );
  XNOR2X1 U74276 ( .A(n71663), .B(n71665), .Y(n71396) );
  XOR2X1 U74277 ( .A(n71654), .B(n71396), .Y(n71467) );
  XNOR2X1 U74278 ( .A(n71397), .B(n71467), .Y(n71398) );
  XNOR2X1 U74279 ( .A(n71469), .B(n71398), .Y(n71438) );
  XNOR2X1 U74280 ( .A(n71438), .B(n72088), .Y(n71399) );
  XNOR2X1 U74281 ( .A(n71689), .B(n43654), .Y(n71400) );
  XNOR2X1 U74282 ( .A(n71690), .B(n71400), .Y(n71401) );
  XNOR2X1 U74283 ( .A(n41073), .B(n71401), .Y(n71428) );
  XNOR2X1 U74284 ( .A(n71402), .B(n71428), .Y(n71403) );
  XNOR2X1 U74285 ( .A(n71413), .B(n71405), .Y(n71713) );
  XNOR2X1 U74286 ( .A(n43715), .B(n72106), .Y(n71406) );
  XNOR2X1 U74287 ( .A(n71407), .B(n71406), .Y(n71412) );
  XNOR2X1 U74288 ( .A(n71408), .B(n36353), .Y(n71409) );
  XNOR2X1 U74289 ( .A(n71410), .B(n71409), .Y(n71411) );
  MX2X1 U74290 ( .A(n71412), .B(n71411), .S0(n43718), .Y(u_muldiv_result_r[28]) );
  NAND2X1 U74291 ( .A(u_muldiv_mult_result_q[28]), .B(n44631), .Y(n13875) );
  XNOR2X1 U74292 ( .A(n43509), .B(n72101), .Y(n71415) );
  NOR2X1 U74293 ( .A(n39922), .B(n40569), .Y(n71416) );
  NAND2X1 U74294 ( .A(n71416), .B(n41019), .Y(n71417) );
  NAND2X1 U74295 ( .A(n71417), .B(n43697), .Y(n71420) );
  NAND2X1 U74296 ( .A(n71418), .B(n43697), .Y(n71419) );
  NAND2X1 U74297 ( .A(n71420), .B(n71419), .Y(n72102) );
  NAND2X1 U74298 ( .A(n71424), .B(n71423), .Y(n71425) );
  NOR2X1 U74299 ( .A(n71426), .B(n71425), .Y(n71427) );
  XNOR2X1 U74300 ( .A(n43524), .B(n71427), .Y(n71429) );
  INVX1 U74301 ( .A(n71428), .Y(n71699) );
  NOR2X1 U74302 ( .A(n43678), .B(n71735), .Y(n71432) );
  NAND2X1 U74303 ( .A(n71434), .B(n71435), .Y(n71436) );
  INVX1 U74304 ( .A(n71735), .Y(n71437) );
  XNOR2X1 U74305 ( .A(n71690), .B(n43673), .Y(n71440) );
  XOR2X1 U74306 ( .A(n71787), .B(n71440), .Y(n71441) );
  NAND2X1 U74307 ( .A(n43642), .B(n71441), .Y(n71764) );
  XNOR2X1 U74308 ( .A(n71662), .B(n72078), .Y(n71443) );
  XNOR2X1 U74309 ( .A(n71467), .B(n71443), .Y(n71444) );
  XNOR2X1 U74310 ( .A(n71444), .B(n71469), .Y(n71445) );
  NAND2X1 U74311 ( .A(n71446), .B(n43632), .Y(n71451) );
  INVX1 U74312 ( .A(n71446), .Y(n71447) );
  NAND2X1 U74313 ( .A(n71447), .B(n43635), .Y(n71448) );
  NAND2X1 U74314 ( .A(n71449), .B(n71448), .Y(n71450) );
  NAND2X1 U74315 ( .A(n71451), .B(n71450), .Y(n72084) );
  NOR2X1 U74316 ( .A(n71461), .B(n71662), .Y(n71458) );
  INVX1 U74317 ( .A(n71654), .Y(n71661) );
  INVX1 U74318 ( .A(n71452), .Y(n71635) );
  XNOR2X1 U74319 ( .A(n71638), .B(n71622), .Y(n71453) );
  XNOR2X1 U74320 ( .A(n71635), .B(n71453), .Y(n71454) );
  XNOR2X1 U74321 ( .A(n71454), .B(n38840), .Y(n71455) );
  XNOR2X1 U74322 ( .A(n71661), .B(n71455), .Y(n71797) );
  INVX1 U74323 ( .A(n71797), .Y(n71456) );
  NAND2X1 U74324 ( .A(n41012), .B(n71456), .Y(n71800) );
  NOR2X1 U74325 ( .A(n71461), .B(n71800), .Y(n71457) );
  NOR2X1 U74326 ( .A(n71458), .B(n71457), .Y(n71466) );
  NOR2X1 U74327 ( .A(n41012), .B(n71459), .Y(n71460) );
  NAND2X1 U74328 ( .A(n71460), .B(n71797), .Y(n71463) );
  NAND2X1 U74329 ( .A(n71461), .B(n71662), .Y(n71462) );
  NAND2X1 U74330 ( .A(n71463), .B(n71462), .Y(n71464) );
  NAND2X1 U74331 ( .A(n71464), .B(n71800), .Y(n71465) );
  NAND2X1 U74332 ( .A(n71466), .B(n71465), .Y(n71474) );
  XNOR2X1 U74333 ( .A(n71467), .B(n71799), .Y(n71470) );
  NAND2X1 U74334 ( .A(n71470), .B(n43623), .Y(n71468) );
  NAND2X1 U74335 ( .A(n71469), .B(n71468), .Y(n71804) );
  INVX1 U74336 ( .A(n71470), .Y(n71471) );
  NAND2X1 U74337 ( .A(n43619), .B(n71471), .Y(n71805) );
  INVX1 U74338 ( .A(n71805), .Y(n71472) );
  NOR2X1 U74339 ( .A(n38863), .B(n71472), .Y(n71473) );
  XNOR2X1 U74340 ( .A(n71474), .B(n71473), .Y(n71659) );
  INVX1 U74341 ( .A(n71475), .Y(n71629) );
  XNOR2X1 U74342 ( .A(n41670), .B(n71629), .Y(n71605) );
  NAND2X1 U74343 ( .A(n43567), .B(n71605), .Y(n71478) );
  INVX1 U74344 ( .A(n71605), .Y(n71612) );
  NAND2X1 U74345 ( .A(n71612), .B(n40670), .Y(n71476) );
  NAND2X1 U74346 ( .A(n41800), .B(n71476), .Y(n71477) );
  NAND2X1 U74347 ( .A(n71478), .B(n71477), .Y(n72031) );
  XNOR2X1 U74348 ( .A(n72031), .B(n43583), .Y(n71621) );
  XNOR2X1 U74349 ( .A(n71479), .B(n41667), .Y(n71590) );
  NAND2X1 U74350 ( .A(n43602), .B(n71590), .Y(n71484) );
  INVX1 U74351 ( .A(n71480), .Y(n71482) );
  INVX1 U74352 ( .A(n71590), .Y(n71591) );
  NAND2X1 U74353 ( .A(n71591), .B(n43597), .Y(n71481) );
  NAND2X1 U74354 ( .A(n71482), .B(n71481), .Y(n71483) );
  NAND2X1 U74355 ( .A(n71484), .B(n71483), .Y(n72012) );
  INVX1 U74356 ( .A(n72012), .Y(n72004) );
  XNOR2X1 U74357 ( .A(n41823), .B(n41734), .Y(n71485) );
  XNOR2X1 U74358 ( .A(n71485), .B(n71578), .Y(n71486) );
  XNOR2X1 U74359 ( .A(n41821), .B(n71486), .Y(n71488) );
  NAND2X1 U74360 ( .A(n72515), .B(n71488), .Y(n71492) );
  INVX1 U74361 ( .A(n71487), .Y(n71597) );
  INVX1 U74362 ( .A(n71488), .Y(n71489) );
  NAND2X1 U74363 ( .A(n71489), .B(n43000), .Y(n71490) );
  NAND2X1 U74364 ( .A(n71597), .B(n71490), .Y(n71491) );
  NAND2X1 U74365 ( .A(n71492), .B(n71491), .Y(n71996) );
  INVX1 U74366 ( .A(n71493), .Y(n71508) );
  XNOR2X1 U74367 ( .A(n71494), .B(n71508), .Y(n71498) );
  NAND2X1 U74368 ( .A(n72212), .B(n71498), .Y(n71497) );
  INVX1 U74369 ( .A(n71498), .Y(n71499) );
  NAND2X1 U74370 ( .A(n71499), .B(n72208), .Y(n71495) );
  NAND2X1 U74371 ( .A(n41832), .B(n71495), .Y(n71496) );
  NAND2X1 U74372 ( .A(n71497), .B(n71496), .Y(n71979) );
  NAND2X1 U74373 ( .A(n72217), .B(n71498), .Y(n71502) );
  NAND2X1 U74374 ( .A(n71499), .B(n72219), .Y(n71500) );
  NAND2X1 U74375 ( .A(n41833), .B(n71500), .Y(n71501) );
  NAND2X1 U74376 ( .A(n71502), .B(n71501), .Y(n71972) );
  INVX1 U74377 ( .A(n71972), .Y(n71963) );
  INVX1 U74378 ( .A(n71504), .Y(n71570) );
  NAND2X1 U74379 ( .A(n72318), .B(n71505), .Y(n71510) );
  INVX1 U74380 ( .A(n71505), .Y(n71506) );
  NAND2X1 U74381 ( .A(n71506), .B(n72225), .Y(n71507) );
  NAND2X1 U74382 ( .A(n71508), .B(n71507), .Y(n71509) );
  NAND2X1 U74383 ( .A(n71510), .B(n71509), .Y(n71956) );
  INVX1 U74384 ( .A(n71956), .Y(n71961) );
  XNOR2X1 U74385 ( .A(n72319), .B(n71961), .Y(n71574) );
  INVX1 U74386 ( .A(n72323), .Y(n72447) );
  NAND2X1 U74387 ( .A(n72447), .B(n71511), .Y(n71514) );
  NAND2X1 U74388 ( .A(n72447), .B(n71512), .Y(n71513) );
  NAND2X1 U74389 ( .A(n71514), .B(n71513), .Y(n71905) );
  INVX1 U74390 ( .A(n71905), .Y(n71910) );
  NAND2X1 U74391 ( .A(n44047), .B(n43607), .Y(n71920) );
  XNOR2X1 U74392 ( .A(n71920), .B(n41737), .Y(n71515) );
  XNOR2X1 U74393 ( .A(n71910), .B(n71515), .Y(n71537) );
  NOR2X1 U74394 ( .A(n72434), .B(n71516), .Y(n71519) );
  NOR2X1 U74395 ( .A(n71517), .B(n72434), .Y(n71518) );
  NAND2X1 U74396 ( .A(n71520), .B(n71893), .Y(n71521) );
  NAND2X1 U74397 ( .A(n71521), .B(n71894), .Y(n71899) );
  XNOR2X1 U74398 ( .A(n71899), .B(n41703), .Y(n71528) );
  XNOR2X1 U74399 ( .A(n41686), .B(n71856), .Y(n71860) );
  XNOR2X1 U74400 ( .A(n71860), .B(n72327), .Y(n71522) );
  XNOR2X1 U74401 ( .A(n71523), .B(n71522), .Y(n71867) );
  XNOR2X1 U74402 ( .A(n71867), .B(n72291), .Y(n71524) );
  XNOR2X1 U74403 ( .A(n72280), .B(n71872), .Y(n71525) );
  XNOR2X1 U74404 ( .A(n41694), .B(n71876), .Y(n71881) );
  XNOR2X1 U74405 ( .A(n41701), .B(n41512), .Y(n71885) );
  XNOR2X1 U74406 ( .A(n72434), .B(n72323), .Y(n71526) );
  XOR2X1 U74407 ( .A(n41511), .B(n71526), .Y(n71527) );
  XNOR2X1 U74408 ( .A(n71528), .B(n71527), .Y(n71529) );
  INVX1 U74409 ( .A(n71530), .Y(n71533) );
  NAND2X1 U74410 ( .A(n71533), .B(n43603), .Y(n72451) );
  INVX1 U74411 ( .A(n72451), .Y(n72456) );
  XNOR2X1 U74412 ( .A(n71904), .B(n72456), .Y(n71909) );
  NAND2X1 U74413 ( .A(n71533), .B(n71531), .Y(n71535) );
  NAND2X1 U74414 ( .A(n71533), .B(n71532), .Y(n71534) );
  XNOR2X1 U74415 ( .A(n71909), .B(n41710), .Y(n71536) );
  XNOR2X1 U74416 ( .A(n71537), .B(n71536), .Y(n71545) );
  INVX1 U74417 ( .A(n71538), .Y(n71540) );
  NAND2X1 U74418 ( .A(n71540), .B(n71539), .Y(n71544) );
  NOR2X1 U74419 ( .A(n71540), .B(n71539), .Y(n71541) );
  NOR2X1 U74420 ( .A(n44053), .B(n71541), .Y(n71542) );
  NAND2X1 U74421 ( .A(n71542), .B(n43517), .Y(n71543) );
  NAND2X1 U74422 ( .A(n71544), .B(n71543), .Y(n71912) );
  INVX1 U74423 ( .A(n71912), .Y(n71915) );
  XNOR2X1 U74424 ( .A(n71545), .B(n71915), .Y(n71929) );
  INVX1 U74425 ( .A(n71929), .Y(n71930) );
  NAND2X1 U74426 ( .A(n43614), .B(n43501), .Y(n72489) );
  INVX1 U74427 ( .A(n72489), .Y(n72486) );
  XNOR2X1 U74428 ( .A(n72317), .B(n72347), .Y(n71555) );
  NAND2X1 U74429 ( .A(n71548), .B(n71547), .Y(n71554) );
  INVX1 U74430 ( .A(n71549), .Y(n71557) );
  NAND2X1 U74431 ( .A(n71551), .B(n71550), .Y(n71552) );
  NAND2X1 U74432 ( .A(n71557), .B(n71552), .Y(n71553) );
  NAND2X1 U74433 ( .A(n71554), .B(n71553), .Y(n71931) );
  INVX1 U74434 ( .A(n71931), .Y(n71936) );
  XNOR2X1 U74435 ( .A(n71555), .B(n71936), .Y(n71556) );
  XNOR2X1 U74436 ( .A(n41706), .B(n71556), .Y(n71563) );
  XNOR2X1 U74437 ( .A(n41254), .B(n71557), .Y(n71564) );
  INVX1 U74438 ( .A(n71564), .Y(n71558) );
  NAND2X1 U74439 ( .A(n72347), .B(n71558), .Y(n71562) );
  NAND2X1 U74440 ( .A(n71564), .B(n72241), .Y(n71560) );
  NAND2X1 U74441 ( .A(n71560), .B(n71559), .Y(n71561) );
  NAND2X1 U74442 ( .A(n71562), .B(n71561), .Y(n71948) );
  INVX1 U74443 ( .A(n71948), .Y(n71938) );
  XNOR2X1 U74444 ( .A(n71563), .B(n71938), .Y(n71573) );
  XNOR2X1 U74445 ( .A(n71564), .B(n72347), .Y(n71565) );
  XNOR2X1 U74446 ( .A(n71566), .B(n71565), .Y(n71567) );
  NAND2X1 U74447 ( .A(n72317), .B(n71567), .Y(n71572) );
  INVX1 U74448 ( .A(n71567), .Y(n71568) );
  NAND2X1 U74449 ( .A(n71568), .B(n72233), .Y(n71569) );
  NAND2X1 U74450 ( .A(n71570), .B(n71569), .Y(n71571) );
  NAND2X1 U74451 ( .A(n71572), .B(n71571), .Y(n71941) );
  INVX1 U74452 ( .A(n71955), .Y(n71954) );
  XNOR2X1 U74453 ( .A(n71574), .B(n41687), .Y(n71575) );
  XNOR2X1 U74454 ( .A(n71963), .B(n71575), .Y(n71978) );
  XNOR2X1 U74455 ( .A(n72202), .B(n71978), .Y(n71576) );
  XOR2X1 U74456 ( .A(n71979), .B(n71576), .Y(n71833) );
  NAND2X1 U74457 ( .A(n72200), .B(n71577), .Y(n71581) );
  NAND2X1 U74458 ( .A(n71578), .B(n72202), .Y(n71579) );
  NAND2X1 U74459 ( .A(n41823), .B(n71579), .Y(n71580) );
  NAND2X1 U74460 ( .A(n71581), .B(n71580), .Y(n71982) );
  XNOR2X1 U74461 ( .A(n71982), .B(n71582), .Y(n71583) );
  XNOR2X1 U74462 ( .A(n71833), .B(n71583), .Y(n71997) );
  XNOR2X1 U74463 ( .A(n41676), .B(n41823), .Y(n71584) );
  NAND2X1 U74464 ( .A(n72510), .B(n71584), .Y(n71588) );
  INVX1 U74465 ( .A(n71584), .Y(n71585) );
  NAND2X1 U74466 ( .A(n71585), .B(n72196), .Y(n71586) );
  NAND2X1 U74467 ( .A(n41821), .B(n71586), .Y(n71587) );
  NAND2X1 U74468 ( .A(n71588), .B(n71587), .Y(n71995) );
  INVX1 U74469 ( .A(n71990), .Y(n71989) );
  XNOR2X1 U74470 ( .A(n39556), .B(n71989), .Y(n71821) );
  INVX1 U74471 ( .A(n71821), .Y(n71589) );
  XNOR2X1 U74472 ( .A(n72004), .B(n71589), .Y(n71595) );
  NAND2X1 U74473 ( .A(n43615), .B(n71590), .Y(n71594) );
  NAND2X1 U74474 ( .A(n71591), .B(n40683), .Y(n71592) );
  NAND2X1 U74475 ( .A(n41784), .B(n71592), .Y(n71593) );
  NAND2X1 U74476 ( .A(n71594), .B(n71593), .Y(n72002) );
  INVX1 U74477 ( .A(n72002), .Y(n72018) );
  XNOR2X1 U74478 ( .A(n71595), .B(n72018), .Y(n71604) );
  NAND2X1 U74479 ( .A(n42187), .B(n71598), .Y(n71602) );
  INVX1 U74480 ( .A(n71598), .Y(n71599) );
  NAND2X1 U74481 ( .A(n71599), .B(n42998), .Y(n71600) );
  NAND2X1 U74482 ( .A(n41667), .B(n71600), .Y(n71601) );
  NAND2X1 U74483 ( .A(n71602), .B(n71601), .Y(n71998) );
  XNOR2X1 U74484 ( .A(n71820), .B(n43618), .Y(n71603) );
  XNOR2X1 U74485 ( .A(n71604), .B(n71603), .Y(n71811) );
  NAND2X1 U74486 ( .A(n71606), .B(n42993), .Y(n71611) );
  NAND2X1 U74487 ( .A(n43592), .B(n71607), .Y(n71609) );
  NAND2X1 U74488 ( .A(n71609), .B(n71608), .Y(n71610) );
  NAND2X1 U74489 ( .A(n71612), .B(n42994), .Y(n71613) );
  XNOR2X1 U74490 ( .A(n71811), .B(n38933), .Y(n71620) );
  NAND2X1 U74491 ( .A(n43617), .B(n71614), .Y(n71618) );
  NAND2X1 U74492 ( .A(n71615), .B(n42997), .Y(n71616) );
  NAND2X1 U74493 ( .A(n41670), .B(n71616), .Y(n71617) );
  NAND2X1 U74494 ( .A(n71618), .B(n71617), .Y(n72021) );
  XNOR2X1 U74495 ( .A(n72021), .B(n72353), .Y(n71619) );
  XNOR2X1 U74496 ( .A(n71620), .B(n71619), .Y(n72045) );
  INVX1 U74497 ( .A(n72045), .Y(n72032) );
  XNOR2X1 U74498 ( .A(n71621), .B(n72032), .Y(n72058) );
  INVX1 U74499 ( .A(n71625), .Y(n71648) );
  NAND2X1 U74500 ( .A(n43577), .B(n71648), .Y(n71628) );
  NAND2X1 U74501 ( .A(n71625), .B(n43573), .Y(n71626) );
  NAND2X1 U74502 ( .A(n38840), .B(n71626), .Y(n71627) );
  NAND2X1 U74503 ( .A(n71628), .B(n71627), .Y(n72061) );
  INVX1 U74504 ( .A(n72061), .Y(n72051) );
  XNOR2X1 U74505 ( .A(n72058), .B(n72051), .Y(n71640) );
  XNOR2X1 U74506 ( .A(n41800), .B(n71631), .Y(n71632) );
  NAND2X1 U74507 ( .A(n43581), .B(n71632), .Y(n71637) );
  INVX1 U74508 ( .A(n71632), .Y(n71633) );
  NAND2X1 U74509 ( .A(n71633), .B(n43585), .Y(n71634) );
  NAND2X1 U74510 ( .A(n71635), .B(n71634), .Y(n71636) );
  NAND2X1 U74511 ( .A(n71637), .B(n71636), .Y(n72048) );
  XNOR2X1 U74512 ( .A(n72048), .B(n71638), .Y(n71639) );
  XNOR2X1 U74513 ( .A(n71640), .B(n71639), .Y(n72039) );
  INVX1 U74514 ( .A(n71641), .Y(n71644) );
  NAND2X1 U74515 ( .A(n71642), .B(n43573), .Y(n71643) );
  NOR2X1 U74516 ( .A(n71644), .B(n71643), .Y(n71646) );
  NAND2X1 U74517 ( .A(n71646), .B(n71645), .Y(n71647) );
  NAND2X1 U74518 ( .A(n71648), .B(n71647), .Y(n71650) );
  INVX1 U74519 ( .A(n71650), .Y(n71649) );
  NAND2X1 U74520 ( .A(n71649), .B(n43536), .Y(n71796) );
  NAND2X1 U74521 ( .A(n71796), .B(n39629), .Y(n71653) );
  NAND2X1 U74522 ( .A(n71650), .B(n43539), .Y(n71651) );
  NAND2X1 U74523 ( .A(n71661), .B(n71651), .Y(n71795) );
  INVX1 U74524 ( .A(n71795), .Y(n71652) );
  NOR2X1 U74525 ( .A(n71653), .B(n71652), .Y(n71658) );
  NOR2X1 U74526 ( .A(n39629), .B(n71654), .Y(n71656) );
  NOR2X1 U74527 ( .A(n39629), .B(n71796), .Y(n71655) );
  OR2X1 U74528 ( .A(n71656), .B(n71655), .Y(n71657) );
  XNOR2X1 U74529 ( .A(n71659), .B(n72079), .Y(n71675) );
  INVX1 U74530 ( .A(n71675), .Y(n71669) );
  XNOR2X1 U74531 ( .A(n71662), .B(n71661), .Y(n71667) );
  XNOR2X1 U74532 ( .A(n43623), .B(n71663), .Y(n71664) );
  XOR2X1 U74533 ( .A(n71665), .B(n71664), .Y(n71666) );
  NOR2X1 U74534 ( .A(n71669), .B(n71672), .Y(n71679) );
  INVX1 U74535 ( .A(n71670), .Y(n71671) );
  NAND2X1 U74536 ( .A(n43544), .B(n71671), .Y(n71673) );
  NAND2X1 U74537 ( .A(n71672), .B(n71673), .Y(n72077) );
  OR2X1 U74538 ( .A(n71675), .B(n72077), .Y(n71677) );
  INVX1 U74539 ( .A(n71673), .Y(n71674) );
  NAND2X1 U74540 ( .A(n71675), .B(n71674), .Y(n71676) );
  NAND2X1 U74541 ( .A(n71677), .B(n71676), .Y(n71678) );
  NOR2X1 U74542 ( .A(n71679), .B(n71678), .Y(n71767) );
  NOR2X1 U74543 ( .A(n38555), .B(n38128), .Y(n71680) );
  NAND2X1 U74544 ( .A(n71680), .B(n71787), .Y(n71683) );
  NOR2X1 U74545 ( .A(n43665), .B(n71787), .Y(n71681) );
  NAND2X1 U74546 ( .A(n71681), .B(n40503), .Y(n71682) );
  NAND2X1 U74547 ( .A(n71683), .B(n71682), .Y(n71768) );
  XNOR2X1 U74548 ( .A(n43524), .B(n43643), .Y(n71684) );
  XNOR2X1 U74549 ( .A(n71684), .B(n43654), .Y(n71685) );
  XNOR2X1 U74550 ( .A(n71768), .B(n71685), .Y(n71686) );
  XNOR2X1 U74551 ( .A(n71791), .B(n71686), .Y(n71687) );
  NAND2X1 U74552 ( .A(n71688), .B(n39725), .Y(n71691) );
  NAND2X1 U74553 ( .A(n71752), .B(n71698), .Y(n71755) );
  NOR2X1 U74554 ( .A(n71695), .B(n71755), .Y(n71694) );
  NOR2X1 U74555 ( .A(n41404), .B(n41340), .Y(n71692) );
  NOR2X1 U74556 ( .A(n71692), .B(n71695), .Y(n71693) );
  INVX1 U74557 ( .A(n71755), .Y(n71773) );
  XNOR2X1 U74558 ( .A(n71700), .B(n43679), .Y(n71701) );
  XNOR2X1 U74559 ( .A(n71733), .B(n71701), .Y(n71702) );
  XNOR2X1 U74560 ( .A(n40143), .B(n71702), .Y(n71730) );
  XNOR2X1 U74561 ( .A(n39866), .B(n72101), .Y(n71723) );
  INVX1 U74562 ( .A(n71723), .Y(n71722) );
  NOR2X1 U74563 ( .A(n39255), .B(n36576), .Y(n71705) );
  NOR2X1 U74564 ( .A(n71723), .B(n41027), .Y(n71708) );
  NOR2X1 U74565 ( .A(n71706), .B(n43512), .Y(n71707) );
  XNOR2X1 U74566 ( .A(n43702), .B(n72097), .Y(n71709) );
  XNOR2X1 U74567 ( .A(n71730), .B(n71709), .Y(n72105) );
  XNOR2X1 U74568 ( .A(n72105), .B(n43707), .Y(n71710) );
  XNOR2X1 U74569 ( .A(n41014), .B(n71710), .Y(n71716) );
  NAND2X1 U74570 ( .A(n41018), .B(n71711), .Y(n71714) );
  NOR2X1 U74571 ( .A(n71713), .B(n71714), .Y(n71712) );
  NAND2X1 U74572 ( .A(n40455), .B(n36565), .Y(n72644) );
  XNOR2X1 U74573 ( .A(n71716), .B(n40192), .Y(n71721) );
  XNOR2X1 U74574 ( .A(n71718), .B(n71717), .Y(n71719) );
  XNOR2X1 U74575 ( .A(n42125), .B(n71719), .Y(n71720) );
  MX2X1 U74576 ( .A(n71721), .B(n71720), .S0(n43718), .Y(u_muldiv_result_r[29]) );
  NAND2X1 U74577 ( .A(u_muldiv_mult_result_q[29]), .B(n44631), .Y(n13864) );
  NOR2X1 U74578 ( .A(n71722), .B(n43512), .Y(n71729) );
  NOR2X1 U74579 ( .A(n43507), .B(n71723), .Y(n71727) );
  INVX1 U74580 ( .A(n71724), .Y(n71725) );
  NOR2X1 U74581 ( .A(n41027), .B(n71725), .Y(n71726) );
  NOR2X1 U74582 ( .A(n71727), .B(n71726), .Y(n71728) );
  NOR2X1 U74583 ( .A(n71729), .B(n71728), .Y(n71732) );
  NAND2X1 U74584 ( .A(n43507), .B(n71730), .Y(n71731) );
  INVX1 U74585 ( .A(n72686), .Y(n72694) );
  NAND2X1 U74586 ( .A(n39227), .B(n71735), .Y(n71738) );
  NAND2X1 U74587 ( .A(n43506), .B(n71736), .Y(n71737) );
  NAND2X1 U74588 ( .A(n71738), .B(n71737), .Y(n71739) );
  NOR2X1 U74589 ( .A(n71740), .B(n71739), .Y(n71743) );
  NAND2X1 U74590 ( .A(n71743), .B(n71742), .Y(n72096) );
  INVX1 U74591 ( .A(n71791), .Y(n72605) );
  XNOR2X1 U74592 ( .A(n71768), .B(n71744), .Y(n71745) );
  XNOR2X1 U74593 ( .A(n72605), .B(n71745), .Y(n71746) );
  XNOR2X1 U74594 ( .A(n38194), .B(n71746), .Y(n71756) );
  NOR2X1 U74595 ( .A(n38930), .B(n71748), .Y(n71750) );
  NAND2X1 U74596 ( .A(n71750), .B(n71749), .Y(n71751) );
  NAND2X1 U74597 ( .A(n71751), .B(n43656), .Y(n71754) );
  NAND2X1 U74598 ( .A(n71752), .B(n43656), .Y(n71753) );
  XNOR2X1 U74599 ( .A(n71756), .B(n41116), .Y(n72132) );
  INVX1 U74600 ( .A(n72132), .Y(n72131) );
  NAND2X1 U74601 ( .A(n43521), .B(n72131), .Y(n71758) );
  NOR2X1 U74602 ( .A(n71758), .B(n71757), .Y(n71761) );
  NAND2X1 U74603 ( .A(n72132), .B(n43527), .Y(n71759) );
  NOR2X1 U74604 ( .A(n39412), .B(n71759), .Y(n71760) );
  NOR2X1 U74605 ( .A(n71761), .B(n71760), .Y(n72095) );
  NAND2X1 U74606 ( .A(n71763), .B(n71764), .Y(n71765) );
  NOR2X1 U74607 ( .A(n38165), .B(n71765), .Y(n71772) );
  XNOR2X1 U74608 ( .A(n72084), .B(n43643), .Y(n71766) );
  XNOR2X1 U74609 ( .A(n71767), .B(n71766), .Y(n71770) );
  INVX1 U74610 ( .A(n71768), .Y(n71769) );
  XNOR2X1 U74611 ( .A(n71770), .B(n71769), .Y(n71771) );
  XNOR2X1 U74612 ( .A(n71772), .B(n71771), .Y(n71778) );
  XNOR2X1 U74613 ( .A(n38047), .B(n43654), .Y(n71777) );
  INVX1 U74614 ( .A(n71777), .Y(n71775) );
  NOR2X1 U74615 ( .A(n71773), .B(n71775), .Y(n71774) );
  NOR2X1 U74616 ( .A(n71777), .B(n38941), .Y(n71780) );
  NAND2X1 U74617 ( .A(n41116), .B(n71779), .Y(n72136) );
  NAND2X1 U74618 ( .A(n71780), .B(n72136), .Y(n71781) );
  NAND2X1 U74619 ( .A(n43643), .B(n71791), .Y(n71785) );
  NAND2X1 U74620 ( .A(n72605), .B(n39301), .Y(n71783) );
  NAND2X1 U74621 ( .A(n71783), .B(n71782), .Y(n71784) );
  NAND2X1 U74622 ( .A(n71785), .B(n71784), .Y(n72669) );
  INVX1 U74623 ( .A(n72669), .Y(n72617) );
  NAND2X1 U74624 ( .A(n43665), .B(n71791), .Y(n72608) );
  INVX1 U74625 ( .A(n71787), .Y(n71786) );
  NAND2X1 U74626 ( .A(n43664), .B(n71786), .Y(n71790) );
  NAND2X1 U74627 ( .A(n71787), .B(n38555), .Y(n71788) );
  NAND2X1 U74628 ( .A(n40503), .B(n71788), .Y(n71789) );
  NAND2X1 U74629 ( .A(n71790), .B(n71789), .Y(n72606) );
  OR2X1 U74630 ( .A(n43667), .B(n71791), .Y(n71792) );
  NAND2X1 U74631 ( .A(n72606), .B(n71792), .Y(n71793) );
  NAND2X1 U74632 ( .A(n72608), .B(n71793), .Y(n72092) );
  XNOR2X1 U74633 ( .A(n71794), .B(n72039), .Y(n71803) );
  NAND2X1 U74634 ( .A(n71796), .B(n71795), .Y(n72054) );
  NAND2X1 U74635 ( .A(n71797), .B(n39629), .Y(n71798) );
  NAND2X1 U74636 ( .A(n71799), .B(n71798), .Y(n71801) );
  XNOR2X1 U74637 ( .A(n72054), .B(n38683), .Y(n71802) );
  XNOR2X1 U74638 ( .A(n71803), .B(n71802), .Y(n71806) );
  NAND2X1 U74639 ( .A(n71805), .B(n71804), .Y(n72560) );
  XNOR2X1 U74640 ( .A(n71806), .B(n38169), .Y(n71807) );
  INVX1 U74641 ( .A(n71807), .Y(n71808) );
  NAND2X1 U74642 ( .A(n71808), .B(n43547), .Y(n71809) );
  XNOR2X1 U74643 ( .A(n71810), .B(n72154), .Y(n72076) );
  INVX1 U74644 ( .A(n71813), .Y(n71812) );
  NAND2X1 U74645 ( .A(n43592), .B(n71812), .Y(n71817) );
  NAND2X1 U74646 ( .A(n71813), .B(n42993), .Y(n71815) );
  NAND2X1 U74647 ( .A(n71815), .B(n71814), .Y(n71816) );
  NAND2X1 U74648 ( .A(n71817), .B(n71816), .Y(n72188) );
  XNOR2X1 U74649 ( .A(n72188), .B(n43594), .Y(n71818) );
  XNOR2X1 U74650 ( .A(n71819), .B(n71818), .Y(n72030) );
  XNOR2X1 U74651 ( .A(n71821), .B(n71820), .Y(n71822) );
  XOR2X1 U74652 ( .A(n72012), .B(n71822), .Y(n72017) );
  XNOR2X1 U74653 ( .A(n42996), .B(n43594), .Y(n71823) );
  XNOR2X1 U74654 ( .A(n72017), .B(n71823), .Y(n71825) );
  XNOR2X1 U74655 ( .A(n72021), .B(n72018), .Y(n71824) );
  XNOR2X1 U74656 ( .A(n71825), .B(n71824), .Y(n71826) );
  XNOR2X1 U74657 ( .A(n38933), .B(n71826), .Y(n71827) );
  NAND2X1 U74658 ( .A(n43567), .B(n71827), .Y(n71831) );
  INVX1 U74659 ( .A(n71827), .Y(n71828) );
  NAND2X1 U74660 ( .A(n71828), .B(n40670), .Y(n71829) );
  NAND2X1 U74661 ( .A(n71829), .B(n72031), .Y(n71830) );
  NAND2X1 U74662 ( .A(n71831), .B(n71830), .Y(n72163) );
  INVX1 U74663 ( .A(n71832), .Y(n72316) );
  INVX1 U74664 ( .A(n71839), .Y(n71838) );
  NAND2X1 U74665 ( .A(n72510), .B(n71838), .Y(n71836) );
  NAND2X1 U74666 ( .A(n71839), .B(n72196), .Y(n71834) );
  NAND2X1 U74667 ( .A(n71834), .B(n71995), .Y(n71835) );
  NAND2X1 U74668 ( .A(n71836), .B(n71835), .Y(n72509) );
  XNOR2X1 U74669 ( .A(n72509), .B(n72510), .Y(n71837) );
  XNOR2X1 U74670 ( .A(n72316), .B(n71837), .Y(n71988) );
  NAND2X1 U74671 ( .A(n72515), .B(n71838), .Y(n71842) );
  NAND2X1 U74672 ( .A(n71839), .B(n43000), .Y(n71840) );
  NAND2X1 U74673 ( .A(n71840), .B(n71996), .Y(n71841) );
  NAND2X1 U74674 ( .A(n71842), .B(n71841), .Y(n72512) );
  INVX1 U74675 ( .A(n71920), .Y(n71923) );
  NAND2X1 U74676 ( .A(n71923), .B(n43603), .Y(n72464) );
  XNOR2X1 U74677 ( .A(n71844), .B(n71843), .Y(n71846) );
  XNOR2X1 U74678 ( .A(n71846), .B(n71845), .Y(n71852) );
  NAND2X1 U74679 ( .A(n71847), .B(n72364), .Y(n71849) );
  NAND2X1 U74680 ( .A(n71849), .B(n71848), .Y(n71850) );
  XNOR2X1 U74681 ( .A(n71850), .B(n72367), .Y(n71851) );
  XNOR2X1 U74682 ( .A(n71852), .B(n71851), .Y(n72374) );
  INVX1 U74683 ( .A(n72308), .Y(n72311) );
  XNOR2X1 U74684 ( .A(n71853), .B(n41520), .Y(n72398) );
  XNOR2X1 U74685 ( .A(n72398), .B(n72397), .Y(n71854) );
  XNOR2X1 U74686 ( .A(n72401), .B(n71854), .Y(n72295) );
  XNOR2X1 U74687 ( .A(n72295), .B(n72327), .Y(n71859) );
  NAND2X1 U74688 ( .A(n71856), .B(n71855), .Y(n71858) );
  NAND2X1 U74689 ( .A(n71858), .B(n71857), .Y(n72298) );
  XNOR2X1 U74690 ( .A(n72289), .B(n72291), .Y(n71864) );
  NAND2X1 U74691 ( .A(n72327), .B(n71860), .Y(n71863) );
  NAND2X1 U74692 ( .A(n72327), .B(n71861), .Y(n71862) );
  XNOR2X1 U74693 ( .A(n71864), .B(n41720), .Y(n72282) );
  XNOR2X1 U74694 ( .A(n72282), .B(n72283), .Y(n71870) );
  INVX1 U74695 ( .A(n71865), .Y(n71866) );
  NOR2X1 U74696 ( .A(n71866), .B(n72288), .Y(n71869) );
  NOR2X1 U74697 ( .A(n71867), .B(n72288), .Y(n71868) );
  NOR2X1 U74698 ( .A(n71869), .B(n71868), .Y(n72285) );
  XNOR2X1 U74699 ( .A(n71870), .B(n72285), .Y(n72275) );
  XNOR2X1 U74700 ( .A(n72275), .B(n72326), .Y(n71875) );
  NAND2X1 U74701 ( .A(n72283), .B(n71871), .Y(n71874) );
  NAND2X1 U74702 ( .A(n72283), .B(n71872), .Y(n71873) );
  XNOR2X1 U74703 ( .A(n71875), .B(n41721), .Y(n72267) );
  XNOR2X1 U74704 ( .A(n72267), .B(n72355), .Y(n71880) );
  NAND2X1 U74705 ( .A(n72326), .B(n71876), .Y(n71879) );
  NAND2X1 U74706 ( .A(n72326), .B(n71877), .Y(n71878) );
  NAND2X1 U74707 ( .A(n71879), .B(n71878), .Y(n72270) );
  XNOR2X1 U74708 ( .A(n72261), .B(n72263), .Y(n71884) );
  NAND2X1 U74709 ( .A(n72355), .B(n71881), .Y(n71883) );
  XNOR2X1 U74710 ( .A(n71884), .B(n41723), .Y(n72423) );
  NAND2X1 U74711 ( .A(n72422), .B(n71885), .Y(n71887) );
  NAND2X1 U74712 ( .A(n71887), .B(n71310), .Y(n72420) );
  XNOR2X1 U74713 ( .A(n72420), .B(n72425), .Y(n71888) );
  XNOR2X1 U74714 ( .A(n72423), .B(n71888), .Y(n71892) );
  NAND2X1 U74715 ( .A(n72263), .B(n41512), .Y(n71890) );
  NAND2X1 U74716 ( .A(n71890), .B(n70997), .Y(n72421) );
  XNOR2X1 U74717 ( .A(n72421), .B(n72422), .Y(n71891) );
  XNOR2X1 U74718 ( .A(n71892), .B(n71891), .Y(n72438) );
  XNOR2X1 U74719 ( .A(n72438), .B(n72439), .Y(n71896) );
  NAND2X1 U74720 ( .A(n41511), .B(n71893), .Y(n71895) );
  NAND2X1 U74721 ( .A(n71895), .B(n71894), .Y(n72436) );
  NAND2X1 U74722 ( .A(n72447), .B(n71897), .Y(n72446) );
  XNOR2X1 U74723 ( .A(n72446), .B(n72456), .Y(n71898) );
  XNOR2X1 U74724 ( .A(n72448), .B(n71898), .Y(n71903) );
  NAND2X1 U74725 ( .A(n72439), .B(n41516), .Y(n71901) );
  NAND2X1 U74726 ( .A(n72439), .B(n71899), .Y(n71900) );
  NAND2X1 U74727 ( .A(n71901), .B(n71900), .Y(n72252) );
  XNOR2X1 U74728 ( .A(n72252), .B(n72447), .Y(n71902) );
  XNOR2X1 U74729 ( .A(n71903), .B(n71902), .Y(n72462) );
  INVX1 U74730 ( .A(n72462), .Y(n72465) );
  XNOR2X1 U74731 ( .A(n72464), .B(n72465), .Y(n71908) );
  NAND2X1 U74732 ( .A(n72456), .B(n71904), .Y(n71907) );
  NAND2X1 U74733 ( .A(n72456), .B(n71905), .Y(n71906) );
  XNOR2X1 U74734 ( .A(n71908), .B(n41717), .Y(n72248) );
  XNOR2X1 U74735 ( .A(n71922), .B(n71923), .Y(n71911) );
  XNOR2X1 U74736 ( .A(n41710), .B(n71911), .Y(n71914) );
  INVX1 U74737 ( .A(n71914), .Y(n71913) );
  NAND2X1 U74738 ( .A(n71913), .B(n71912), .Y(n71918) );
  NAND2X1 U74739 ( .A(n71915), .B(n71914), .Y(n71916) );
  NAND2X1 U74740 ( .A(n41737), .B(n71916), .Y(n71917) );
  NAND2X1 U74741 ( .A(n71918), .B(n71917), .Y(n72472) );
  NAND2X1 U74742 ( .A(n43614), .B(n39844), .Y(n72480) );
  INVX1 U74743 ( .A(n72480), .Y(n72477) );
  XNOR2X1 U74744 ( .A(n72472), .B(n72477), .Y(n71919) );
  XNOR2X1 U74745 ( .A(n72248), .B(n71919), .Y(n71928) );
  INVX1 U74746 ( .A(n71922), .Y(n71921) );
  NAND2X1 U74747 ( .A(n71921), .B(n71920), .Y(n71926) );
  NAND2X1 U74748 ( .A(n71923), .B(n71922), .Y(n71924) );
  NAND2X1 U74749 ( .A(n41710), .B(n71924), .Y(n71925) );
  NAND2X1 U74750 ( .A(n71926), .B(n71925), .Y(n72473) );
  NAND2X1 U74751 ( .A(n44054), .B(n43607), .Y(n72475) );
  INVX1 U74752 ( .A(n72475), .Y(n72337) );
  XNOR2X1 U74753 ( .A(n72473), .B(n72337), .Y(n71927) );
  XNOR2X1 U74754 ( .A(n71928), .B(n71927), .Y(n72488) );
  XNOR2X1 U74755 ( .A(n72488), .B(n72486), .Y(n71935) );
  NAND2X1 U74756 ( .A(n72486), .B(n71929), .Y(n71934) );
  NAND2X1 U74757 ( .A(n72489), .B(n71930), .Y(n71932) );
  NAND2X1 U74758 ( .A(n71932), .B(n71931), .Y(n71933) );
  XNOR2X1 U74759 ( .A(n71935), .B(n41712), .Y(n72242) );
  XNOR2X1 U74760 ( .A(n41706), .B(n71936), .Y(n71947) );
  XNOR2X1 U74761 ( .A(n71947), .B(n72347), .Y(n71937) );
  XNOR2X1 U74762 ( .A(n71938), .B(n71937), .Y(n71939) );
  NAND2X1 U74763 ( .A(n72317), .B(n71939), .Y(n71944) );
  INVX1 U74764 ( .A(n71939), .Y(n71940) );
  NAND2X1 U74765 ( .A(n71940), .B(n72233), .Y(n71942) );
  NAND2X1 U74766 ( .A(n71942), .B(n71941), .Y(n71943) );
  NAND2X1 U74767 ( .A(n71944), .B(n71943), .Y(n72235) );
  XNOR2X1 U74768 ( .A(n72235), .B(n72317), .Y(n71945) );
  XNOR2X1 U74769 ( .A(n72242), .B(n71945), .Y(n71953) );
  INVX1 U74770 ( .A(n71947), .Y(n71946) );
  NAND2X1 U74771 ( .A(n72347), .B(n71946), .Y(n71951) );
  NAND2X1 U74772 ( .A(n71947), .B(n72241), .Y(n71949) );
  NAND2X1 U74773 ( .A(n71949), .B(n71948), .Y(n71950) );
  NAND2X1 U74774 ( .A(n71951), .B(n71950), .Y(n72231) );
  XNOR2X1 U74775 ( .A(n72231), .B(n72347), .Y(n71952) );
  XNOR2X1 U74776 ( .A(n71953), .B(n71952), .Y(n72226) );
  XNOR2X1 U74777 ( .A(n72226), .B(n72318), .Y(n71960) );
  NAND2X1 U74778 ( .A(n72318), .B(n71954), .Y(n71959) );
  NAND2X1 U74779 ( .A(n71955), .B(n72225), .Y(n71957) );
  NAND2X1 U74780 ( .A(n71957), .B(n71956), .Y(n71958) );
  XNOR2X1 U74781 ( .A(n71960), .B(n41699), .Y(n72218) );
  XNOR2X1 U74782 ( .A(n41687), .B(n71961), .Y(n71970) );
  XNOR2X1 U74783 ( .A(n71970), .B(n72217), .Y(n71962) );
  XNOR2X1 U74784 ( .A(n71963), .B(n71962), .Y(n71965) );
  INVX1 U74785 ( .A(n71965), .Y(n71964) );
  NAND2X1 U74786 ( .A(n72212), .B(n71964), .Y(n71968) );
  NAND2X1 U74787 ( .A(n71965), .B(n72208), .Y(n71966) );
  NAND2X1 U74788 ( .A(n71966), .B(n71979), .Y(n71967) );
  NAND2X1 U74789 ( .A(n71968), .B(n71967), .Y(n72209) );
  XNOR2X1 U74790 ( .A(n72209), .B(n72212), .Y(n71969) );
  XNOR2X1 U74791 ( .A(n72218), .B(n71969), .Y(n71977) );
  NAND2X1 U74792 ( .A(n72217), .B(n71970), .Y(n71975) );
  INVX1 U74793 ( .A(n71970), .Y(n71971) );
  NAND2X1 U74794 ( .A(n71971), .B(n72219), .Y(n71973) );
  NAND2X1 U74795 ( .A(n71973), .B(n71972), .Y(n71974) );
  NAND2X1 U74796 ( .A(n71975), .B(n71974), .Y(n72221) );
  XNOR2X1 U74797 ( .A(n72221), .B(n72217), .Y(n71976) );
  XNOR2X1 U74798 ( .A(n71977), .B(n71976), .Y(n72201) );
  XNOR2X1 U74799 ( .A(n72201), .B(n72200), .Y(n71986) );
  NAND2X1 U74800 ( .A(n72200), .B(n71980), .Y(n71985) );
  INVX1 U74801 ( .A(n71980), .Y(n71981) );
  NAND2X1 U74802 ( .A(n71981), .B(n72202), .Y(n71983) );
  NAND2X1 U74803 ( .A(n71983), .B(n71982), .Y(n71984) );
  NAND2X1 U74804 ( .A(n71985), .B(n71984), .Y(n72204) );
  INVX1 U74805 ( .A(n72520), .Y(n72523) );
  XNOR2X1 U74806 ( .A(n72512), .B(n72523), .Y(n71987) );
  XNOR2X1 U74807 ( .A(n71988), .B(n71987), .Y(n71994) );
  NAND2X1 U74808 ( .A(n42187), .B(n71989), .Y(n71993) );
  NAND2X1 U74809 ( .A(n71990), .B(n42999), .Y(n71991) );
  NAND2X1 U74810 ( .A(n71991), .B(n71998), .Y(n71992) );
  NAND2X1 U74811 ( .A(n71993), .B(n71992), .Y(n72521) );
  XNOR2X1 U74812 ( .A(n71995), .B(n42187), .Y(n72000) );
  XNOR2X1 U74813 ( .A(n72000), .B(n71999), .Y(n72010) );
  INVX1 U74814 ( .A(n72010), .Y(n72011) );
  XNOR2X1 U74815 ( .A(n43602), .B(n72011), .Y(n72005) );
  INVX1 U74816 ( .A(n72005), .Y(n72001) );
  NAND2X1 U74817 ( .A(n72001), .B(n40683), .Y(n72003) );
  NAND2X1 U74818 ( .A(n72003), .B(n72002), .Y(n72008) );
  XNOR2X1 U74819 ( .A(n72005), .B(n72004), .Y(n72006) );
  NAND2X1 U74820 ( .A(n43615), .B(n72006), .Y(n72007) );
  NAND2X1 U74821 ( .A(n72008), .B(n72007), .Y(n72530) );
  XNOR2X1 U74822 ( .A(n72530), .B(n43616), .Y(n72009) );
  XNOR2X1 U74823 ( .A(n72545), .B(n72009), .Y(n72028) );
  NAND2X1 U74824 ( .A(n43599), .B(n72010), .Y(n72015) );
  NAND2X1 U74825 ( .A(n72011), .B(n43597), .Y(n72013) );
  NAND2X1 U74826 ( .A(n72013), .B(n72012), .Y(n72014) );
  NAND2X1 U74827 ( .A(n72015), .B(n72014), .Y(n72192) );
  XNOR2X1 U74828 ( .A(n72192), .B(n43602), .Y(n72016) );
  XNOR2X1 U74829 ( .A(n43618), .B(n72016), .Y(n72026) );
  XNOR2X1 U74830 ( .A(n72018), .B(n72017), .Y(n72019) );
  NAND2X1 U74831 ( .A(n43617), .B(n72019), .Y(n72024) );
  INVX1 U74832 ( .A(n72019), .Y(n72020) );
  NAND2X1 U74833 ( .A(n72020), .B(n42995), .Y(n72022) );
  NAND2X1 U74834 ( .A(n72022), .B(n72021), .Y(n72023) );
  NAND2X1 U74835 ( .A(n72024), .B(n72023), .Y(n72543) );
  INVX1 U74836 ( .A(n72543), .Y(n72025) );
  XNOR2X1 U74837 ( .A(n72026), .B(n72025), .Y(n72027) );
  XNOR2X1 U74838 ( .A(n72028), .B(n72027), .Y(n72187) );
  INVX1 U74839 ( .A(n72187), .Y(n72186) );
  XNOR2X1 U74840 ( .A(n72163), .B(n72186), .Y(n72029) );
  XNOR2X1 U74841 ( .A(n72030), .B(n72029), .Y(n72038) );
  INVX1 U74842 ( .A(n72031), .Y(n72047) );
  XNOR2X1 U74843 ( .A(n72047), .B(n72032), .Y(n72034) );
  INVX1 U74844 ( .A(n72034), .Y(n72033) );
  NAND2X1 U74845 ( .A(n43581), .B(n72033), .Y(n72037) );
  NAND2X1 U74846 ( .A(n72034), .B(n43585), .Y(n72035) );
  NAND2X1 U74847 ( .A(n72035), .B(n72048), .Y(n72036) );
  XNOR2X1 U74848 ( .A(n72038), .B(n41238), .Y(n72177) );
  NAND2X1 U74849 ( .A(n41012), .B(n72040), .Y(n72044) );
  NAND2X1 U74850 ( .A(n72042), .B(n72041), .Y(n72043) );
  NAND2X1 U74851 ( .A(n72044), .B(n72043), .Y(n72159) );
  XNOR2X1 U74852 ( .A(n72045), .B(n72152), .Y(n72046) );
  XNOR2X1 U74853 ( .A(n72047), .B(n72046), .Y(n72049) );
  INVX1 U74854 ( .A(n72048), .Y(n72059) );
  XNOR2X1 U74855 ( .A(n72049), .B(n72059), .Y(n72050) );
  XNOR2X1 U74856 ( .A(n72051), .B(n72050), .Y(n72053) );
  INVX1 U74857 ( .A(n72053), .Y(n72052) );
  NAND2X1 U74858 ( .A(n43535), .B(n72052), .Y(n72057) );
  NAND2X1 U74859 ( .A(n72053), .B(n43539), .Y(n72055) );
  NAND2X1 U74860 ( .A(n72055), .B(n72054), .Y(n72056) );
  NAND2X1 U74861 ( .A(n72057), .B(n72056), .Y(n72146) );
  XNOR2X1 U74862 ( .A(n43580), .B(n72149), .Y(n72065) );
  NAND2X1 U74863 ( .A(n43577), .B(n72060), .Y(n72174) );
  NOR2X1 U74864 ( .A(n72065), .B(n72174), .Y(n72064) );
  NAND2X1 U74865 ( .A(n72062), .B(n72061), .Y(n72173) );
  NOR2X1 U74866 ( .A(n72064), .B(n72063), .Y(n72067) );
  OR2X1 U74867 ( .A(n72065), .B(n72173), .Y(n72066) );
  NAND2X1 U74868 ( .A(n72067), .B(n72066), .Y(n72068) );
  XOR2X1 U74869 ( .A(n72146), .B(n72068), .Y(n72069) );
  XOR2X1 U74870 ( .A(n72177), .B(n72070), .Y(n72595) );
  XNOR2X1 U74871 ( .A(n72079), .B(n38683), .Y(n72072) );
  INVX1 U74872 ( .A(n72072), .Y(n72559) );
  NAND2X1 U74873 ( .A(n72560), .B(n43623), .Y(n72071) );
  NOR2X1 U74874 ( .A(n72559), .B(n72071), .Y(n72074) );
  NAND2X1 U74875 ( .A(n43619), .B(n72072), .Y(n72562) );
  NOR2X1 U74876 ( .A(n72074), .B(n72073), .Y(n72075) );
  INVX1 U74877 ( .A(n72611), .Y(n72090) );
  XNOR2X1 U74878 ( .A(n72078), .B(n38683), .Y(n72081) );
  XNOR2X1 U74879 ( .A(n72560), .B(n72079), .Y(n72080) );
  NAND2X1 U74880 ( .A(n43631), .B(n72082), .Y(n72087) );
  INVX1 U74881 ( .A(n72082), .Y(n72083) );
  NAND2X1 U74882 ( .A(n72083), .B(n43635), .Y(n72085) );
  NAND2X1 U74883 ( .A(n72085), .B(n72084), .Y(n72086) );
  NAND2X1 U74884 ( .A(n72087), .B(n72086), .Y(n72610) );
  XNOR2X1 U74885 ( .A(n72610), .B(n72088), .Y(n72089) );
  XNOR2X1 U74886 ( .A(n72090), .B(n72089), .Y(n72091) );
  XNOR2X1 U74887 ( .A(n72092), .B(n72091), .Y(n72671) );
  XNOR2X1 U74888 ( .A(n72617), .B(n72671), .Y(n72621) );
  INVX1 U74889 ( .A(n72621), .Y(n72622) );
  XNOR2X1 U74890 ( .A(n72093), .B(n72622), .Y(n72094) );
  XNOR2X1 U74891 ( .A(n72095), .B(n72094), .Y(n72685) );
  INVX1 U74892 ( .A(n72685), .Y(n72692) );
  INVX1 U74893 ( .A(n72666), .Y(n72665) );
  NAND2X1 U74894 ( .A(n72099), .B(n72098), .Y(n72100) );
  INVX1 U74895 ( .A(n72646), .Y(n72657) );
  INVX1 U74896 ( .A(n72106), .Y(n72109) );
  NAND2X1 U74897 ( .A(n43707), .B(n72107), .Y(n72108) );
  NOR2X1 U74898 ( .A(n72109), .B(n72108), .Y(n72110) );
  NAND2X1 U74899 ( .A(n72111), .B(n41070), .Y(n72117) );
  XNOR2X1 U74900 ( .A(n72113), .B(n72112), .Y(n72114) );
  XOR2X1 U74901 ( .A(n42129), .B(n72114), .Y(n72115) );
  NAND2X1 U74902 ( .A(n43718), .B(n72115), .Y(n72116) );
  NAND2X1 U74903 ( .A(n72117), .B(n72116), .Y(n72121) );
  NAND2X1 U74904 ( .A(n40192), .B(n40456), .Y(n72122) );
  NAND2X1 U74905 ( .A(n72657), .B(n72732), .Y(n72118) );
  NOR2X1 U74906 ( .A(n38580), .B(n72118), .Y(n72119) );
  NAND2X1 U74907 ( .A(n40457), .B(n72732), .Y(n72125) );
  NAND2X1 U74908 ( .A(n41070), .B(n72719), .Y(n72123) );
  NAND2X1 U74909 ( .A(n72123), .B(n72122), .Y(n72124) );
  OR2X1 U74910 ( .A(n72125), .B(n72124), .Y(n72126) );
  NAND2X1 U74911 ( .A(u_muldiv_mult_result_q[30]), .B(n44631), .Y(n13855) );
  XNOR2X1 U74912 ( .A(n72128), .B(n72127), .Y(n72129) );
  XNOR2X1 U74913 ( .A(n72129), .B(n42130), .Y(n72130) );
  NAND2X1 U74914 ( .A(n43718), .B(n72130), .Y(n72713) );
  INVX1 U74915 ( .A(n72713), .Y(n72660) );
  NAND2X1 U74916 ( .A(n72131), .B(n43527), .Y(n72135) );
  NAND2X1 U74917 ( .A(n43521), .B(n72132), .Y(n72133) );
  NAND2X1 U74918 ( .A(n39412), .B(n72133), .Y(n72134) );
  AND2X1 U74919 ( .A(n72135), .B(n72134), .Y(n72674) );
  XNOR2X1 U74920 ( .A(n72621), .B(n43655), .Y(n72138) );
  XNOR2X1 U74921 ( .A(n41142), .B(n72138), .Y(n72142) );
  INVX1 U74922 ( .A(n72142), .Y(n72140) );
  NAND2X1 U74923 ( .A(n72140), .B(n43530), .Y(n72141) );
  NAND2X1 U74924 ( .A(n72674), .B(n72141), .Y(n72144) );
  NAND2X1 U74925 ( .A(n43522), .B(n72142), .Y(n72143) );
  NAND2X1 U74926 ( .A(n72144), .B(n72143), .Y(n72639) );
  INVX1 U74927 ( .A(n72177), .Y(n72172) );
  NAND2X1 U74928 ( .A(n72172), .B(n43539), .Y(n72148) );
  NAND2X1 U74929 ( .A(n72148), .B(n72147), .Y(n72150) );
  XNOR2X1 U74930 ( .A(n72150), .B(n72149), .Y(n72151) );
  XNOR2X1 U74931 ( .A(n72152), .B(n72151), .Y(n72157) );
  INVX1 U74932 ( .A(n72157), .Y(n72156) );
  NAND2X1 U74933 ( .A(n41241), .B(n72156), .Y(n72572) );
  INVX1 U74934 ( .A(n72595), .Y(n72592) );
  NAND2X1 U74935 ( .A(n72592), .B(n43549), .Y(n72155) );
  NAND2X1 U74936 ( .A(n41481), .B(n72156), .Y(n72576) );
  NAND2X1 U74937 ( .A(n72572), .B(n72576), .Y(n72571) );
  NOR2X1 U74938 ( .A(n41481), .B(n41241), .Y(n72158) );
  NAND2X1 U74939 ( .A(n72158), .B(n72157), .Y(n72575) );
  NAND2X1 U74940 ( .A(n41012), .B(n72177), .Y(n72162) );
  NAND2X1 U74941 ( .A(n72172), .B(n43559), .Y(n72160) );
  NAND2X1 U74942 ( .A(n72160), .B(n72159), .Y(n72161) );
  NAND2X1 U74943 ( .A(n72162), .B(n72161), .Y(n72557) );
  INVX1 U74944 ( .A(n72163), .Y(n72166) );
  XNOR2X1 U74945 ( .A(n72187), .B(n43594), .Y(n72164) );
  NOR2X1 U74946 ( .A(n43568), .B(n72167), .Y(n72165) );
  NOR2X1 U74947 ( .A(n72166), .B(n72165), .Y(n72171) );
  INVX1 U74948 ( .A(n72167), .Y(n72169) );
  NOR2X1 U74949 ( .A(n72169), .B(n40670), .Y(n72170) );
  NOR2X1 U74950 ( .A(n72171), .B(n72170), .Y(n72181) );
  NOR2X1 U74951 ( .A(n72172), .B(n43574), .Y(n72176) );
  NAND2X1 U74952 ( .A(n72174), .B(n72173), .Y(n72175) );
  NOR2X1 U74953 ( .A(n72176), .B(n72175), .Y(n72179) );
  NOR2X1 U74954 ( .A(n43578), .B(n72177), .Y(n72178) );
  NOR2X1 U74955 ( .A(n72179), .B(n72178), .Y(n72180) );
  XNOR2X1 U74956 ( .A(n72181), .B(n72180), .Y(n72555) );
  NAND2X1 U74957 ( .A(n72187), .B(n43585), .Y(n72185) );
  NAND2X1 U74958 ( .A(n43582), .B(n72186), .Y(n72183) );
  NAND2X1 U74959 ( .A(n41238), .B(n72183), .Y(n72184) );
  NAND2X1 U74960 ( .A(n72185), .B(n72184), .Y(n72553) );
  NAND2X1 U74961 ( .A(n43592), .B(n72186), .Y(n72191) );
  NAND2X1 U74962 ( .A(n72187), .B(n42994), .Y(n72189) );
  NAND2X1 U74963 ( .A(n72189), .B(n72188), .Y(n72190) );
  NAND2X1 U74964 ( .A(n72191), .B(n72190), .Y(n72551) );
  INVX1 U74965 ( .A(n72545), .Y(n72542) );
  NAND2X1 U74966 ( .A(n72542), .B(n43597), .Y(n72195) );
  INVX1 U74967 ( .A(n72192), .Y(n72532) );
  NAND2X1 U74968 ( .A(n43602), .B(n72545), .Y(n72193) );
  NAND2X1 U74969 ( .A(n72532), .B(n72193), .Y(n72194) );
  NAND2X1 U74970 ( .A(n72195), .B(n72194), .Y(n72529) );
  NAND2X1 U74971 ( .A(n72510), .B(n72523), .Y(n72199) );
  NAND2X1 U74972 ( .A(n72520), .B(n72196), .Y(n72197) );
  NAND2X1 U74973 ( .A(n72197), .B(n72509), .Y(n72198) );
  NAND2X1 U74974 ( .A(n72199), .B(n72198), .Y(n72508) );
  NAND2X1 U74975 ( .A(n72200), .B(n72201), .Y(n72207) );
  INVX1 U74976 ( .A(n72201), .Y(n72203) );
  NAND2X1 U74977 ( .A(n72203), .B(n72202), .Y(n72205) );
  NAND2X1 U74978 ( .A(n72205), .B(n72204), .Y(n72206) );
  NAND2X1 U74979 ( .A(n72207), .B(n72206), .Y(n72506) );
  NAND2X1 U74980 ( .A(n72210), .B(n72208), .Y(n72216) );
  INVX1 U74981 ( .A(n72209), .Y(n72214) );
  INVX1 U74982 ( .A(n72210), .Y(n72211) );
  NAND2X1 U74983 ( .A(n72212), .B(n72211), .Y(n72213) );
  NAND2X1 U74984 ( .A(n72214), .B(n72213), .Y(n72215) );
  NAND2X1 U74985 ( .A(n72216), .B(n72215), .Y(n72504) );
  NAND2X1 U74986 ( .A(n72217), .B(n72218), .Y(n72224) );
  INVX1 U74987 ( .A(n72218), .Y(n72220) );
  NAND2X1 U74988 ( .A(n72220), .B(n72219), .Y(n72222) );
  NAND2X1 U74989 ( .A(n72222), .B(n72221), .Y(n72223) );
  NAND2X1 U74990 ( .A(n72224), .B(n72223), .Y(n72502) );
  NAND2X1 U74991 ( .A(n72226), .B(n72225), .Y(n72230) );
  INVX1 U74992 ( .A(n72226), .Y(n72227) );
  NAND2X1 U74993 ( .A(n72318), .B(n72227), .Y(n72228) );
  NAND2X1 U74994 ( .A(n41699), .B(n72228), .Y(n72229) );
  NAND2X1 U74995 ( .A(n72230), .B(n72229), .Y(n72500) );
  INVX1 U74996 ( .A(n72231), .Y(n72245) );
  XNOR2X1 U74997 ( .A(n72242), .B(n72347), .Y(n72232) );
  XNOR2X1 U74998 ( .A(n72245), .B(n72232), .Y(n72236) );
  INVX1 U74999 ( .A(n72236), .Y(n72234) );
  NAND2X1 U75000 ( .A(n72234), .B(n72233), .Y(n72240) );
  INVX1 U75001 ( .A(n72235), .Y(n72238) );
  NAND2X1 U75002 ( .A(n72317), .B(n72236), .Y(n72237) );
  NAND2X1 U75003 ( .A(n72238), .B(n72237), .Y(n72239) );
  NAND2X1 U75004 ( .A(n72240), .B(n72239), .Y(n72498) );
  NAND2X1 U75005 ( .A(n72242), .B(n72241), .Y(n72247) );
  INVX1 U75006 ( .A(n72242), .Y(n72243) );
  NAND2X1 U75007 ( .A(n72347), .B(n72243), .Y(n72244) );
  NAND2X1 U75008 ( .A(n72245), .B(n72244), .Y(n72246) );
  NAND2X1 U75009 ( .A(n72247), .B(n72246), .Y(n72496) );
  NAND2X1 U75010 ( .A(n72248), .B(n72475), .Y(n72251) );
  INVX1 U75011 ( .A(n72248), .Y(n72474) );
  NAND2X1 U75012 ( .A(n72337), .B(n72474), .Y(n72249) );
  NAND2X1 U75013 ( .A(n72249), .B(n72473), .Y(n72250) );
  NAND2X1 U75014 ( .A(n72251), .B(n72250), .Y(n72471) );
  NAND2X1 U75015 ( .A(n72448), .B(n72323), .Y(n72256) );
  INVX1 U75016 ( .A(n72252), .Y(n72450) );
  INVX1 U75017 ( .A(n72448), .Y(n72253) );
  NAND2X1 U75018 ( .A(n72447), .B(n72253), .Y(n72254) );
  NAND2X1 U75019 ( .A(n72450), .B(n72254), .Y(n72255) );
  NAND2X1 U75020 ( .A(n72256), .B(n72255), .Y(n72445) );
  NAND2X1 U75021 ( .A(n72422), .B(n72423), .Y(n72260) );
  INVX1 U75022 ( .A(n72423), .Y(n72257) );
  NAND2X1 U75023 ( .A(n72257), .B(n72356), .Y(n72258) );
  NAND2X1 U75024 ( .A(n72258), .B(n72421), .Y(n72259) );
  NAND2X1 U75025 ( .A(n72260), .B(n72259), .Y(n72419) );
  NAND2X1 U75026 ( .A(n72261), .B(n72328), .Y(n72266) );
  INVX1 U75027 ( .A(n72261), .Y(n72262) );
  NAND2X1 U75028 ( .A(n72263), .B(n72262), .Y(n72264) );
  NAND2X1 U75029 ( .A(n41723), .B(n72264), .Y(n72265) );
  NAND2X1 U75030 ( .A(n72266), .B(n72265), .Y(n72417) );
  NAND2X1 U75031 ( .A(n72355), .B(n72267), .Y(n72273) );
  INVX1 U75032 ( .A(n72267), .Y(n72269) );
  NAND2X1 U75033 ( .A(n72269), .B(n72268), .Y(n72271) );
  NAND2X1 U75034 ( .A(n72271), .B(n72270), .Y(n72272) );
  NAND2X1 U75035 ( .A(n72273), .B(n72272), .Y(n72415) );
  NAND2X1 U75036 ( .A(n72275), .B(n72274), .Y(n72279) );
  INVX1 U75037 ( .A(n72275), .Y(n72276) );
  NAND2X1 U75038 ( .A(n72326), .B(n72276), .Y(n72277) );
  NAND2X1 U75039 ( .A(n41721), .B(n72277), .Y(n72278) );
  NAND2X1 U75040 ( .A(n72279), .B(n72278), .Y(n72413) );
  INVX1 U75041 ( .A(n72282), .Y(n72281) );
  NAND2X1 U75042 ( .A(n72281), .B(n72280), .Y(n72287) );
  NAND2X1 U75043 ( .A(n72283), .B(n72282), .Y(n72284) );
  NAND2X1 U75044 ( .A(n72285), .B(n72284), .Y(n72286) );
  NAND2X1 U75045 ( .A(n72287), .B(n72286), .Y(n72411) );
  NAND2X1 U75046 ( .A(n72289), .B(n72288), .Y(n72294) );
  INVX1 U75047 ( .A(n72289), .Y(n72290) );
  NAND2X1 U75048 ( .A(n72291), .B(n72290), .Y(n72292) );
  NAND2X1 U75049 ( .A(n41720), .B(n72292), .Y(n72293) );
  NAND2X1 U75050 ( .A(n72294), .B(n72293), .Y(n72409) );
  NAND2X1 U75051 ( .A(n72327), .B(n72295), .Y(n72301) );
  INVX1 U75052 ( .A(n72295), .Y(n72297) );
  NAND2X1 U75053 ( .A(n72297), .B(n72296), .Y(n72299) );
  NAND2X1 U75054 ( .A(n72299), .B(n72298), .Y(n72300) );
  NAND2X1 U75055 ( .A(n72301), .B(n72300), .Y(n72407) );
  NOR2X1 U75056 ( .A(n72303), .B(n72302), .Y(n72307) );
  INVX1 U75057 ( .A(n72304), .Y(n72305) );
  NOR2X1 U75058 ( .A(n72305), .B(n41520), .Y(n72306) );
  NOR2X1 U75059 ( .A(n72307), .B(n72306), .Y(n72395) );
  NAND2X1 U75060 ( .A(n72333), .B(n72308), .Y(n72315) );
  INVX1 U75061 ( .A(n72309), .Y(n72313) );
  NAND2X1 U75062 ( .A(n72311), .B(n72310), .Y(n72312) );
  NAND2X1 U75063 ( .A(n72313), .B(n72312), .Y(n72314) );
  NAND2X1 U75064 ( .A(n72315), .B(n72314), .Y(n72393) );
  XNOR2X1 U75065 ( .A(n72316), .B(n41734), .Y(n72322) );
  XNOR2X1 U75066 ( .A(n72318), .B(n72317), .Y(n72320) );
  XNOR2X1 U75067 ( .A(n72320), .B(n72319), .Y(n72321) );
  XNOR2X1 U75068 ( .A(n72322), .B(n72321), .Y(n72346) );
  XNOR2X1 U75069 ( .A(n72425), .B(n72439), .Y(n72325) );
  XNOR2X1 U75070 ( .A(n72323), .B(n72370), .Y(n72324) );
  XNOR2X1 U75071 ( .A(n72325), .B(n72324), .Y(n72332) );
  XNOR2X1 U75072 ( .A(n72397), .B(n72326), .Y(n72330) );
  XNOR2X1 U75073 ( .A(n72328), .B(n72327), .Y(n72329) );
  XNOR2X1 U75074 ( .A(n72330), .B(n72329), .Y(n72331) );
  XNOR2X1 U75075 ( .A(n72332), .B(n72331), .Y(n72344) );
  XNOR2X1 U75076 ( .A(n72334), .B(n72333), .Y(n72335) );
  XNOR2X1 U75077 ( .A(n43599), .B(n72335), .Y(n72342) );
  XNOR2X1 U75078 ( .A(n72387), .B(n72456), .Y(n72340) );
  NAND2X1 U75079 ( .A(n72337), .B(n43604), .Y(n72338) );
  INVX1 U75080 ( .A(n72464), .Y(n72461) );
  XNOR2X1 U75081 ( .A(n72338), .B(n72461), .Y(n72339) );
  XNOR2X1 U75082 ( .A(n72340), .B(n72339), .Y(n72341) );
  XNOR2X1 U75083 ( .A(n72342), .B(n72341), .Y(n72343) );
  XNOR2X1 U75084 ( .A(n72344), .B(n72343), .Y(n72345) );
  XNOR2X1 U75085 ( .A(n72346), .B(n72345), .Y(n72363) );
  XNOR2X1 U75086 ( .A(n72347), .B(n72486), .Y(n72351) );
  NAND2X1 U75087 ( .A(n43614), .B(n43607), .Y(n72349) );
  XNOR2X1 U75088 ( .A(n72349), .B(n72477), .Y(n72350) );
  XNOR2X1 U75089 ( .A(n72351), .B(n72350), .Y(n72352) );
  XNOR2X1 U75090 ( .A(n72353), .B(n72352), .Y(n72361) );
  XNOR2X1 U75091 ( .A(n72356), .B(n72355), .Y(n72357) );
  XNOR2X1 U75092 ( .A(n72359), .B(n72358), .Y(n72360) );
  XNOR2X1 U75093 ( .A(n72361), .B(n72360), .Y(n72362) );
  XNOR2X1 U75094 ( .A(n72363), .B(n72362), .Y(n72381) );
  NAND2X1 U75095 ( .A(n72365), .B(n72364), .Y(n72369) );
  NAND2X1 U75096 ( .A(n72367), .B(n72366), .Y(n72368) );
  NOR2X1 U75097 ( .A(n72369), .B(n72368), .Y(n72379) );
  NAND2X1 U75098 ( .A(n72371), .B(n72370), .Y(n72377) );
  NAND2X1 U75099 ( .A(n72373), .B(n72372), .Y(n72375) );
  NAND2X1 U75100 ( .A(n72375), .B(n72374), .Y(n72376) );
  NAND2X1 U75101 ( .A(n72377), .B(n72376), .Y(n72378) );
  NOR2X1 U75102 ( .A(n72379), .B(n72378), .Y(n72380) );
  XNOR2X1 U75103 ( .A(n72381), .B(n72380), .Y(n72391) );
  NOR2X1 U75104 ( .A(n72383), .B(n72382), .Y(n72385) );
  NOR2X1 U75105 ( .A(n72385), .B(n72384), .Y(n72389) );
  NOR2X1 U75106 ( .A(n72387), .B(n72386), .Y(n72388) );
  NOR2X1 U75107 ( .A(n72389), .B(n72388), .Y(n72390) );
  XNOR2X1 U75108 ( .A(n72391), .B(n72390), .Y(n72392) );
  XNOR2X1 U75109 ( .A(n72393), .B(n72392), .Y(n72394) );
  XNOR2X1 U75110 ( .A(n72395), .B(n72394), .Y(n72405) );
  NOR2X1 U75111 ( .A(n72397), .B(n72396), .Y(n72399) );
  NOR2X1 U75112 ( .A(n72399), .B(n72398), .Y(n72403) );
  NOR2X1 U75113 ( .A(n72401), .B(n72400), .Y(n72402) );
  NOR2X1 U75114 ( .A(n72403), .B(n72402), .Y(n72404) );
  XNOR2X1 U75115 ( .A(n72405), .B(n72404), .Y(n72406) );
  XNOR2X1 U75116 ( .A(n72407), .B(n72406), .Y(n72408) );
  XNOR2X1 U75117 ( .A(n72409), .B(n72408), .Y(n72410) );
  XNOR2X1 U75118 ( .A(n72411), .B(n72410), .Y(n72412) );
  XNOR2X1 U75119 ( .A(n72413), .B(n72412), .Y(n72414) );
  XNOR2X1 U75120 ( .A(n72415), .B(n72414), .Y(n72416) );
  XNOR2X1 U75121 ( .A(n72417), .B(n72416), .Y(n72418) );
  XNOR2X1 U75122 ( .A(n72419), .B(n72418), .Y(n72433) );
  INVX1 U75123 ( .A(n72420), .Y(n72427) );
  INVX1 U75124 ( .A(n72429), .Y(n72424) );
  NOR2X1 U75125 ( .A(n72425), .B(n72424), .Y(n72426) );
  NOR2X1 U75126 ( .A(n72427), .B(n72426), .Y(n72431) );
  NOR2X1 U75127 ( .A(n72429), .B(n72428), .Y(n72430) );
  NOR2X1 U75128 ( .A(n72431), .B(n72430), .Y(n72432) );
  XNOR2X1 U75129 ( .A(n72433), .B(n72432), .Y(n72443) );
  INVX1 U75130 ( .A(n72438), .Y(n72435) );
  NOR2X1 U75131 ( .A(n72435), .B(n72434), .Y(n72437) );
  NOR2X1 U75132 ( .A(n72437), .B(n72436), .Y(n72441) );
  NOR2X1 U75133 ( .A(n72439), .B(n72438), .Y(n72440) );
  NOR2X1 U75134 ( .A(n72441), .B(n72440), .Y(n72442) );
  XNOR2X1 U75135 ( .A(n72443), .B(n72442), .Y(n72444) );
  XNOR2X1 U75136 ( .A(n72445), .B(n72444), .Y(n72460) );
  INVX1 U75137 ( .A(n72446), .Y(n72454) );
  XNOR2X1 U75138 ( .A(n72448), .B(n72447), .Y(n72449) );
  XNOR2X1 U75139 ( .A(n72450), .B(n72449), .Y(n72455) );
  INVX1 U75140 ( .A(n72455), .Y(n72452) );
  NOR2X1 U75141 ( .A(n72452), .B(n72451), .Y(n72453) );
  NOR2X1 U75142 ( .A(n72454), .B(n72453), .Y(n72458) );
  NOR2X1 U75143 ( .A(n72456), .B(n72455), .Y(n72457) );
  NOR2X1 U75144 ( .A(n72458), .B(n72457), .Y(n72459) );
  XNOR2X1 U75145 ( .A(n72460), .B(n72459), .Y(n72469) );
  NOR2X1 U75146 ( .A(n72462), .B(n72461), .Y(n72463) );
  NOR2X1 U75147 ( .A(n41717), .B(n72463), .Y(n72467) );
  NOR2X1 U75148 ( .A(n72465), .B(n72464), .Y(n72466) );
  NOR2X1 U75149 ( .A(n72467), .B(n72466), .Y(n72468) );
  XNOR2X1 U75150 ( .A(n72469), .B(n72468), .Y(n72470) );
  XNOR2X1 U75151 ( .A(n72471), .B(n72470), .Y(n72485) );
  INVX1 U75152 ( .A(n72472), .Y(n72479) );
  INVX1 U75153 ( .A(n72481), .Y(n72476) );
  NOR2X1 U75154 ( .A(n72477), .B(n72476), .Y(n72478) );
  NOR2X1 U75155 ( .A(n72479), .B(n72478), .Y(n72483) );
  NOR2X1 U75156 ( .A(n72481), .B(n72480), .Y(n72482) );
  NOR2X1 U75157 ( .A(n72483), .B(n72482), .Y(n72484) );
  XNOR2X1 U75158 ( .A(n72485), .B(n72484), .Y(n72494) );
  NOR2X1 U75159 ( .A(n72486), .B(n72488), .Y(n72487) );
  NOR2X1 U75160 ( .A(n41712), .B(n72487), .Y(n72492) );
  INVX1 U75161 ( .A(n72488), .Y(n72490) );
  NOR2X1 U75162 ( .A(n72490), .B(n72489), .Y(n72491) );
  NOR2X1 U75163 ( .A(n72492), .B(n72491), .Y(n72493) );
  XNOR2X1 U75164 ( .A(n72494), .B(n72493), .Y(n72495) );
  XNOR2X1 U75165 ( .A(n72496), .B(n72495), .Y(n72497) );
  XNOR2X1 U75166 ( .A(n72498), .B(n72497), .Y(n72499) );
  XNOR2X1 U75167 ( .A(n72500), .B(n72499), .Y(n72501) );
  XNOR2X1 U75168 ( .A(n72502), .B(n72501), .Y(n72503) );
  XNOR2X1 U75169 ( .A(n72504), .B(n72503), .Y(n72505) );
  XNOR2X1 U75170 ( .A(n72506), .B(n72505), .Y(n72507) );
  XNOR2X1 U75171 ( .A(n72508), .B(n72507), .Y(n72519) );
  INVX1 U75172 ( .A(n72514), .Y(n72511) );
  NOR2X1 U75173 ( .A(n72511), .B(n43000), .Y(n72513) );
  NOR2X1 U75174 ( .A(n72513), .B(n72512), .Y(n72517) );
  NOR2X1 U75175 ( .A(n72515), .B(n72514), .Y(n72516) );
  NOR2X1 U75176 ( .A(n72517), .B(n72516), .Y(n72518) );
  XNOR2X1 U75177 ( .A(n72519), .B(n72518), .Y(n72527) );
  NOR2X1 U75178 ( .A(n72520), .B(n42998), .Y(n72522) );
  NOR2X1 U75179 ( .A(n72522), .B(n72521), .Y(n72525) );
  NOR2X1 U75180 ( .A(n42187), .B(n72523), .Y(n72524) );
  NOR2X1 U75181 ( .A(n72525), .B(n72524), .Y(n72526) );
  XNOR2X1 U75182 ( .A(n72527), .B(n72526), .Y(n72528) );
  XNOR2X1 U75183 ( .A(n72529), .B(n72528), .Y(n72541) );
  INVX1 U75184 ( .A(n72530), .Y(n72535) );
  XNOR2X1 U75185 ( .A(n72545), .B(n43602), .Y(n72531) );
  XNOR2X1 U75186 ( .A(n72532), .B(n72531), .Y(n72537) );
  INVX1 U75187 ( .A(n72537), .Y(n72533) );
  NOR2X1 U75188 ( .A(n43616), .B(n72533), .Y(n72534) );
  NOR2X1 U75189 ( .A(n72535), .B(n72534), .Y(n72539) );
  NOR2X1 U75190 ( .A(n72537), .B(n40683), .Y(n72538) );
  NOR2X1 U75191 ( .A(n72539), .B(n72538), .Y(n72540) );
  XNOR2X1 U75192 ( .A(n72541), .B(n72540), .Y(n72549) );
  NOR2X1 U75193 ( .A(n72542), .B(n42997), .Y(n72544) );
  NOR2X1 U75194 ( .A(n72544), .B(n72543), .Y(n72547) );
  NOR2X1 U75195 ( .A(n43617), .B(n72545), .Y(n72546) );
  NOR2X1 U75196 ( .A(n72547), .B(n72546), .Y(n72548) );
  XNOR2X1 U75197 ( .A(n72549), .B(n72548), .Y(n72550) );
  XNOR2X1 U75198 ( .A(n72551), .B(n72550), .Y(n72552) );
  XNOR2X1 U75199 ( .A(n72553), .B(n72552), .Y(n72554) );
  XNOR2X1 U75200 ( .A(n72555), .B(n72554), .Y(n72556) );
  XNOR2X1 U75201 ( .A(n72557), .B(n72556), .Y(n72569) );
  NOR2X1 U75202 ( .A(n72592), .B(n43628), .Y(n72565) );
  NAND2X1 U75203 ( .A(n72559), .B(n43624), .Y(n72561) );
  NAND2X1 U75204 ( .A(n72561), .B(n72560), .Y(n72563) );
  NAND2X1 U75205 ( .A(n72563), .B(n72562), .Y(n72564) );
  NOR2X1 U75206 ( .A(n72565), .B(n72564), .Y(n72567) );
  NOR2X1 U75207 ( .A(n43620), .B(n72595), .Y(n72566) );
  NOR2X1 U75208 ( .A(n72567), .B(n72566), .Y(n72568) );
  XNOR2X1 U75209 ( .A(n72569), .B(n72568), .Y(n72577) );
  NAND2X1 U75210 ( .A(n72575), .B(n72577), .Y(n72570) );
  NOR2X1 U75211 ( .A(n72571), .B(n72570), .Y(n72574) );
  NOR2X1 U75212 ( .A(n72577), .B(n72572), .Y(n72573) );
  NOR2X1 U75213 ( .A(n72574), .B(n72573), .Y(n72581) );
  NOR2X1 U75214 ( .A(n72577), .B(n72575), .Y(n72579) );
  NOR2X1 U75215 ( .A(n72577), .B(n72576), .Y(n72578) );
  NOR2X1 U75216 ( .A(n72579), .B(n72578), .Y(n72580) );
  NAND2X1 U75217 ( .A(n72581), .B(n72580), .Y(n72604) );
  XNOR2X1 U75218 ( .A(n43673), .B(n43707), .Y(n72582) );
  XNOR2X1 U75219 ( .A(n43644), .B(n72582), .Y(n72585) );
  XNOR2X1 U75220 ( .A(n72583), .B(n43692), .Y(n72584) );
  XNOR2X1 U75221 ( .A(n72585), .B(n72584), .Y(n72590) );
  INVX1 U75222 ( .A(n72586), .Y(n72668) );
  XNOR2X1 U75223 ( .A(n43621), .B(n72668), .Y(n72588) );
  XNOR2X1 U75224 ( .A(n72588), .B(n72587), .Y(n72589) );
  XNOR2X1 U75225 ( .A(n72590), .B(n72589), .Y(n72594) );
  NAND2X1 U75226 ( .A(n72592), .B(n43637), .Y(n72593) );
  NAND2X1 U75227 ( .A(n72593), .B(n72610), .Y(n72596) );
  NOR2X1 U75228 ( .A(n72594), .B(n72596), .Y(n72602) );
  INVX1 U75229 ( .A(n72594), .Y(n72598) );
  NOR2X1 U75230 ( .A(n72598), .B(n41489), .Y(n72597) );
  NAND2X1 U75231 ( .A(n72597), .B(n72596), .Y(n72600) );
  NAND2X1 U75232 ( .A(n41489), .B(n72598), .Y(n72599) );
  NAND2X1 U75233 ( .A(n72600), .B(n72599), .Y(n72601) );
  NOR2X1 U75234 ( .A(n72602), .B(n72601), .Y(n72603) );
  XNOR2X1 U75235 ( .A(n72604), .B(n72603), .Y(n72638) );
  NAND2X1 U75236 ( .A(n72605), .B(n38555), .Y(n72607) );
  NAND2X1 U75237 ( .A(n72607), .B(n72606), .Y(n72609) );
  NAND2X1 U75238 ( .A(n72609), .B(n72608), .Y(n72627) );
  XNOR2X1 U75239 ( .A(n72629), .B(n43666), .Y(n72612) );
  INVX1 U75240 ( .A(n72615), .Y(n72614) );
  NAND2X1 U75241 ( .A(n72614), .B(n39301), .Y(n72619) );
  NAND2X1 U75242 ( .A(n40142), .B(n72615), .Y(n72616) );
  NAND2X1 U75243 ( .A(n72617), .B(n72616), .Y(n72618) );
  NAND2X1 U75244 ( .A(n72619), .B(n72618), .Y(n72636) );
  NAND2X1 U75245 ( .A(n72621), .B(n43656), .Y(n72625) );
  NAND2X1 U75246 ( .A(n43653), .B(n72622), .Y(n72623) );
  NAND2X1 U75247 ( .A(n41142), .B(n72623), .Y(n72624) );
  NAND2X1 U75248 ( .A(n72625), .B(n72624), .Y(n72634) );
  NOR2X1 U75249 ( .A(n72629), .B(n43672), .Y(n72628) );
  NOR2X1 U75250 ( .A(n72628), .B(n72627), .Y(n72632) );
  INVX1 U75251 ( .A(n72629), .Y(n72630) );
  NOR2X1 U75252 ( .A(n43666), .B(n72630), .Y(n72631) );
  NOR2X1 U75253 ( .A(n72632), .B(n72631), .Y(n72633) );
  XNOR2X1 U75254 ( .A(n72634), .B(n72633), .Y(n72635) );
  XNOR2X1 U75255 ( .A(n72636), .B(n72635), .Y(n72637) );
  XNOR2X1 U75256 ( .A(n72638), .B(n72637), .Y(n72640) );
  NAND2X1 U75257 ( .A(n72639), .B(n72640), .Y(n72642) );
  OR2X1 U75258 ( .A(n72640), .B(n72639), .Y(n72641) );
  NAND2X1 U75259 ( .A(n72642), .B(n72641), .Y(n72709) );
  INVX1 U75260 ( .A(n72709), .Y(n72720) );
  NOR2X1 U75261 ( .A(n72660), .B(n72720), .Y(n72643) );
  NAND2X1 U75262 ( .A(n72643), .B(n72719), .Y(n72651) );
  NOR2X1 U75263 ( .A(n39427), .B(n38189), .Y(n72648) );
  NAND2X1 U75264 ( .A(n72646), .B(n40456), .Y(n72647) );
  NAND2X1 U75265 ( .A(n72648), .B(n72647), .Y(n72649) );
  NAND2X1 U75266 ( .A(n72721), .B(n72649), .Y(n72650) );
  NOR2X1 U75267 ( .A(n72651), .B(n72650), .Y(n72664) );
  NOR2X1 U75268 ( .A(n38818), .B(n43715), .Y(n72659) );
  NOR2X1 U75269 ( .A(n43707), .B(n72665), .Y(n72652) );
  NOR2X1 U75270 ( .A(n38189), .B(n72652), .Y(n72656) );
  NOR2X1 U75271 ( .A(n36569), .B(n41273), .Y(n72653) );
  NAND2X1 U75272 ( .A(n72653), .B(n38887), .Y(n72654) );
  NAND2X1 U75273 ( .A(n40455), .B(n72654), .Y(n72655) );
  NOR2X1 U75274 ( .A(n72659), .B(n72658), .Y(n72662) );
  NOR2X1 U75275 ( .A(n72661), .B(n72662), .Y(n72663) );
  NAND2X1 U75276 ( .A(n72666), .B(n43697), .Y(n72667) );
  XNOR2X1 U75277 ( .A(n72669), .B(n72668), .Y(n72670) );
  XNOR2X1 U75278 ( .A(n72671), .B(n72670), .Y(n72672) );
  XNOR2X1 U75279 ( .A(n72672), .B(n41142), .Y(n72673) );
  XNOR2X1 U75280 ( .A(n72674), .B(n72673), .Y(n72681) );
  INVX1 U75281 ( .A(n72681), .Y(n72676) );
  NOR2X1 U75282 ( .A(n43678), .B(n39177), .Y(n72679) );
  NOR2X1 U75283 ( .A(n72679), .B(n72678), .Y(n72680) );
  NOR2X1 U75284 ( .A(n40304), .B(n72680), .Y(n72683) );
  NAND2X1 U75285 ( .A(n43677), .B(n72681), .Y(n72682) );
  NAND2X1 U75286 ( .A(n43506), .B(n72692), .Y(n72684) );
  NOR2X1 U75287 ( .A(n39252), .B(n72684), .Y(n72691) );
  NAND2X1 U75288 ( .A(n43506), .B(n72685), .Y(n72687) );
  NAND2X1 U75289 ( .A(n72687), .B(n72686), .Y(n72688) );
  NOR2X1 U75290 ( .A(n72689), .B(n72688), .Y(n72690) );
  NOR2X1 U75291 ( .A(n43507), .B(n72692), .Y(n72693) );
  NOR2X1 U75292 ( .A(n39252), .B(n72693), .Y(n72695) );
  NAND2X1 U75293 ( .A(n72703), .B(n72697), .Y(n72696) );
  NOR2X1 U75294 ( .A(n72701), .B(n72696), .Y(n72707) );
  NOR2X1 U75295 ( .A(n72703), .B(n72697), .Y(n72705) );
  NAND2X1 U75296 ( .A(n72699), .B(n43698), .Y(n72700) );
  NAND2X1 U75297 ( .A(n72701), .B(n72700), .Y(n72702) );
  NOR2X1 U75298 ( .A(n72703), .B(n72702), .Y(n72704) );
  OR2X1 U75299 ( .A(n72705), .B(n72704), .Y(n72706) );
  NOR2X1 U75300 ( .A(n72707), .B(n72706), .Y(n72727) );
  NAND2X1 U75301 ( .A(n72709), .B(n43711), .Y(n72710) );
  NOR2X1 U75302 ( .A(n40457), .B(n72710), .Y(n72711) );
  NOR2X1 U75303 ( .A(n43718), .B(n72711), .Y(n72712) );
  NAND2X1 U75304 ( .A(n72712), .B(n72727), .Y(n72714) );
  NOR2X1 U75305 ( .A(n36551), .B(n72716), .Y(n72717) );
  NOR2X1 U75306 ( .A(n72720), .B(n72718), .Y(n72726) );
  NAND2X1 U75307 ( .A(n72720), .B(n72719), .Y(n72724) );
  NAND2X1 U75308 ( .A(n72722), .B(n72721), .Y(n72723) );
  NOR2X1 U75309 ( .A(n72724), .B(n72723), .Y(n72725) );
  NAND2X1 U75310 ( .A(n38972), .B(n44631), .Y(n13841) );
  NAND2X1 U75311 ( .A(n72732), .B(n72731), .Y(n10607) );
  NOR2X1 U75312 ( .A(n36719), .B(n72732), .Y(n72733) );
  NAND2X1 U75313 ( .A(n43729), .B(n72733), .Y(n10608) );
  NOR2X1 U75314 ( .A(n43520), .B(n72796), .Y(n72735) );
  NOR2X1 U75315 ( .A(n43722), .B(n72797), .Y(n72734) );
  NOR2X1 U75316 ( .A(n72735), .B(n72734), .Y(n72738) );
  INVX1 U75317 ( .A(n72736), .Y(n72800) );
  NAND2X1 U75318 ( .A(n72800), .B(n43791), .Y(n72737) );
  NAND2X1 U75319 ( .A(n72738), .B(n72737), .Y(u_lsu_N224) );
  INVX1 U75320 ( .A(n72739), .Y(n72824) );
  NAND2X1 U75321 ( .A(n72824), .B(n43792), .Y(n72743) );
  INVX1 U75322 ( .A(n72740), .Y(n72826) );
  NAND2X1 U75323 ( .A(n72826), .B(n40488), .Y(n72742) );
  NAND2X1 U75324 ( .A(n72743), .B(n72742), .Y(u_lsu_N208) );
  NOR2X1 U75325 ( .A(n43503), .B(n72796), .Y(n72745) );
  NOR2X1 U75326 ( .A(n40477), .B(n72797), .Y(n72744) );
  NOR2X1 U75327 ( .A(n72745), .B(n72744), .Y(n72747) );
  NAND2X1 U75328 ( .A(n72800), .B(n43744), .Y(n72746) );
  NAND2X1 U75329 ( .A(n72747), .B(n72746), .Y(u_lsu_N223) );
  NOR2X1 U75330 ( .A(n43498), .B(n72796), .Y(n72749) );
  NOR2X1 U75331 ( .A(n40460), .B(n72797), .Y(n72748) );
  NOR2X1 U75332 ( .A(n72749), .B(n72748), .Y(n72751) );
  NAND2X1 U75333 ( .A(n72800), .B(n43766), .Y(n72750) );
  NAND2X1 U75334 ( .A(n72751), .B(n72750), .Y(u_lsu_N222) );
  NOR2X1 U75335 ( .A(n43480), .B(n72796), .Y(n72753) );
  NOR2X1 U75336 ( .A(n43740), .B(n72797), .Y(n72752) );
  NOR2X1 U75337 ( .A(n72753), .B(n72752), .Y(n72755) );
  NAND2X1 U75338 ( .A(n72800), .B(n43732), .Y(n72754) );
  NAND2X1 U75339 ( .A(n72755), .B(n72754), .Y(u_lsu_N218) );
  INVX1 U75340 ( .A(n72756), .Y(n72814) );
  NAND2X1 U75341 ( .A(n72814), .B(n43732), .Y(n72758) );
  NAND2X1 U75342 ( .A(n72816), .B(n43725), .Y(n72757) );
  NAND2X1 U75343 ( .A(n72758), .B(n72757), .Y(u_lsu_N210) );
  NAND2X1 U75344 ( .A(n72824), .B(n43731), .Y(n72762) );
  NAND2X1 U75345 ( .A(n72826), .B(n43736), .Y(n72761) );
  NAND2X1 U75346 ( .A(n72762), .B(n72761), .Y(u_lsu_N202) );
  NAND2X1 U75347 ( .A(n72814), .B(n43744), .Y(n72764) );
  NAND2X1 U75348 ( .A(n72816), .B(n42712), .Y(n72763) );
  NAND2X1 U75349 ( .A(n72764), .B(n72763), .Y(u_lsu_N215) );
  NAND2X1 U75350 ( .A(n72824), .B(n43742), .Y(n72768) );
  NAND2X1 U75351 ( .A(n72826), .B(n40470), .Y(n72767) );
  NAND2X1 U75352 ( .A(n72768), .B(n72767), .Y(u_lsu_N207) );
  NAND2X1 U75353 ( .A(n72814), .B(n43752), .Y(n72770) );
  NAND2X1 U75354 ( .A(n72816), .B(n42636), .Y(n72769) );
  NAND2X1 U75355 ( .A(n72770), .B(n72769), .Y(u_lsu_N211) );
  NOR2X1 U75356 ( .A(n43485), .B(n72796), .Y(n72772) );
  NOR2X1 U75357 ( .A(n43760), .B(n72797), .Y(n72771) );
  NOR2X1 U75358 ( .A(n72772), .B(n72771), .Y(n72774) );
  NAND2X1 U75359 ( .A(n72800), .B(n43752), .Y(n72773) );
  NAND2X1 U75360 ( .A(n72774), .B(n72773), .Y(u_lsu_N219) );
  NOR2X1 U75361 ( .A(n43495), .B(n72796), .Y(n72776) );
  NOR2X1 U75362 ( .A(n43813), .B(n72797), .Y(n72775) );
  NOR2X1 U75363 ( .A(n72776), .B(n72775), .Y(n72778) );
  NAND2X1 U75364 ( .A(n72800), .B(n43805), .Y(n72777) );
  NAND2X1 U75365 ( .A(n72778), .B(n72777), .Y(u_lsu_N221) );
  NAND2X1 U75366 ( .A(n72824), .B(n43752), .Y(n72782) );
  NAND2X1 U75367 ( .A(n72826), .B(n43759), .Y(n72781) );
  NAND2X1 U75368 ( .A(n72782), .B(n72781), .Y(u_lsu_N203) );
  NAND2X1 U75369 ( .A(n72814), .B(n43766), .Y(n72785) );
  NAND2X1 U75370 ( .A(n72816), .B(n42653), .Y(n72784) );
  NAND2X1 U75371 ( .A(n72785), .B(n72784), .Y(u_lsu_N214) );
  NAND2X1 U75372 ( .A(n72824), .B(n39525), .Y(n72789) );
  NAND2X1 U75373 ( .A(n72826), .B(n40466), .Y(n72788) );
  NAND2X1 U75374 ( .A(n72789), .B(n72788), .Y(u_lsu_N206) );
  NAND2X1 U75375 ( .A(n72814), .B(n43815), .Y(n72791) );
  NAND2X1 U75376 ( .A(n72816), .B(n40259), .Y(n72790) );
  NAND2X1 U75377 ( .A(n72791), .B(n72790), .Y(u_lsu_N212) );
  NOR2X1 U75378 ( .A(n43489), .B(n72796), .Y(n72793) );
  NOR2X1 U75379 ( .A(n43822), .B(n72797), .Y(n72792) );
  NOR2X1 U75380 ( .A(n72793), .B(n72792), .Y(n72795) );
  NAND2X1 U75381 ( .A(n72800), .B(n43816), .Y(n72794) );
  NAND2X1 U75382 ( .A(n72795), .B(n72794), .Y(u_lsu_N220) );
  NOR2X1 U75383 ( .A(n39083), .B(n72796), .Y(n72799) );
  NOR2X1 U75384 ( .A(n43789), .B(n72797), .Y(n72798) );
  NOR2X1 U75385 ( .A(n72799), .B(n72798), .Y(n72802) );
  NAND2X1 U75386 ( .A(n72800), .B(n43781), .Y(n72801) );
  NAND2X1 U75387 ( .A(n72802), .B(n72801), .Y(u_lsu_N225) );
  NAND2X1 U75388 ( .A(n72814), .B(n39163), .Y(n72805) );
  NAND2X1 U75389 ( .A(n72816), .B(n43774), .Y(n72804) );
  NAND2X1 U75390 ( .A(n72805), .B(n72804), .Y(u_lsu_N217) );
  NAND2X1 U75391 ( .A(n72824), .B(n43780), .Y(n72809) );
  NAND2X1 U75392 ( .A(n72826), .B(n43788), .Y(n72808) );
  NAND2X1 U75393 ( .A(n72809), .B(n72808), .Y(u_lsu_N209) );
  NAND2X1 U75394 ( .A(n72814), .B(n43792), .Y(n72813) );
  NAND2X1 U75395 ( .A(n72816), .B(n43796), .Y(n72812) );
  NAND2X1 U75396 ( .A(n72813), .B(n72812), .Y(u_lsu_N216) );
  NAND2X1 U75397 ( .A(n72814), .B(n43805), .Y(n72818) );
  NAND2X1 U75398 ( .A(n72816), .B(n43798), .Y(n72817) );
  NAND2X1 U75399 ( .A(n72818), .B(n72817), .Y(u_lsu_N213) );
  NAND2X1 U75400 ( .A(n72824), .B(n43804), .Y(n72822) );
  NAND2X1 U75401 ( .A(n72826), .B(n72820), .Y(n72821) );
  NAND2X1 U75402 ( .A(n72822), .B(n72821), .Y(u_lsu_N205) );
  NAND2X1 U75403 ( .A(n72824), .B(n43815), .Y(n72828) );
  NAND2X1 U75404 ( .A(n72826), .B(n43820), .Y(n72827) );
  NAND2X1 U75405 ( .A(n72828), .B(n72827), .Y(u_lsu_N204) );
  NAND2X1 U75406 ( .A(n43825), .B(n73274), .Y(n72830) );
  NAND2X1 U75407 ( .A(u_csr_csr_stvec_q[11]), .B(n72830), .Y(n72832) );
  NAND2X1 U75408 ( .A(n42140), .B(n43963), .Y(n72831) );
  NAND2X1 U75409 ( .A(n72832), .B(n72831), .Y(u_csr_csr_stvec_r[11]) );
  OR2X1 U75410 ( .A(n72834), .B(n72833), .Y(n72835) );
  NAND2X1 U75411 ( .A(n43829), .B(n73274), .Y(n72836) );
  NAND2X1 U75412 ( .A(u_csr_csr_sscratch_q[11]), .B(n72836), .Y(n72838) );
  NAND2X1 U75413 ( .A(n42212), .B(n43963), .Y(n72837) );
  NAND2X1 U75414 ( .A(n72838), .B(n72837), .Y(u_csr_csr_sscratch_r[11]) );
  NOR2X1 U75415 ( .A(n72839), .B(n37353), .Y(n72845) );
  NAND2X1 U75416 ( .A(n72840), .B(n28235), .Y(n72841) );
  NAND2X1 U75417 ( .A(n72841), .B(n474), .Y(n72843) );
  NAND2X1 U75418 ( .A(n72843), .B(n72842), .Y(n72844) );
  NAND2X1 U75419 ( .A(n72845), .B(n72844), .Y(u_csr_N3472) );
  NAND2X1 U75420 ( .A(n43825), .B(n73186), .Y(n72846) );
  NAND2X1 U75421 ( .A(u_csr_csr_stvec_q[10]), .B(n72846), .Y(n72848) );
  NAND2X1 U75422 ( .A(n42140), .B(n43861), .Y(n72847) );
  NAND2X1 U75423 ( .A(n72848), .B(n72847), .Y(u_csr_csr_stvec_r[10]) );
  NAND2X1 U75424 ( .A(n43825), .B(n73267), .Y(n72849) );
  NAND2X1 U75425 ( .A(u_csr_csr_stvec_q[12]), .B(n72849), .Y(n72851) );
  NAND2X1 U75426 ( .A(n42140), .B(n43953), .Y(n72850) );
  NAND2X1 U75427 ( .A(n72851), .B(n72850), .Y(u_csr_csr_stvec_r[12]) );
  NAND2X1 U75428 ( .A(n43824), .B(n73193), .Y(n72852) );
  NAND2X1 U75429 ( .A(u_csr_csr_stvec_q[13]), .B(n72852), .Y(n72854) );
  NAND2X1 U75430 ( .A(n43827), .B(n43871), .Y(n72853) );
  NAND2X1 U75431 ( .A(n72854), .B(n72853), .Y(u_csr_csr_stvec_r[13]) );
  NAND2X1 U75432 ( .A(n43824), .B(n73200), .Y(n72855) );
  NAND2X1 U75433 ( .A(u_csr_csr_stvec_q[14]), .B(n72855), .Y(n72857) );
  NAND2X1 U75434 ( .A(n43827), .B(n43880), .Y(n72856) );
  NAND2X1 U75435 ( .A(n72857), .B(n72856), .Y(u_csr_csr_stvec_r[14]) );
  NAND2X1 U75436 ( .A(n43824), .B(n73207), .Y(n72858) );
  NAND2X1 U75437 ( .A(u_csr_csr_stvec_q[15]), .B(n72858), .Y(n72860) );
  NAND2X1 U75438 ( .A(n43827), .B(n43890), .Y(n72859) );
  NAND2X1 U75439 ( .A(n72860), .B(n72859), .Y(u_csr_csr_stvec_r[15]) );
  NAND2X1 U75440 ( .A(n43824), .B(n73214), .Y(n72861) );
  NAND2X1 U75441 ( .A(u_csr_csr_stvec_q[16]), .B(n72861), .Y(n72863) );
  NAND2X1 U75442 ( .A(n43827), .B(n43899), .Y(n72862) );
  NAND2X1 U75443 ( .A(n72863), .B(n72862), .Y(u_csr_csr_stvec_r[16]) );
  NAND2X1 U75444 ( .A(n43824), .B(n73222), .Y(n72864) );
  NAND2X1 U75445 ( .A(u_csr_csr_stvec_q[17]), .B(n72864), .Y(n72866) );
  NAND2X1 U75446 ( .A(n43827), .B(n43904), .Y(n72865) );
  NAND2X1 U75447 ( .A(n72866), .B(n72865), .Y(u_csr_csr_stvec_r[17]) );
  NAND2X1 U75448 ( .A(n43824), .B(n73230), .Y(n72867) );
  NAND2X1 U75449 ( .A(u_csr_csr_stvec_q[18]), .B(n72867), .Y(n72869) );
  NAND2X1 U75450 ( .A(n43827), .B(n43912), .Y(n72868) );
  NAND2X1 U75451 ( .A(n72869), .B(n72868), .Y(u_csr_csr_stvec_r[18]) );
  NAND2X1 U75452 ( .A(n43824), .B(n73238), .Y(n72870) );
  NAND2X1 U75453 ( .A(u_csr_csr_stvec_q[19]), .B(n72870), .Y(n72872) );
  NAND2X1 U75454 ( .A(n43827), .B(n43921), .Y(n72871) );
  NAND2X1 U75455 ( .A(n72872), .B(n72871), .Y(u_csr_csr_stvec_r[19]) );
  NAND2X1 U75456 ( .A(n43824), .B(n73245), .Y(n72873) );
  NAND2X1 U75457 ( .A(u_csr_csr_stvec_q[20]), .B(n72873), .Y(n72875) );
  NAND2X1 U75458 ( .A(n43827), .B(n43928), .Y(n72874) );
  NAND2X1 U75459 ( .A(n72875), .B(n72874), .Y(u_csr_csr_stvec_r[20]) );
  NAND2X1 U75460 ( .A(n43824), .B(n73252), .Y(n72876) );
  NAND2X1 U75461 ( .A(u_csr_csr_stvec_q[21]), .B(n72876), .Y(n72878) );
  NAND2X1 U75462 ( .A(n43827), .B(n43934), .Y(n72877) );
  NAND2X1 U75463 ( .A(n72878), .B(n72877), .Y(u_csr_csr_stvec_r[21]) );
  NAND2X1 U75464 ( .A(n43947), .B(n44083), .Y(n73260) );
  NAND2X1 U75465 ( .A(n43824), .B(n73260), .Y(n72879) );
  NAND2X1 U75466 ( .A(u_csr_csr_stvec_q[22]), .B(n72879), .Y(n72881) );
  NAND2X1 U75467 ( .A(n43827), .B(n43943), .Y(n72880) );
  NAND2X1 U75468 ( .A(n72881), .B(n72880), .Y(u_csr_csr_stvec_r[22]) );
  NAND2X1 U75469 ( .A(n43978), .B(n44083), .Y(n73281) );
  NAND2X1 U75470 ( .A(n43824), .B(n73281), .Y(n72882) );
  NAND2X1 U75471 ( .A(u_csr_csr_stvec_q[23]), .B(n72882), .Y(n72884) );
  NAND2X1 U75472 ( .A(n43827), .B(n43972), .Y(n72883) );
  NAND2X1 U75473 ( .A(n72884), .B(n72883), .Y(u_csr_csr_stvec_r[23]) );
  NAND2X1 U75474 ( .A(n43987), .B(n44083), .Y(n73288) );
  NAND2X1 U75475 ( .A(n43824), .B(n73288), .Y(n72885) );
  NAND2X1 U75476 ( .A(u_csr_csr_stvec_q[24]), .B(n72885), .Y(n72887) );
  NAND2X1 U75477 ( .A(n43827), .B(n43983), .Y(n72886) );
  NAND2X1 U75478 ( .A(n72887), .B(n72886), .Y(u_csr_csr_stvec_r[24]) );
  NAND2X1 U75479 ( .A(n43996), .B(n44083), .Y(n73295) );
  NAND2X1 U75480 ( .A(n43823), .B(n73295), .Y(n72888) );
  NAND2X1 U75481 ( .A(u_csr_csr_stvec_q[25]), .B(n72888), .Y(n72890) );
  NAND2X1 U75482 ( .A(n43826), .B(n43992), .Y(n72889) );
  NAND2X1 U75483 ( .A(n72890), .B(n72889), .Y(u_csr_csr_stvec_r[25]) );
  NAND2X1 U75484 ( .A(n44006), .B(n44082), .Y(n73302) );
  NAND2X1 U75485 ( .A(n43823), .B(n73302), .Y(n72891) );
  NAND2X1 U75486 ( .A(u_csr_csr_stvec_q[26]), .B(n72891), .Y(n72893) );
  NAND2X1 U75487 ( .A(n43826), .B(n43999), .Y(n72892) );
  NAND2X1 U75488 ( .A(n72893), .B(n72892), .Y(u_csr_csr_stvec_r[26]) );
  NAND2X1 U75489 ( .A(n44013), .B(n44082), .Y(n73309) );
  NAND2X1 U75490 ( .A(n43823), .B(n73309), .Y(n72894) );
  NAND2X1 U75491 ( .A(u_csr_csr_stvec_q[27]), .B(n72894), .Y(n72896) );
  NAND2X1 U75492 ( .A(n43826), .B(n44007), .Y(n72895) );
  NAND2X1 U75493 ( .A(n72896), .B(n72895), .Y(u_csr_csr_stvec_r[27]) );
  NAND2X1 U75494 ( .A(n44020), .B(n44082), .Y(n73317) );
  NAND2X1 U75495 ( .A(n43823), .B(n73317), .Y(n72897) );
  NAND2X1 U75496 ( .A(u_csr_csr_stvec_q[28]), .B(n72897), .Y(n72899) );
  NAND2X1 U75497 ( .A(n43826), .B(n44016), .Y(n72898) );
  NAND2X1 U75498 ( .A(n72899), .B(n72898), .Y(u_csr_csr_stvec_r[28]) );
  NAND2X1 U75499 ( .A(n44028), .B(n44082), .Y(n73324) );
  NAND2X1 U75500 ( .A(n43823), .B(n73324), .Y(n72900) );
  NAND2X1 U75501 ( .A(u_csr_csr_stvec_q[29]), .B(n72900), .Y(n72902) );
  NAND2X1 U75502 ( .A(n43826), .B(n44024), .Y(n72901) );
  NAND2X1 U75503 ( .A(n72902), .B(n72901), .Y(u_csr_csr_stvec_r[29]) );
  NAND2X1 U75504 ( .A(n44053), .B(n44082), .Y(n73331) );
  NAND2X1 U75505 ( .A(n43823), .B(n73331), .Y(n72903) );
  NAND2X1 U75506 ( .A(u_csr_csr_stvec_q[30]), .B(n72903), .Y(n72905) );
  NAND2X1 U75507 ( .A(n43826), .B(n44047), .Y(n72904) );
  NAND2X1 U75508 ( .A(n72905), .B(n72904), .Y(u_csr_csr_stvec_r[30]) );
  NAND2X1 U75509 ( .A(n43823), .B(n73338), .Y(n72906) );
  NAND2X1 U75510 ( .A(u_csr_csr_stvec_q[31]), .B(n72906), .Y(n72908) );
  NAND2X1 U75511 ( .A(n43826), .B(n44054), .Y(n72907) );
  NAND2X1 U75512 ( .A(n72908), .B(n72907), .Y(u_csr_csr_stvec_r[31]) );
  NAND2X1 U75513 ( .A(n43823), .B(n73345), .Y(n72909) );
  NAND2X1 U75514 ( .A(u_csr_csr_stvec_q[5]), .B(n72909), .Y(n72911) );
  NAND2X1 U75515 ( .A(n43826), .B(n39942), .Y(n72910) );
  NAND2X1 U75516 ( .A(n72911), .B(n72910), .Y(u_csr_csr_stvec_r[5]) );
  NAND2X1 U75517 ( .A(n43823), .B(n73170), .Y(n72912) );
  NAND2X1 U75518 ( .A(u_csr_csr_stvec_q[6]), .B(n72912), .Y(n72914) );
  NAND2X1 U75519 ( .A(n43826), .B(n43841), .Y(n72913) );
  NAND2X1 U75520 ( .A(n72914), .B(n72913), .Y(u_csr_csr_stvec_r[6]) );
  NAND2X1 U75521 ( .A(n43823), .B(n73352), .Y(n72915) );
  NAND2X1 U75522 ( .A(u_csr_csr_stvec_q[7]), .B(n72915), .Y(n72917) );
  NAND2X1 U75523 ( .A(n43826), .B(n38382), .Y(n72916) );
  NAND2X1 U75524 ( .A(n72917), .B(n72916), .Y(u_csr_csr_stvec_r[7]) );
  NAND2X1 U75525 ( .A(n43823), .B(n73359), .Y(n72918) );
  NAND2X1 U75526 ( .A(u_csr_csr_stvec_q[8]), .B(n72918), .Y(n72920) );
  NAND2X1 U75527 ( .A(n43826), .B(n44036), .Y(n72919) );
  NAND2X1 U75528 ( .A(n72920), .B(n72919), .Y(u_csr_csr_stvec_r[8]) );
  NAND2X1 U75529 ( .A(n43823), .B(n73179), .Y(n72921) );
  NAND2X1 U75530 ( .A(u_csr_csr_stvec_q[9]), .B(n72921), .Y(n72923) );
  NAND2X1 U75531 ( .A(n43826), .B(n43852), .Y(n72922) );
  NAND2X1 U75532 ( .A(n72923), .B(n72922), .Y(u_csr_csr_stvec_r[9]) );
  NAND2X1 U75533 ( .A(n43829), .B(n73186), .Y(n72924) );
  NAND2X1 U75534 ( .A(u_csr_csr_sscratch_q[10]), .B(n72924), .Y(n72926) );
  NAND2X1 U75535 ( .A(n42212), .B(n43861), .Y(n72925) );
  NAND2X1 U75536 ( .A(n72926), .B(n72925), .Y(u_csr_csr_sscratch_r[10]) );
  NAND2X1 U75537 ( .A(n43829), .B(n73267), .Y(n72927) );
  NAND2X1 U75538 ( .A(u_csr_csr_sscratch_q[12]), .B(n72927), .Y(n72929) );
  NAND2X1 U75539 ( .A(n42212), .B(n43953), .Y(n72928) );
  NAND2X1 U75540 ( .A(n72929), .B(n72928), .Y(u_csr_csr_sscratch_r[12]) );
  NAND2X1 U75541 ( .A(n43829), .B(n73193), .Y(n72930) );
  NAND2X1 U75542 ( .A(u_csr_csr_sscratch_q[13]), .B(n72930), .Y(n72932) );
  NAND2X1 U75543 ( .A(n43833), .B(n43871), .Y(n72931) );
  NAND2X1 U75544 ( .A(n72932), .B(n72931), .Y(u_csr_csr_sscratch_r[13]) );
  NAND2X1 U75545 ( .A(n43829), .B(n73200), .Y(n72933) );
  NAND2X1 U75546 ( .A(u_csr_csr_sscratch_q[14]), .B(n72933), .Y(n72935) );
  NAND2X1 U75547 ( .A(n43833), .B(n43880), .Y(n72934) );
  NAND2X1 U75548 ( .A(n72935), .B(n72934), .Y(u_csr_csr_sscratch_r[14]) );
  NAND2X1 U75549 ( .A(n43829), .B(n73207), .Y(n72936) );
  NAND2X1 U75550 ( .A(u_csr_csr_sscratch_q[15]), .B(n72936), .Y(n72938) );
  NAND2X1 U75551 ( .A(n43833), .B(n43890), .Y(n72937) );
  NAND2X1 U75552 ( .A(n72938), .B(n72937), .Y(u_csr_csr_sscratch_r[15]) );
  NAND2X1 U75553 ( .A(n43829), .B(n73214), .Y(n72939) );
  NAND2X1 U75554 ( .A(u_csr_csr_sscratch_q[16]), .B(n72939), .Y(n72941) );
  NAND2X1 U75555 ( .A(n43833), .B(n43899), .Y(n72940) );
  NAND2X1 U75556 ( .A(n72941), .B(n72940), .Y(u_csr_csr_sscratch_r[16]) );
  NAND2X1 U75557 ( .A(n43829), .B(n73222), .Y(n72942) );
  NAND2X1 U75558 ( .A(u_csr_csr_sscratch_q[17]), .B(n72942), .Y(n72944) );
  NAND2X1 U75559 ( .A(n43833), .B(n43904), .Y(n72943) );
  NAND2X1 U75560 ( .A(n72944), .B(n72943), .Y(u_csr_csr_sscratch_r[17]) );
  NAND2X1 U75561 ( .A(n43829), .B(n73230), .Y(n72945) );
  NAND2X1 U75562 ( .A(u_csr_csr_sscratch_q[18]), .B(n72945), .Y(n72947) );
  NAND2X1 U75563 ( .A(n43833), .B(n43912), .Y(n72946) );
  NAND2X1 U75564 ( .A(n72947), .B(n72946), .Y(u_csr_csr_sscratch_r[18]) );
  NAND2X1 U75565 ( .A(n43829), .B(n73238), .Y(n72948) );
  NAND2X1 U75566 ( .A(u_csr_csr_sscratch_q[19]), .B(n72948), .Y(n72950) );
  NAND2X1 U75567 ( .A(n43833), .B(n43921), .Y(n72949) );
  NAND2X1 U75568 ( .A(n72950), .B(n72949), .Y(u_csr_csr_sscratch_r[19]) );
  NAND2X1 U75569 ( .A(n43829), .B(n73245), .Y(n72951) );
  NAND2X1 U75570 ( .A(u_csr_csr_sscratch_q[20]), .B(n72951), .Y(n72953) );
  NAND2X1 U75571 ( .A(n43833), .B(n43929), .Y(n72952) );
  NAND2X1 U75572 ( .A(n72953), .B(n72952), .Y(u_csr_csr_sscratch_r[20]) );
  NAND2X1 U75573 ( .A(n43829), .B(n73252), .Y(n72954) );
  NAND2X1 U75574 ( .A(u_csr_csr_sscratch_q[21]), .B(n72954), .Y(n72956) );
  NAND2X1 U75575 ( .A(n43833), .B(n43933), .Y(n72955) );
  NAND2X1 U75576 ( .A(n72956), .B(n72955), .Y(u_csr_csr_sscratch_r[21]) );
  NAND2X1 U75577 ( .A(n43830), .B(n73260), .Y(n72957) );
  NAND2X1 U75578 ( .A(u_csr_csr_sscratch_q[22]), .B(n72957), .Y(n72959) );
  NAND2X1 U75579 ( .A(n43833), .B(n43943), .Y(n72958) );
  NAND2X1 U75580 ( .A(n72959), .B(n72958), .Y(u_csr_csr_sscratch_r[22]) );
  NAND2X1 U75581 ( .A(n43830), .B(n73281), .Y(n72960) );
  NAND2X1 U75582 ( .A(u_csr_csr_sscratch_q[23]), .B(n72960), .Y(n72962) );
  NAND2X1 U75583 ( .A(n43833), .B(n43972), .Y(n72961) );
  NAND2X1 U75584 ( .A(n72962), .B(n72961), .Y(u_csr_csr_sscratch_r[23]) );
  NAND2X1 U75585 ( .A(n43830), .B(n73288), .Y(n72963) );
  NAND2X1 U75586 ( .A(u_csr_csr_sscratch_q[24]), .B(n72963), .Y(n72965) );
  NAND2X1 U75587 ( .A(n43833), .B(n43982), .Y(n72964) );
  NAND2X1 U75588 ( .A(n72965), .B(n72964), .Y(u_csr_csr_sscratch_r[24]) );
  NAND2X1 U75589 ( .A(n43830), .B(n73295), .Y(n72966) );
  NAND2X1 U75590 ( .A(u_csr_csr_sscratch_q[25]), .B(n72966), .Y(n72968) );
  NAND2X1 U75591 ( .A(n43832), .B(n43991), .Y(n72967) );
  NAND2X1 U75592 ( .A(n72968), .B(n72967), .Y(u_csr_csr_sscratch_r[25]) );
  NAND2X1 U75593 ( .A(n43830), .B(n73302), .Y(n72969) );
  NAND2X1 U75594 ( .A(u_csr_csr_sscratch_q[26]), .B(n72969), .Y(n72971) );
  NAND2X1 U75595 ( .A(n43832), .B(n43999), .Y(n72970) );
  NAND2X1 U75596 ( .A(n72971), .B(n72970), .Y(u_csr_csr_sscratch_r[26]) );
  NAND2X1 U75597 ( .A(n43830), .B(n73309), .Y(n72972) );
  NAND2X1 U75598 ( .A(u_csr_csr_sscratch_q[27]), .B(n72972), .Y(n72974) );
  NAND2X1 U75599 ( .A(n43832), .B(n44007), .Y(n72973) );
  NAND2X1 U75600 ( .A(n72974), .B(n72973), .Y(u_csr_csr_sscratch_r[27]) );
  NAND2X1 U75601 ( .A(n43830), .B(n73317), .Y(n72975) );
  NAND2X1 U75602 ( .A(u_csr_csr_sscratch_q[28]), .B(n72975), .Y(n72977) );
  NAND2X1 U75603 ( .A(n43832), .B(n44016), .Y(n72976) );
  NAND2X1 U75604 ( .A(n72977), .B(n72976), .Y(u_csr_csr_sscratch_r[28]) );
  NAND2X1 U75605 ( .A(n43830), .B(n73324), .Y(n72978) );
  NAND2X1 U75606 ( .A(u_csr_csr_sscratch_q[29]), .B(n72978), .Y(n72980) );
  NAND2X1 U75607 ( .A(n43832), .B(n44024), .Y(n72979) );
  NAND2X1 U75608 ( .A(n72980), .B(n72979), .Y(u_csr_csr_sscratch_r[29]) );
  NAND2X1 U75609 ( .A(n43830), .B(n73331), .Y(n72981) );
  NAND2X1 U75610 ( .A(u_csr_csr_sscratch_q[30]), .B(n72981), .Y(n72983) );
  NAND2X1 U75611 ( .A(n43832), .B(n44047), .Y(n72982) );
  NAND2X1 U75612 ( .A(n72983), .B(n72982), .Y(u_csr_csr_sscratch_r[30]) );
  NAND2X1 U75613 ( .A(n43830), .B(n73338), .Y(n72984) );
  NAND2X1 U75614 ( .A(u_csr_csr_sscratch_q[31]), .B(n72984), .Y(n72986) );
  NAND2X1 U75615 ( .A(n43832), .B(n44054), .Y(n72985) );
  NAND2X1 U75616 ( .A(n72986), .B(n72985), .Y(u_csr_csr_sscratch_r[31]) );
  NAND2X1 U75617 ( .A(n43830), .B(n73345), .Y(n72987) );
  NAND2X1 U75618 ( .A(u_csr_csr_sscratch_q[5]), .B(n72987), .Y(n72989) );
  NAND2X1 U75619 ( .A(n43832), .B(n39942), .Y(n72988) );
  NAND2X1 U75620 ( .A(n72989), .B(n72988), .Y(u_csr_csr_sscratch_r[5]) );
  NAND2X1 U75621 ( .A(n43830), .B(n73170), .Y(n72990) );
  NAND2X1 U75622 ( .A(u_csr_csr_sscratch_q[6]), .B(n72990), .Y(n72992) );
  NAND2X1 U75623 ( .A(n43832), .B(n43842), .Y(n72991) );
  NAND2X1 U75624 ( .A(n72992), .B(n72991), .Y(u_csr_csr_sscratch_r[6]) );
  NAND2X1 U75625 ( .A(n43831), .B(n73352), .Y(n72993) );
  NAND2X1 U75626 ( .A(u_csr_csr_sscratch_q[7]), .B(n72993), .Y(n72995) );
  NAND2X1 U75627 ( .A(n43832), .B(n38381), .Y(n72994) );
  NAND2X1 U75628 ( .A(n72995), .B(n72994), .Y(u_csr_csr_sscratch_r[7]) );
  NAND2X1 U75629 ( .A(n43831), .B(n73359), .Y(n72996) );
  NAND2X1 U75630 ( .A(u_csr_csr_sscratch_q[8]), .B(n72996), .Y(n72998) );
  NAND2X1 U75631 ( .A(n43832), .B(n44037), .Y(n72997) );
  NAND2X1 U75632 ( .A(n72998), .B(n72997), .Y(u_csr_csr_sscratch_r[8]) );
  NAND2X1 U75633 ( .A(n43831), .B(n73179), .Y(n72999) );
  NAND2X1 U75634 ( .A(u_csr_csr_sscratch_q[9]), .B(n72999), .Y(n73001) );
  NAND2X1 U75635 ( .A(n43832), .B(n43852), .Y(n73000) );
  NAND2X1 U75636 ( .A(n73001), .B(n73000), .Y(u_csr_csr_sscratch_r[9]) );
  NAND2X1 U75637 ( .A(n26335), .B(n73281), .Y(n73002) );
  NAND2X1 U75638 ( .A(u_csr_csr_sr_q_23), .B(n73002), .Y(n73005) );
  INVX1 U75639 ( .A(n73003), .Y(n73028) );
  NAND2X1 U75640 ( .A(n73028), .B(n43972), .Y(n73004) );
  NAND2X1 U75641 ( .A(n73005), .B(n73004), .Y(u_csr_csr_sr_r[23]) );
  NAND2X1 U75642 ( .A(n26335), .B(n73288), .Y(n73006) );
  NAND2X1 U75643 ( .A(u_csr_csr_sr_q_24), .B(n73006), .Y(n73008) );
  NAND2X1 U75644 ( .A(n73028), .B(n43983), .Y(n73007) );
  NAND2X1 U75645 ( .A(n73008), .B(n73007), .Y(u_csr_csr_sr_r[24]) );
  NAND2X1 U75646 ( .A(n26335), .B(n73295), .Y(n73009) );
  NAND2X1 U75647 ( .A(u_csr_csr_sr_q_25), .B(n73009), .Y(n73011) );
  NAND2X1 U75648 ( .A(n73028), .B(n43991), .Y(n73010) );
  NAND2X1 U75649 ( .A(n73011), .B(n73010), .Y(u_csr_csr_sr_r[25]) );
  NAND2X1 U75650 ( .A(n26335), .B(n73302), .Y(n73012) );
  NAND2X1 U75651 ( .A(u_csr_csr_sr_q_26), .B(n73012), .Y(n73014) );
  NAND2X1 U75652 ( .A(n73028), .B(n43999), .Y(n73013) );
  NAND2X1 U75653 ( .A(n73014), .B(n73013), .Y(u_csr_csr_sr_r[26]) );
  NAND2X1 U75654 ( .A(n26335), .B(n73309), .Y(n73015) );
  NAND2X1 U75655 ( .A(u_csr_csr_sr_q_27), .B(n73015), .Y(n73017) );
  NAND2X1 U75656 ( .A(n73028), .B(n44007), .Y(n73016) );
  NAND2X1 U75657 ( .A(n73017), .B(n73016), .Y(u_csr_csr_sr_r[27]) );
  NAND2X1 U75658 ( .A(n26335), .B(n73317), .Y(n73018) );
  NAND2X1 U75659 ( .A(u_csr_csr_sr_q_28), .B(n73018), .Y(n73020) );
  NAND2X1 U75660 ( .A(n73028), .B(n44016), .Y(n73019) );
  NAND2X1 U75661 ( .A(n73020), .B(n73019), .Y(u_csr_csr_sr_r[28]) );
  NAND2X1 U75662 ( .A(n26335), .B(n73324), .Y(n73021) );
  NAND2X1 U75663 ( .A(u_csr_csr_sr_q_29), .B(n73021), .Y(n73023) );
  NAND2X1 U75664 ( .A(n73028), .B(n44024), .Y(n73022) );
  NAND2X1 U75665 ( .A(n73023), .B(n73022), .Y(u_csr_csr_sr_r[29]) );
  NAND2X1 U75666 ( .A(n26335), .B(n73331), .Y(n73024) );
  NAND2X1 U75667 ( .A(u_csr_csr_sr_q_30), .B(n73024), .Y(n73026) );
  NAND2X1 U75668 ( .A(n73028), .B(n44047), .Y(n73025) );
  NAND2X1 U75669 ( .A(n73026), .B(n73025), .Y(u_csr_csr_sr_r[30]) );
  NAND2X1 U75670 ( .A(n26335), .B(n73338), .Y(n73027) );
  NAND2X1 U75671 ( .A(u_csr_csr_sr_q_31), .B(n73027), .Y(n73030) );
  NAND2X1 U75672 ( .A(n73028), .B(n44054), .Y(n73029) );
  NAND2X1 U75673 ( .A(n73030), .B(n73029), .Y(u_csr_csr_sr_r[31]) );
  NAND2X1 U75674 ( .A(n44278), .B(n73245), .Y(n73032) );
  NAND2X1 U75675 ( .A(n73032), .B(n73031), .Y(n73034) );
  NAND2X1 U75676 ( .A(n43835), .B(n43928), .Y(n73033) );
  NAND2X1 U75677 ( .A(n73034), .B(n73033), .Y(u_csr_csr_satp_r[20]) );
  NAND2X1 U75678 ( .A(n44278), .B(n73252), .Y(n73035) );
  NAND2X1 U75679 ( .A(n73035), .B(n73567), .Y(n73037) );
  NAND2X1 U75680 ( .A(n43835), .B(n43933), .Y(n73036) );
  NAND2X1 U75681 ( .A(n73037), .B(n73036), .Y(u_csr_csr_satp_r[21]) );
  NAND2X1 U75682 ( .A(n44278), .B(n73260), .Y(n73038) );
  NAND2X1 U75683 ( .A(n73038), .B(n73566), .Y(n73040) );
  NAND2X1 U75684 ( .A(n43835), .B(n43943), .Y(n73039) );
  NAND2X1 U75685 ( .A(n73040), .B(n73039), .Y(u_csr_csr_satp_r[22]) );
  NAND2X1 U75686 ( .A(n44278), .B(n73281), .Y(n73041) );
  NAND2X1 U75687 ( .A(n73041), .B(n73565), .Y(n73043) );
  NAND2X1 U75688 ( .A(n43835), .B(n43973), .Y(n73042) );
  NAND2X1 U75689 ( .A(n73043), .B(n73042), .Y(u_csr_csr_satp_r[23]) );
  NAND2X1 U75690 ( .A(n44278), .B(n73288), .Y(n73044) );
  NAND2X1 U75691 ( .A(n73044), .B(n73564), .Y(n73046) );
  NAND2X1 U75692 ( .A(n43835), .B(n43982), .Y(n73045) );
  NAND2X1 U75693 ( .A(n73046), .B(n73045), .Y(u_csr_csr_satp_r[24]) );
  NAND2X1 U75694 ( .A(n44278), .B(n73295), .Y(n73047) );
  NAND2X1 U75695 ( .A(n73047), .B(n73563), .Y(n73049) );
  NAND2X1 U75696 ( .A(n43835), .B(n43991), .Y(n73048) );
  NAND2X1 U75697 ( .A(n73049), .B(n73048), .Y(u_csr_csr_satp_r[25]) );
  NAND2X1 U75698 ( .A(n44278), .B(n73302), .Y(n73050) );
  NAND2X1 U75699 ( .A(n73050), .B(n73562), .Y(n73052) );
  NAND2X1 U75700 ( .A(n43835), .B(n43999), .Y(n73051) );
  NAND2X1 U75701 ( .A(n73052), .B(n73051), .Y(u_csr_csr_satp_r[26]) );
  NAND2X1 U75702 ( .A(n44278), .B(n73309), .Y(n73053) );
  NAND2X1 U75703 ( .A(n73053), .B(n73561), .Y(n73055) );
  NAND2X1 U75704 ( .A(n43835), .B(n44007), .Y(n73054) );
  NAND2X1 U75705 ( .A(n73055), .B(n73054), .Y(u_csr_csr_satp_r[27]) );
  NAND2X1 U75706 ( .A(n44278), .B(n73317), .Y(n73056) );
  NAND2X1 U75707 ( .A(n73056), .B(n73560), .Y(n73058) );
  NAND2X1 U75708 ( .A(n43835), .B(n44016), .Y(n73057) );
  NAND2X1 U75709 ( .A(n73058), .B(n73057), .Y(u_csr_csr_satp_r[28]) );
  NAND2X1 U75710 ( .A(n44278), .B(n73324), .Y(n73059) );
  NAND2X1 U75711 ( .A(n73059), .B(n73559), .Y(n73061) );
  NAND2X1 U75712 ( .A(n43835), .B(n44024), .Y(n73060) );
  NAND2X1 U75713 ( .A(n73061), .B(n73060), .Y(u_csr_csr_satp_r[29]) );
  NAND2X1 U75714 ( .A(n44278), .B(n73331), .Y(n73063) );
  NAND2X1 U75715 ( .A(n73063), .B(n73062), .Y(n73065) );
  NAND2X1 U75716 ( .A(n43835), .B(n44047), .Y(n73064) );
  NAND2X1 U75717 ( .A(n73065), .B(n73064), .Y(u_csr_csr_satp_r[30]) );
  NAND2X1 U75718 ( .A(n28567), .B(n73170), .Y(n73066) );
  NAND2X1 U75719 ( .A(u_csr_csr_sr_q[6]), .B(n73066), .Y(n73068) );
  NAND2X1 U75720 ( .A(n37344), .B(n43842), .Y(n73067) );
  NAND2X1 U75721 ( .A(n73068), .B(n73067), .Y(u_csr_N2379) );
  NAND2X1 U75722 ( .A(n28567), .B(n73179), .Y(n73069) );
  NAND2X1 U75723 ( .A(u_csr_csr_sr_q[9]), .B(n73069), .Y(n73071) );
  NAND2X1 U75724 ( .A(n37344), .B(n43852), .Y(n73070) );
  NAND2X1 U75725 ( .A(n73071), .B(n73070), .Y(u_csr_N2382) );
  NAND2X1 U75726 ( .A(n28567), .B(n73186), .Y(n73072) );
  NAND2X1 U75727 ( .A(u_csr_csr_sr_q[10]), .B(n73072), .Y(n73074) );
  NAND2X1 U75728 ( .A(n37344), .B(n43861), .Y(n73073) );
  NAND2X1 U75729 ( .A(n73074), .B(n73073), .Y(u_csr_N2383) );
  NAND2X1 U75730 ( .A(n28567), .B(n73193), .Y(n73075) );
  NAND2X1 U75731 ( .A(u_csr_csr_sr_q[13]), .B(n73075), .Y(n73077) );
  NAND2X1 U75732 ( .A(n37344), .B(n43871), .Y(n73076) );
  NAND2X1 U75733 ( .A(n73077), .B(n73076), .Y(u_csr_N2386) );
  NAND2X1 U75734 ( .A(n28567), .B(n73200), .Y(n73078) );
  NAND2X1 U75735 ( .A(u_csr_csr_sr_q[14]), .B(n73078), .Y(n73080) );
  NAND2X1 U75736 ( .A(n37344), .B(n43880), .Y(n73079) );
  NAND2X1 U75737 ( .A(n73080), .B(n73079), .Y(u_csr_N2387) );
  NAND2X1 U75738 ( .A(n28567), .B(n73207), .Y(n73081) );
  NAND2X1 U75739 ( .A(u_csr_csr_sr_q[15]), .B(n73081), .Y(n73083) );
  NAND2X1 U75740 ( .A(n37344), .B(n43890), .Y(n73082) );
  NAND2X1 U75741 ( .A(n73083), .B(n73082), .Y(u_csr_N2388) );
  NAND2X1 U75742 ( .A(n28567), .B(n73214), .Y(n73084) );
  NAND2X1 U75743 ( .A(u_csr_csr_sr_q[16]), .B(n73084), .Y(n73086) );
  NAND2X1 U75744 ( .A(n37344), .B(n43899), .Y(n73085) );
  NAND2X1 U75745 ( .A(n73086), .B(n73085), .Y(u_csr_N2389) );
  NAND2X1 U75746 ( .A(n28567), .B(n73222), .Y(n73087) );
  NAND2X1 U75747 ( .A(u_csr_csr_sr_q[17]), .B(n73087), .Y(n73089) );
  NAND2X1 U75748 ( .A(n37344), .B(n43904), .Y(n73088) );
  NAND2X1 U75749 ( .A(n73089), .B(n73088), .Y(u_csr_N2390) );
  NAND2X1 U75750 ( .A(n28567), .B(n73238), .Y(n73090) );
  NAND2X1 U75751 ( .A(u_csr_csr_sr_q_19), .B(n73090), .Y(n73092) );
  NAND2X1 U75752 ( .A(n37344), .B(n43921), .Y(n73091) );
  NAND2X1 U75753 ( .A(n73092), .B(n73091), .Y(u_csr_N2392) );
  NAND2X1 U75754 ( .A(n28567), .B(n73245), .Y(n73093) );
  NAND2X1 U75755 ( .A(u_csr_csr_sr_q_20), .B(n73093), .Y(n73095) );
  NAND2X1 U75756 ( .A(n37344), .B(n43928), .Y(n73094) );
  NAND2X1 U75757 ( .A(n73095), .B(n73094), .Y(u_csr_N2393) );
  NAND2X1 U75758 ( .A(n28567), .B(n73252), .Y(n73096) );
  NAND2X1 U75759 ( .A(u_csr_csr_sr_q_21), .B(n73096), .Y(n73098) );
  NAND2X1 U75760 ( .A(n37344), .B(n43934), .Y(n73097) );
  NAND2X1 U75761 ( .A(n73098), .B(n73097), .Y(u_csr_N2394) );
  NAND2X1 U75762 ( .A(n28567), .B(n73260), .Y(n73099) );
  NAND2X1 U75763 ( .A(u_csr_csr_sr_q_22), .B(n73099), .Y(n73101) );
  NAND2X1 U75764 ( .A(n37344), .B(n43942), .Y(n73100) );
  NAND2X1 U75765 ( .A(n73101), .B(n73100), .Y(u_csr_N2395) );
  NAND2X1 U75766 ( .A(n27407), .B(n73134), .Y(n73102) );
  NAND2X1 U75767 ( .A(u_csr_csr_mideleg_q[9]), .B(n73102), .Y(n73104) );
  NAND2X1 U75768 ( .A(n42214), .B(n43851), .Y(n73103) );
  NAND2X1 U75769 ( .A(n73104), .B(n73103), .Y(u_csr_csr_mideleg_r[9]) );
  NAND2X1 U75770 ( .A(n43003), .B(n44040), .Y(n73138) );
  NAND2X1 U75771 ( .A(n27407), .B(n73138), .Y(n73105) );
  NAND2X1 U75772 ( .A(u_csr_csr_mideleg_q[8]), .B(n73105), .Y(n73107) );
  NAND2X1 U75773 ( .A(n42214), .B(n44036), .Y(n73106) );
  NAND2X1 U75774 ( .A(n73107), .B(n73106), .Y(u_csr_csr_mideleg_r[8]) );
  NAND2X1 U75775 ( .A(n27407), .B(n73142), .Y(n73108) );
  NAND2X1 U75776 ( .A(u_csr_csr_mideleg_q[7]), .B(n73108), .Y(n73110) );
  NAND2X1 U75777 ( .A(n42214), .B(n38378), .Y(n73109) );
  NAND2X1 U75778 ( .A(n73110), .B(n73109), .Y(u_csr_csr_mideleg_r[7]) );
  NAND2X1 U75779 ( .A(n43004), .B(n43847), .Y(n73146) );
  NAND2X1 U75780 ( .A(n27407), .B(n73146), .Y(n73111) );
  NAND2X1 U75781 ( .A(u_csr_csr_mideleg_q[6]), .B(n73111), .Y(n73113) );
  NAND2X1 U75782 ( .A(n42214), .B(n43841), .Y(n73112) );
  NAND2X1 U75783 ( .A(n73113), .B(n73112), .Y(u_csr_csr_mideleg_r[6]) );
  NAND2X1 U75784 ( .A(n27407), .B(n73114), .Y(n73115) );
  NAND2X1 U75785 ( .A(u_csr_csr_mideleg_q[15]), .B(n73115), .Y(n73117) );
  NAND2X1 U75786 ( .A(n42214), .B(n43890), .Y(n73116) );
  NAND2X1 U75787 ( .A(n73117), .B(n73116), .Y(u_csr_csr_mideleg_r[15]) );
  NAND2X1 U75788 ( .A(n43002), .B(n43885), .Y(n73150) );
  NAND2X1 U75789 ( .A(n27407), .B(n73150), .Y(n73118) );
  NAND2X1 U75790 ( .A(u_csr_csr_mideleg_q[14]), .B(n73118), .Y(n73120) );
  NAND2X1 U75791 ( .A(n42214), .B(n43880), .Y(n73119) );
  NAND2X1 U75792 ( .A(n73120), .B(n73119), .Y(u_csr_csr_mideleg_r[14]) );
  NAND2X1 U75793 ( .A(n27407), .B(n73121), .Y(n73122) );
  NAND2X1 U75794 ( .A(u_csr_csr_mideleg_q[13]), .B(n73122), .Y(n73124) );
  NAND2X1 U75795 ( .A(n42214), .B(n43871), .Y(n73123) );
  NAND2X1 U75796 ( .A(n73124), .B(n73123), .Y(u_csr_csr_mideleg_r[13]) );
  NAND2X1 U75797 ( .A(n43003), .B(n43958), .Y(n73154) );
  NAND2X1 U75798 ( .A(n27407), .B(n73154), .Y(n73125) );
  NAND2X1 U75799 ( .A(u_csr_csr_mideleg_q[12]), .B(n73125), .Y(n73127) );
  NAND2X1 U75800 ( .A(n42214), .B(n43953), .Y(n73126) );
  NAND2X1 U75801 ( .A(n73127), .B(n73126), .Y(u_csr_csr_mideleg_r[12]) );
  NAND2X1 U75802 ( .A(n27407), .B(n73158), .Y(n73128) );
  NAND2X1 U75803 ( .A(u_csr_csr_mideleg_q[11]), .B(n73128), .Y(n73130) );
  NAND2X1 U75804 ( .A(n42214), .B(n43963), .Y(n73129) );
  NAND2X1 U75805 ( .A(n73130), .B(n73129), .Y(u_csr_csr_mideleg_r[11]) );
  NAND2X1 U75806 ( .A(n43004), .B(n43866), .Y(n73162) );
  NAND2X1 U75807 ( .A(n27407), .B(n73162), .Y(n73131) );
  NAND2X1 U75808 ( .A(u_csr_csr_mideleg_q[10]), .B(n73131), .Y(n73133) );
  NAND2X1 U75809 ( .A(n42214), .B(n43861), .Y(n73132) );
  NAND2X1 U75810 ( .A(n73133), .B(n73132), .Y(u_csr_csr_mideleg_r[10]) );
  NAND2X1 U75811 ( .A(n28045), .B(n73134), .Y(n73135) );
  NAND2X1 U75812 ( .A(u_csr_csr_medeleg_q[9]), .B(n73135), .Y(n73137) );
  NAND2X1 U75813 ( .A(n42143), .B(n43851), .Y(n73136) );
  NAND2X1 U75814 ( .A(n73137), .B(n73136), .Y(u_csr_csr_medeleg_r[9]) );
  NAND2X1 U75815 ( .A(n28045), .B(n73138), .Y(n73139) );
  NAND2X1 U75816 ( .A(u_csr_csr_medeleg_q[8]), .B(n73139), .Y(n73141) );
  NAND2X1 U75817 ( .A(n42143), .B(n44036), .Y(n73140) );
  NAND2X1 U75818 ( .A(n73141), .B(n73140), .Y(u_csr_csr_medeleg_r[8]) );
  NAND2X1 U75819 ( .A(n28045), .B(n73142), .Y(n73143) );
  NAND2X1 U75820 ( .A(u_csr_csr_medeleg_q[7]), .B(n73143), .Y(n73145) );
  NAND2X1 U75821 ( .A(n42143), .B(n38379), .Y(n73144) );
  NAND2X1 U75822 ( .A(n73145), .B(n73144), .Y(u_csr_csr_medeleg_r[7]) );
  NAND2X1 U75823 ( .A(n28045), .B(n73146), .Y(n73147) );
  NAND2X1 U75824 ( .A(u_csr_csr_medeleg_q[6]), .B(n73147), .Y(n73149) );
  NAND2X1 U75825 ( .A(n42143), .B(n43842), .Y(n73148) );
  NAND2X1 U75826 ( .A(n73149), .B(n73148), .Y(u_csr_csr_medeleg_r[6]) );
  NAND2X1 U75827 ( .A(n28045), .B(n73150), .Y(n73151) );
  NAND2X1 U75828 ( .A(u_csr_csr_medeleg_q[14]), .B(n73151), .Y(n73153) );
  NAND2X1 U75829 ( .A(n42143), .B(n43880), .Y(n73152) );
  NAND2X1 U75830 ( .A(n73153), .B(n73152), .Y(u_csr_csr_medeleg_r[14]) );
  NAND2X1 U75831 ( .A(n28045), .B(n73154), .Y(n73155) );
  NAND2X1 U75832 ( .A(u_csr_csr_medeleg_q[12]), .B(n73155), .Y(n73157) );
  NAND2X1 U75833 ( .A(n42143), .B(n43953), .Y(n73156) );
  NAND2X1 U75834 ( .A(n73157), .B(n73156), .Y(u_csr_csr_medeleg_r[12]) );
  NAND2X1 U75835 ( .A(n28045), .B(n73158), .Y(n73159) );
  NAND2X1 U75836 ( .A(u_csr_csr_medeleg_q[11]), .B(n73159), .Y(n73161) );
  NAND2X1 U75837 ( .A(n42143), .B(n43963), .Y(n73160) );
  NAND2X1 U75838 ( .A(n73161), .B(n73160), .Y(u_csr_csr_medeleg_r[11]) );
  NAND2X1 U75839 ( .A(n28045), .B(n73162), .Y(n73163) );
  NAND2X1 U75840 ( .A(u_csr_csr_medeleg_q[10]), .B(n73163), .Y(n73165) );
  NAND2X1 U75841 ( .A(n42143), .B(n43861), .Y(n73164) );
  NAND2X1 U75842 ( .A(n73165), .B(n73164), .Y(u_csr_csr_medeleg_r[10]) );
  NAND2X1 U75843 ( .A(n44274), .B(n73170), .Y(n73166) );
  NAND2X1 U75844 ( .A(u_csr_csr_mscratch_q[6]), .B(n73166), .Y(n73169) );
  NAND2X1 U75845 ( .A(n42141), .B(n43841), .Y(n73168) );
  NAND2X1 U75846 ( .A(n73169), .B(n73168), .Y(u_csr_csr_mscratch_r[6]) );
  NAND2X1 U75847 ( .A(n44277), .B(n73170), .Y(n73171) );
  NAND2X1 U75848 ( .A(u_csr_csr_mtvec_q[6]), .B(n73171), .Y(n73175) );
  NAND2X1 U75849 ( .A(n42139), .B(n43842), .Y(n73174) );
  NAND2X1 U75850 ( .A(n73175), .B(n73174), .Y(u_csr_csr_mtvec_r[6]) );
  NAND2X1 U75851 ( .A(n44274), .B(n73179), .Y(n73176) );
  NAND2X1 U75852 ( .A(u_csr_csr_mscratch_q[9]), .B(n73176), .Y(n73178) );
  NAND2X1 U75853 ( .A(n42141), .B(n43851), .Y(n73177) );
  NAND2X1 U75854 ( .A(n73178), .B(n73177), .Y(u_csr_csr_mscratch_r[9]) );
  NAND2X1 U75855 ( .A(n44277), .B(n73179), .Y(n73180) );
  NAND2X1 U75856 ( .A(u_csr_csr_mtvec_q[9]), .B(n73180), .Y(n73182) );
  NAND2X1 U75857 ( .A(n42139), .B(n43852), .Y(n73181) );
  NAND2X1 U75858 ( .A(n73182), .B(n73181), .Y(u_csr_csr_mtvec_r[9]) );
  NAND2X1 U75859 ( .A(n44274), .B(n73186), .Y(n73183) );
  NAND2X1 U75860 ( .A(u_csr_csr_mscratch_q[10]), .B(n73183), .Y(n73185) );
  NAND2X1 U75861 ( .A(n42141), .B(n43861), .Y(n73184) );
  NAND2X1 U75862 ( .A(n73185), .B(n73184), .Y(u_csr_csr_mscratch_r[10]) );
  NAND2X1 U75863 ( .A(n44277), .B(n73186), .Y(n73187) );
  NAND2X1 U75864 ( .A(u_csr_csr_mtvec_q[10]), .B(n73187), .Y(n73189) );
  NAND2X1 U75865 ( .A(n42139), .B(n43861), .Y(n73188) );
  NAND2X1 U75866 ( .A(n73189), .B(n73188), .Y(u_csr_csr_mtvec_r[10]) );
  NAND2X1 U75867 ( .A(n44273), .B(n73193), .Y(n73190) );
  NAND2X1 U75868 ( .A(u_csr_csr_mscratch_q[13]), .B(n73190), .Y(n73192) );
  NAND2X1 U75869 ( .A(n44031), .B(n43871), .Y(n73191) );
  NAND2X1 U75870 ( .A(n73192), .B(n73191), .Y(u_csr_csr_mscratch_r[13]) );
  NAND2X1 U75871 ( .A(n44276), .B(n73193), .Y(n73194) );
  NAND2X1 U75872 ( .A(u_csr_csr_mtvec_q[13]), .B(n73194), .Y(n73196) );
  NAND2X1 U75873 ( .A(n44043), .B(n43871), .Y(n73195) );
  NAND2X1 U75874 ( .A(n73196), .B(n73195), .Y(u_csr_csr_mtvec_r[13]) );
  NAND2X1 U75875 ( .A(n44273), .B(n73200), .Y(n73197) );
  NAND2X1 U75876 ( .A(u_csr_csr_mscratch_q[14]), .B(n73197), .Y(n73199) );
  NAND2X1 U75877 ( .A(n44031), .B(n43880), .Y(n73198) );
  NAND2X1 U75878 ( .A(n73199), .B(n73198), .Y(u_csr_csr_mscratch_r[14]) );
  NAND2X1 U75879 ( .A(n44276), .B(n73200), .Y(n73201) );
  NAND2X1 U75880 ( .A(u_csr_csr_mtvec_q[14]), .B(n73201), .Y(n73203) );
  NAND2X1 U75881 ( .A(n44043), .B(n43880), .Y(n73202) );
  NAND2X1 U75882 ( .A(n73203), .B(n73202), .Y(u_csr_csr_mtvec_r[14]) );
  NAND2X1 U75883 ( .A(n44273), .B(n73207), .Y(n73204) );
  NAND2X1 U75884 ( .A(u_csr_csr_mscratch_q[15]), .B(n73204), .Y(n73206) );
  NAND2X1 U75885 ( .A(n44031), .B(n43890), .Y(n73205) );
  NAND2X1 U75886 ( .A(n73206), .B(n73205), .Y(u_csr_csr_mscratch_r[15]) );
  NAND2X1 U75887 ( .A(n44276), .B(n73207), .Y(n73208) );
  NAND2X1 U75888 ( .A(u_csr_csr_mtvec_q[15]), .B(n73208), .Y(n73210) );
  NAND2X1 U75889 ( .A(n44043), .B(n43891), .Y(n73209) );
  NAND2X1 U75890 ( .A(n73210), .B(n73209), .Y(u_csr_csr_mtvec_r[15]) );
  NAND2X1 U75891 ( .A(n44273), .B(n73214), .Y(n73211) );
  NAND2X1 U75892 ( .A(u_csr_csr_mscratch_q[16]), .B(n73211), .Y(n73213) );
  NAND2X1 U75893 ( .A(n44031), .B(n43899), .Y(n73212) );
  NAND2X1 U75894 ( .A(n73213), .B(n73212), .Y(u_csr_csr_mscratch_r[16]) );
  NAND2X1 U75895 ( .A(n44276), .B(n73214), .Y(n73215) );
  NAND2X1 U75896 ( .A(u_csr_csr_mtvec_q[16]), .B(n73215), .Y(n73218) );
  NAND2X1 U75897 ( .A(n44043), .B(n43898), .Y(n73217) );
  NAND2X1 U75898 ( .A(n73218), .B(n73217), .Y(u_csr_csr_mtvec_r[16]) );
  NAND2X1 U75899 ( .A(n44273), .B(n73222), .Y(n73219) );
  NAND2X1 U75900 ( .A(u_csr_csr_mscratch_q[17]), .B(n73219), .Y(n73221) );
  NAND2X1 U75901 ( .A(n44031), .B(n43904), .Y(n73220) );
  NAND2X1 U75902 ( .A(n73221), .B(n73220), .Y(u_csr_csr_mscratch_r[17]) );
  NAND2X1 U75903 ( .A(n44276), .B(n73222), .Y(n73223) );
  NAND2X1 U75904 ( .A(u_csr_csr_mtvec_q[17]), .B(n73223), .Y(n73226) );
  NAND2X1 U75905 ( .A(n44043), .B(n43903), .Y(n73225) );
  NAND2X1 U75906 ( .A(n73226), .B(n73225), .Y(u_csr_csr_mtvec_r[17]) );
  NAND2X1 U75907 ( .A(n44273), .B(n73230), .Y(n73227) );
  NAND2X1 U75908 ( .A(u_csr_csr_mscratch_q[18]), .B(n73227), .Y(n73229) );
  NAND2X1 U75909 ( .A(n44031), .B(n43912), .Y(n73228) );
  NAND2X1 U75910 ( .A(n73229), .B(n73228), .Y(u_csr_csr_mscratch_r[18]) );
  NAND2X1 U75911 ( .A(n44276), .B(n73230), .Y(n73231) );
  NAND2X1 U75912 ( .A(u_csr_csr_mtvec_q[18]), .B(n73231), .Y(n73234) );
  NAND2X1 U75913 ( .A(n44043), .B(n43911), .Y(n73233) );
  NAND2X1 U75914 ( .A(n73234), .B(n73233), .Y(u_csr_csr_mtvec_r[18]) );
  NAND2X1 U75915 ( .A(n44273), .B(n73238), .Y(n73235) );
  NAND2X1 U75916 ( .A(u_csr_csr_mscratch_q[19]), .B(n73235), .Y(n73237) );
  NAND2X1 U75917 ( .A(n44031), .B(n43921), .Y(n73236) );
  NAND2X1 U75918 ( .A(n73237), .B(n73236), .Y(u_csr_csr_mscratch_r[19]) );
  NAND2X1 U75919 ( .A(n44276), .B(n73238), .Y(n73239) );
  NAND2X1 U75920 ( .A(u_csr_csr_mtvec_q[19]), .B(n73239), .Y(n73241) );
  NAND2X1 U75921 ( .A(n44043), .B(n43920), .Y(n73240) );
  NAND2X1 U75922 ( .A(n73241), .B(n73240), .Y(u_csr_csr_mtvec_r[19]) );
  NAND2X1 U75923 ( .A(n44273), .B(n73245), .Y(n73242) );
  NAND2X1 U75924 ( .A(u_csr_csr_mscratch_q[20]), .B(n73242), .Y(n73244) );
  NAND2X1 U75925 ( .A(n44031), .B(n43928), .Y(n73243) );
  NAND2X1 U75926 ( .A(n73244), .B(n73243), .Y(u_csr_csr_mscratch_r[20]) );
  NAND2X1 U75927 ( .A(n44276), .B(n73245), .Y(n73246) );
  NAND2X1 U75928 ( .A(u_csr_csr_mtvec_q[20]), .B(n73246), .Y(n73248) );
  NAND2X1 U75929 ( .A(n44043), .B(n43929), .Y(n73247) );
  NAND2X1 U75930 ( .A(n73248), .B(n73247), .Y(u_csr_csr_mtvec_r[20]) );
  NAND2X1 U75931 ( .A(n44273), .B(n73252), .Y(n73249) );
  NAND2X1 U75932 ( .A(u_csr_csr_mscratch_q[21]), .B(n73249), .Y(n73251) );
  NAND2X1 U75933 ( .A(n44031), .B(n43933), .Y(n73250) );
  NAND2X1 U75934 ( .A(n73251), .B(n73250), .Y(u_csr_csr_mscratch_r[21]) );
  NAND2X1 U75935 ( .A(n44276), .B(n73252), .Y(n73253) );
  NAND2X1 U75936 ( .A(u_csr_csr_mtvec_q[21]), .B(n73253), .Y(n73256) );
  NAND2X1 U75937 ( .A(n44043), .B(n43934), .Y(n73255) );
  NAND2X1 U75938 ( .A(n73256), .B(n73255), .Y(u_csr_csr_mtvec_r[21]) );
  NAND2X1 U75939 ( .A(n44273), .B(n73260), .Y(n73257) );
  NAND2X1 U75940 ( .A(u_csr_csr_mscratch_q[22]), .B(n73257), .Y(n73259) );
  NAND2X1 U75941 ( .A(n44031), .B(n43942), .Y(n73258) );
  NAND2X1 U75942 ( .A(n73259), .B(n73258), .Y(u_csr_csr_mscratch_r[22]) );
  NAND2X1 U75943 ( .A(n44276), .B(n73260), .Y(n73261) );
  NAND2X1 U75944 ( .A(u_csr_csr_mtvec_q[22]), .B(n73261), .Y(n73263) );
  NAND2X1 U75945 ( .A(n44043), .B(n43943), .Y(n73262) );
  NAND2X1 U75946 ( .A(n73263), .B(n73262), .Y(u_csr_csr_mtvec_r[22]) );
  NAND2X1 U75947 ( .A(n44273), .B(n73267), .Y(n73264) );
  NAND2X1 U75948 ( .A(u_csr_csr_mscratch_q[12]), .B(n73264), .Y(n73266) );
  NAND2X1 U75949 ( .A(n44031), .B(n43953), .Y(n73265) );
  NAND2X1 U75950 ( .A(n73266), .B(n73265), .Y(u_csr_csr_mscratch_r[12]) );
  NAND2X1 U75951 ( .A(n44276), .B(n73267), .Y(n73268) );
  NAND2X1 U75952 ( .A(u_csr_csr_mtvec_q[12]), .B(n73268), .Y(n73270) );
  NAND2X1 U75953 ( .A(n44043), .B(n43954), .Y(n73269) );
  NAND2X1 U75954 ( .A(n73270), .B(n73269), .Y(u_csr_csr_mtvec_r[12]) );
  NAND2X1 U75955 ( .A(n44273), .B(n73274), .Y(n73271) );
  NAND2X1 U75956 ( .A(u_csr_csr_mscratch_q[11]), .B(n73271), .Y(n73273) );
  NAND2X1 U75957 ( .A(n44031), .B(n43963), .Y(n73272) );
  NAND2X1 U75958 ( .A(n73273), .B(n73272), .Y(u_csr_csr_mscratch_r[11]) );
  NAND2X1 U75959 ( .A(n44276), .B(n73274), .Y(n73275) );
  NAND2X1 U75960 ( .A(u_csr_csr_mtvec_q[11]), .B(n73275), .Y(n73277) );
  NAND2X1 U75961 ( .A(n44043), .B(n43964), .Y(n73276) );
  NAND2X1 U75962 ( .A(n73277), .B(n73276), .Y(u_csr_csr_mtvec_r[11]) );
  NAND2X1 U75963 ( .A(n44272), .B(n73281), .Y(n73278) );
  NAND2X1 U75964 ( .A(u_csr_csr_mscratch_q[23]), .B(n73278), .Y(n73280) );
  NAND2X1 U75965 ( .A(n44030), .B(n43972), .Y(n73279) );
  NAND2X1 U75966 ( .A(n73280), .B(n73279), .Y(u_csr_csr_mscratch_r[23]) );
  NAND2X1 U75967 ( .A(n44275), .B(n73281), .Y(n73282) );
  NAND2X1 U75968 ( .A(u_csr_csr_mtvec_q[23]), .B(n73282), .Y(n73284) );
  NAND2X1 U75969 ( .A(n44042), .B(n43973), .Y(n73283) );
  NAND2X1 U75970 ( .A(n73284), .B(n73283), .Y(u_csr_csr_mtvec_r[23]) );
  NAND2X1 U75971 ( .A(n44272), .B(n73288), .Y(n73285) );
  NAND2X1 U75972 ( .A(u_csr_csr_mscratch_q[24]), .B(n73285), .Y(n73287) );
  NAND2X1 U75973 ( .A(n44030), .B(n43982), .Y(n73286) );
  NAND2X1 U75974 ( .A(n73287), .B(n73286), .Y(u_csr_csr_mscratch_r[24]) );
  NAND2X1 U75975 ( .A(n44275), .B(n73288), .Y(n73289) );
  NAND2X1 U75976 ( .A(u_csr_csr_mtvec_q[24]), .B(n73289), .Y(n73291) );
  NAND2X1 U75977 ( .A(n44042), .B(n43982), .Y(n73290) );
  NAND2X1 U75978 ( .A(n73291), .B(n73290), .Y(u_csr_csr_mtvec_r[24]) );
  NAND2X1 U75979 ( .A(n44272), .B(n73295), .Y(n73292) );
  NAND2X1 U75980 ( .A(u_csr_csr_mscratch_q[25]), .B(n73292), .Y(n73294) );
  NAND2X1 U75981 ( .A(n44030), .B(n43991), .Y(n73293) );
  NAND2X1 U75982 ( .A(n73294), .B(n73293), .Y(u_csr_csr_mscratch_r[25]) );
  NAND2X1 U75983 ( .A(n44275), .B(n73295), .Y(n73296) );
  NAND2X1 U75984 ( .A(u_csr_csr_mtvec_q[25]), .B(n73296), .Y(n73298) );
  NAND2X1 U75985 ( .A(n44042), .B(n43993), .Y(n73297) );
  NAND2X1 U75986 ( .A(n73298), .B(n73297), .Y(u_csr_csr_mtvec_r[25]) );
  NAND2X1 U75987 ( .A(n44272), .B(n73302), .Y(n73299) );
  NAND2X1 U75988 ( .A(u_csr_csr_mscratch_q[26]), .B(n73299), .Y(n73301) );
  NAND2X1 U75989 ( .A(n44030), .B(n43999), .Y(n73300) );
  NAND2X1 U75990 ( .A(n73301), .B(n73300), .Y(u_csr_csr_mscratch_r[26]) );
  NAND2X1 U75991 ( .A(n44275), .B(n73302), .Y(n73303) );
  NAND2X1 U75992 ( .A(u_csr_csr_mtvec_q[26]), .B(n73303), .Y(n73305) );
  NAND2X1 U75993 ( .A(n44042), .B(n44001), .Y(n73304) );
  NAND2X1 U75994 ( .A(n73305), .B(n73304), .Y(u_csr_csr_mtvec_r[26]) );
  NAND2X1 U75995 ( .A(n44272), .B(n73309), .Y(n73306) );
  NAND2X1 U75996 ( .A(u_csr_csr_mscratch_q[27]), .B(n73306), .Y(n73308) );
  NAND2X1 U75997 ( .A(n44030), .B(n44007), .Y(n73307) );
  NAND2X1 U75998 ( .A(n73308), .B(n73307), .Y(u_csr_csr_mscratch_r[27]) );
  NAND2X1 U75999 ( .A(n44275), .B(n73309), .Y(n73310) );
  NAND2X1 U76000 ( .A(u_csr_csr_mtvec_q[27]), .B(n73310), .Y(n73313) );
  NAND2X1 U76001 ( .A(n44042), .B(n44009), .Y(n73312) );
  NAND2X1 U76002 ( .A(n73313), .B(n73312), .Y(u_csr_csr_mtvec_r[27]) );
  NAND2X1 U76003 ( .A(n44272), .B(n73317), .Y(n73314) );
  NAND2X1 U76004 ( .A(u_csr_csr_mscratch_q[28]), .B(n73314), .Y(n73316) );
  NAND2X1 U76005 ( .A(n44030), .B(n44016), .Y(n73315) );
  NAND2X1 U76006 ( .A(n73316), .B(n73315), .Y(u_csr_csr_mscratch_r[28]) );
  NAND2X1 U76007 ( .A(n44275), .B(n73317), .Y(n73318) );
  NAND2X1 U76008 ( .A(u_csr_csr_mtvec_q[28]), .B(n73318), .Y(n73320) );
  NAND2X1 U76009 ( .A(n44042), .B(n44018), .Y(n73319) );
  NAND2X1 U76010 ( .A(n73320), .B(n73319), .Y(u_csr_csr_mtvec_r[28]) );
  NAND2X1 U76011 ( .A(n44272), .B(n73324), .Y(n73321) );
  NAND2X1 U76012 ( .A(u_csr_csr_mscratch_q[29]), .B(n73321), .Y(n73323) );
  NAND2X1 U76013 ( .A(n44030), .B(n44024), .Y(n73322) );
  NAND2X1 U76014 ( .A(n73323), .B(n73322), .Y(u_csr_csr_mscratch_r[29]) );
  NAND2X1 U76015 ( .A(n44275), .B(n73324), .Y(n73325) );
  NAND2X1 U76016 ( .A(u_csr_csr_mtvec_q[29]), .B(n73325), .Y(n73327) );
  NAND2X1 U76017 ( .A(n44042), .B(n44026), .Y(n73326) );
  NAND2X1 U76018 ( .A(n73327), .B(n73326), .Y(u_csr_csr_mtvec_r[29]) );
  NAND2X1 U76019 ( .A(n44272), .B(n73331), .Y(n73328) );
  NAND2X1 U76020 ( .A(u_csr_csr_mscratch_q[30]), .B(n73328), .Y(n73330) );
  NAND2X1 U76021 ( .A(n44030), .B(n44047), .Y(n73329) );
  NAND2X1 U76022 ( .A(n73330), .B(n73329), .Y(u_csr_csr_mscratch_r[30]) );
  NAND2X1 U76023 ( .A(n44275), .B(n73331), .Y(n73332) );
  NAND2X1 U76024 ( .A(u_csr_csr_mtvec_q[30]), .B(n73332), .Y(n73334) );
  NAND2X1 U76025 ( .A(n44042), .B(n44047), .Y(n73333) );
  NAND2X1 U76026 ( .A(n73334), .B(n73333), .Y(u_csr_csr_mtvec_r[30]) );
  NAND2X1 U76027 ( .A(n44272), .B(n73338), .Y(n73335) );
  NAND2X1 U76028 ( .A(u_csr_csr_mscratch_q[31]), .B(n73335), .Y(n73337) );
  NAND2X1 U76029 ( .A(n44030), .B(n44054), .Y(n73336) );
  NAND2X1 U76030 ( .A(n73337), .B(n73336), .Y(u_csr_csr_mscratch_r[31]) );
  NAND2X1 U76031 ( .A(n44275), .B(n73338), .Y(n73339) );
  NAND2X1 U76032 ( .A(u_csr_csr_mtvec_q[31]), .B(n73339), .Y(n73341) );
  NAND2X1 U76033 ( .A(n44042), .B(n44054), .Y(n73340) );
  NAND2X1 U76034 ( .A(n73341), .B(n73340), .Y(u_csr_csr_mtvec_r[31]) );
  NAND2X1 U76035 ( .A(n44272), .B(n73345), .Y(n73342) );
  NAND2X1 U76036 ( .A(u_csr_csr_mscratch_q[5]), .B(n73342), .Y(n73344) );
  NAND2X1 U76037 ( .A(n44030), .B(n39943), .Y(n73343) );
  NAND2X1 U76038 ( .A(n73344), .B(n73343), .Y(u_csr_csr_mscratch_r[5]) );
  NAND2X1 U76039 ( .A(n44275), .B(n73345), .Y(n73346) );
  NAND2X1 U76040 ( .A(u_csr_csr_mtvec_q[5]), .B(n73346), .Y(n73348) );
  NAND2X1 U76041 ( .A(n44042), .B(n39938), .Y(n73347) );
  NAND2X1 U76042 ( .A(n73348), .B(n73347), .Y(u_csr_csr_mtvec_r[5]) );
  NAND2X1 U76043 ( .A(n44272), .B(n73352), .Y(n73349) );
  NAND2X1 U76044 ( .A(u_csr_csr_mscratch_q[7]), .B(n73349), .Y(n73351) );
  NAND2X1 U76045 ( .A(n44030), .B(n38380), .Y(n73350) );
  NAND2X1 U76046 ( .A(n73351), .B(n73350), .Y(u_csr_csr_mscratch_r[7]) );
  NAND2X1 U76047 ( .A(n44275), .B(n73352), .Y(n73353) );
  NAND2X1 U76048 ( .A(u_csr_csr_mtvec_q[7]), .B(n73353), .Y(n73355) );
  NAND2X1 U76049 ( .A(n44042), .B(n38383), .Y(n73354) );
  NAND2X1 U76050 ( .A(n73355), .B(n73354), .Y(u_csr_csr_mtvec_r[7]) );
  NAND2X1 U76051 ( .A(n44272), .B(n73359), .Y(n73356) );
  NAND2X1 U76052 ( .A(u_csr_csr_mscratch_q[8]), .B(n73356), .Y(n73358) );
  NAND2X1 U76053 ( .A(n44030), .B(n44036), .Y(n73357) );
  NAND2X1 U76054 ( .A(n73358), .B(n73357), .Y(u_csr_csr_mscratch_r[8]) );
  NAND2X1 U76055 ( .A(n44275), .B(n73359), .Y(n73360) );
  NAND2X1 U76056 ( .A(u_csr_csr_mtvec_q[8]), .B(n73360), .Y(n73362) );
  NAND2X1 U76057 ( .A(n44042), .B(n44037), .Y(n73361) );
  NAND2X1 U76058 ( .A(n73362), .B(n73361), .Y(u_csr_csr_mtvec_r[8]) );
  NAND2X1 U76059 ( .A(n17098), .B(n73363), .Y(n4705) );
  NAND2X1 U76060 ( .A(n73365), .B(n73364), .Y(n73371) );
  NOR2X1 U76061 ( .A(n73367), .B(n73366), .Y(n73369) );
  NAND2X1 U76062 ( .A(n73369), .B(n42675), .Y(n73370) );
  NOR2X1 U76063 ( .A(n73371), .B(n73370), .Y(u_lsu_N230) );
  NAND2X1 U76064 ( .A(opcode_opcode_w[7]), .B(n73374), .Y(n73372) );
  NAND2X1 U76065 ( .A(n28905), .B(n73372), .Y(n8510) );
  NAND2X1 U76066 ( .A(opcode_opcode_w[10]), .B(n73374), .Y(n73373) );
  NAND2X1 U76067 ( .A(n28911), .B(n73373), .Y(n8507) );
  NAND2X1 U76068 ( .A(opcode_opcode_w[11]), .B(n73374), .Y(n73375) );
  NAND2X1 U76069 ( .A(n28913), .B(n73375), .Y(n8506) );
  NOR2X1 U76070 ( .A(n44047), .B(n73376), .Y(n73377) );
  NAND2X1 U76071 ( .A(n44063), .B(n73377), .Y(n73378) );
  NAND2X1 U76072 ( .A(n73378), .B(n73383), .Y(n73380) );
  NAND2X1 U76073 ( .A(n73380), .B(n44056), .Y(n73381) );
  NAND2X1 U76074 ( .A(n14449), .B(n73381), .Y(u_muldiv_N263) );
  NAND2X1 U76075 ( .A(n73383), .B(n44064), .Y(n73385) );
  NAND2X1 U76076 ( .A(n73385), .B(n73384), .Y(n73386) );
  NAND2X1 U76077 ( .A(n14890), .B(n73386), .Y(u_muldiv_N232) );
  MX2X1 U76078 ( .A(n21), .B(u_mmu_itlb_entry_q[12]), .S0(n44073), .Y(
        mem_i_pc_o[12]) );
  MX2X1 U76079 ( .A(n9), .B(u_mmu_itlb_entry_q[13]), .S0(n44073), .Y(
        mem_i_pc_o[13]) );
  MX2X1 U76080 ( .A(n24), .B(u_mmu_itlb_entry_q[14]), .S0(n44073), .Y(
        mem_i_pc_o[14]) );
  MX2X1 U76081 ( .A(n22), .B(u_mmu_itlb_entry_q[15]), .S0(n44073), .Y(
        mem_i_pc_o[15]) );
  MX2X1 U76082 ( .A(n8), .B(u_mmu_itlb_entry_q[16]), .S0(n44073), .Y(
        mem_i_pc_o[16]) );
  MX2X1 U76083 ( .A(n6), .B(u_mmu_itlb_entry_q[17]), .S0(n44074), .Y(
        mem_i_pc_o[17]) );
  MX2X1 U76084 ( .A(n10), .B(u_mmu_itlb_entry_q[18]), .S0(n44074), .Y(
        mem_i_pc_o[18]) );
  MX2X1 U76085 ( .A(n20), .B(u_mmu_itlb_entry_q[19]), .S0(n44074), .Y(
        mem_i_pc_o[19]) );
  MX2X1 U76086 ( .A(n7), .B(u_mmu_itlb_entry_q[20]), .S0(n44074), .Y(
        mem_i_pc_o[20]) );
  MX2X1 U76087 ( .A(n12), .B(u_mmu_itlb_entry_q[21]), .S0(n44074), .Y(
        mem_i_pc_o[21]) );
  MX2X1 U76088 ( .A(n17), .B(u_mmu_itlb_entry_q[22]), .S0(n44074), .Y(
        mem_i_pc_o[22]) );
  MX2X1 U76089 ( .A(n15), .B(u_mmu_itlb_entry_q[23]), .S0(n44074), .Y(
        mem_i_pc_o[23]) );
  MX2X1 U76090 ( .A(n11), .B(u_mmu_itlb_entry_q[24]), .S0(n44074), .Y(
        mem_i_pc_o[24]) );
  MX2X1 U76091 ( .A(n23), .B(u_mmu_itlb_entry_q[25]), .S0(n44074), .Y(
        mem_i_pc_o[25]) );
  MX2X1 U76092 ( .A(n13), .B(u_mmu_itlb_entry_q[26]), .S0(n44074), .Y(
        mem_i_pc_o[26]) );
  MX2X1 U76093 ( .A(n19), .B(u_mmu_itlb_entry_q[27]), .S0(n44074), .Y(
        mem_i_pc_o[27]) );
  MX2X1 U76094 ( .A(n18), .B(u_mmu_itlb_entry_q[28]), .S0(n44074), .Y(
        mem_i_pc_o[28]) );
  MX2X1 U76095 ( .A(n16), .B(u_mmu_itlb_entry_q[30]), .S0(n44073), .Y(
        mem_i_pc_o[30]) );
  MX2X1 U76096 ( .A(\mmu_ifetch_pc_w[31] ), .B(u_mmu_itlb_entry_q[31]), .S0(
        n44074), .Y(mem_i_pc_o[31]) );
  NAND2X1 U76097 ( .A(n73387), .B(n24429), .Y(n73393) );
  NOR2X1 U76098 ( .A(n73389), .B(n73388), .Y(n73391) );
  NAND2X1 U76099 ( .A(n73391), .B(n73390), .Y(n73392) );
  NOR2X1 U76100 ( .A(n73393), .B(n73392), .Y(u_decode_N180) );
  NOR2X1 U76101 ( .A(n1877), .B(n44256), .Y(mem_d_req_tag_o[0]) );
  NOR2X1 U76102 ( .A(n1880), .B(n44256), .Y(mem_d_req_tag_o[3]) );
  NOR2X1 U76103 ( .A(n1881), .B(n44256), .Y(mem_d_req_tag_o[4]) );
endmodule
